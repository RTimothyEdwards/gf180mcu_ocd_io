magic
tech gf180mcuD
magscale 1 10
timestamp 1484609607
<< polysilicon >>
rect 73 65 157 84
rect 73 19 92 65
rect 138 19 157 65
rect 73 -76 157 19
<< polycontact >>
rect 92 19 138 65
<< metal1 >>
rect 0 65 236 76
rect 0 19 92 65
rect 138 19 236 65
rect 0 8 236 19
<< end >>
