magic
tech gf180mcuD
magscale 1 10
timestamp 1758818771
<< metal5 >>
rect 14000 70000 17000 71000
rect 17200 70000 20200 71000
rect 20400 70000 23400 71000
rect 23600 70000 25000 71000
rect 25200 70000 26600 71000
rect 26800 70000 29800 71000
rect 30000 70000 33000 71000
rect 33200 70000 36200 71000
rect 36400 70000 39400 71000
rect 39600 70000 41000 71000
rect 41200 70000 42600 71000
rect 42800 70000 45800 71000
rect 46000 70000 49000 71000
rect 49200 70000 50600 71000
rect 50800 70000 52200 71000
rect 52400 70000 53800 71000
rect 54000 70000 55400 71000
rect 55600 70000 57000 71000
rect 57200 70000 58600 71000
rect 58800 70000 60200 71000
rect 60400 70000 61800 71000
rect 62000 70000 63400 71000
rect 63600 70000 65000 71000
rect 65200 70000 66600 71000
rect 66800 70000 68200 71000
rect 68400 70000 69678 71000
rect 70000 68400 71000 69678
rect 70000 66800 71000 68200
rect 70000 65200 71000 66600
rect 70000 63600 71000 65000
rect 70000 62000 71000 63400
rect 70000 60400 71000 61800
rect 70000 58800 71000 60200
rect 70000 57200 71000 58600
rect 70000 55600 71000 57000
rect 70000 54000 71000 55400
rect 70000 52400 71000 53800
rect 70000 50800 71000 52200
rect 70000 49200 71000 50600
rect 70000 46000 71000 49000
rect 70000 42800 71000 45799
rect 70000 41200 71000 42600
rect 70000 39600 71000 41000
rect 70000 36400 71000 39400
rect 70000 33200 71000 36200
rect 70000 30000 71000 33000
rect 70000 26800 71000 29800
rect 70000 25200 71000 26600
rect 70000 23600 71000 25000
rect 70000 20400 71000 23400
rect 70000 17200 71000 20200
rect 70000 14000 71000 17000
use GF_NI_COR_BASE  GF_NI_COR_BASE_0
timestamp 1758749514
transform 1 0 12 0 1 0
box 13436 13361 70889 70890
use POWER_RAIL_COR  POWER_RAIL_COR_0
timestamp 1758726819
transform 1 0 0 0 1 0
box 13097 13097 71000 71000
<< labels >>
flabel metal5 s 70000 33200 71000 36200 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 70000 30000 71000 33000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 70000 26800 71000 29800 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 70000 23600 71000 25000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 70000 39600 71000 41000 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 70000 25200 71000 26600 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 70000 20400 71000 23400 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 70000 14000 71000 17000 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 70000 17200 71000 20200 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 70000 41200 71000 42600 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 70000 36400 71000 39400 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 36400 70000 39400 71000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 33200 70000 36200 71000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 30000 70000 33000 71000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 26800 70000 29800 71000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 25200 70000 26600 71000 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 23600 70000 25000 71000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 20400 70000 23400 71000 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 17200 70000 20200 71000 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 14000 70000 17000 71000 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 41200 70000 42600 71000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 39600 70000 41000 71000 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 65200 70000 66600 71000 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 63600 70000 65000 71000 0 FreeSans 1600 0 0 0 VSS
port 4 nsew ground bidirectional
flabel metal5 s 62000 70000 63400 71000 0 FreeSans 1600 0 0 0 VDD
port 3 nsew power bidirectional
flabel metal5 s 60400 70000 61800 71000 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 58800 70000 60200 71000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 57200 70000 58600 71000 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 55600 70000 57000 71000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 54000 70000 55400 71000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 52400 70000 53800 71000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 50800 70000 52200 71000 0 FreeSans 1600 0 0 0 VDD
port 3 nsew power bidirectional
flabel metal5 s 49200 70000 50600 71000 0 FreeSans 1600 0 0 0 VSS
port 4 nsew ground bidirectional
flabel metal5 s 46000 70000 49000 71000 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 42800 70000 45800 71000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 70000 66800 71000 68200 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 70000 62000 71000 63400 0 FreeSans 1600 0 0 0 VDD
port 3 nsew power bidirectional
flabel metal5 s 70000 58800 71000 60200 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 70000 55600 71000 57000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 70000 54000 71000 55400 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 70000 52400 71000 53800 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 70000 42800 71000 45799 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 70000 68400 71000 69678 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 70000 65200 71000 66600 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 70000 60400 71000 61800 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 70000 57200 71000 58600 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 70000 46000 71000 49000 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 68400 70000 69678 71000 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 66800 70000 68200 71000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 70000 50800 71000 52200 0 FreeSans 1600 0 0 0 VDD
port 3 nsew power bidirectional
flabel metal5 s 70000 49200 71000 50600 0 FreeSans 1600 0 0 0 VSS
port 4 nsew ground bidirectional
flabel metal5 s 70000 63600 71000 65000 0 FreeSans 1600 0 0 0 VSS
port 4 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 71000 71000
string LEFclass PAD SPACER
string LEFsymmetry X Y R90
string LEFsite GF_IO_Site
<< end >>
