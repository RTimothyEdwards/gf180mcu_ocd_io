magic
tech gf180mcuD
magscale 1 10
timestamp 1758724778
<< nwell >>
rect -3895 53660 -2673 54997
<< nsubdiff >>
rect -3812 54892 -2756 54914
rect -3812 53812 -3790 54892
rect -3744 54846 -3636 54892
rect -2932 54846 -2824 54892
rect -3744 54824 -2824 54846
rect -3744 53880 -3722 54824
rect -2846 53880 -2824 54824
rect -3744 53858 -2824 53880
rect -3744 53812 -3636 53858
rect -2932 53812 -2824 53858
rect -2778 53812 -2756 54892
rect -3812 53790 -2756 53812
<< nsubdiffcont >>
rect -3790 53812 -3744 54892
rect -3636 54846 -2932 54892
rect -3636 53812 -2932 53858
rect -2824 53812 -2778 54892
<< polysilicon >>
rect -3504 54601 -3344 54614
rect -3504 54555 -3447 54601
rect -3401 54555 -3344 54601
rect -3504 54512 -3344 54555
rect -3504 54149 -3344 54192
rect -3504 54103 -3447 54149
rect -3401 54103 -3344 54149
rect -3504 54090 -3344 54103
rect -3224 54601 -3064 54614
rect -3224 54555 -3167 54601
rect -3121 54555 -3064 54601
rect -3224 54512 -3064 54555
rect -3224 54149 -3064 54192
rect -3224 54103 -3167 54149
rect -3121 54103 -3064 54149
rect -3224 54090 -3064 54103
<< polycontact >>
rect -3447 54555 -3401 54601
rect -3447 54103 -3401 54149
rect -3167 54555 -3121 54601
rect -3167 54103 -3121 54149
<< ppolyres >>
rect -3504 54192 -3344 54512
rect -3224 54192 -3064 54512
<< metal1 >>
rect -3801 54892 -2767 54903
rect -3801 53869 -3790 54892
rect -3850 53812 -3790 53869
rect -3744 54846 -3636 54892
rect -2932 54846 -2824 54892
rect -3744 54835 -2824 54846
rect -3744 54160 -3733 54835
rect -3502 54601 -3320 54612
rect -3502 54555 -3447 54601
rect -3401 54555 -3320 54601
rect -3502 54544 -3320 54555
rect -3396 54432 -3320 54544
rect -3254 54601 -3066 54612
rect -3254 54555 -3167 54601
rect -3121 54555 -3066 54601
rect -3254 54544 -3066 54555
rect -3254 54432 -3178 54544
rect -2835 54160 -2824 54835
rect -3744 54149 -2824 54160
rect -3744 54103 -3447 54149
rect -3401 54103 -3167 54149
rect -3121 54103 -2824 54149
rect -3744 54092 -2824 54103
rect -3744 53869 -3733 54092
rect -2835 53869 -2824 54092
rect -3744 53858 -2824 53869
rect -3744 53812 -3636 53858
rect -2932 53812 -2824 53858
rect -2778 53869 -2767 54892
rect -2778 53812 -2720 53869
rect -3850 53660 -2720 53812
<< end >>
