magic
tech gf180mcuB
magscale 1 10
timestamp 1758807451
use 4LM_METAL_RAIL  4LM_METAL_RAIL_0
timestamp 1484609606
transform 1 0 0 0 1 0
box -32 13097 15032 69968
use Bondpad_4LM  Bondpad_4LM_0
timestamp 1484609606
transform 1 0 1100 0 1 0
box -400 0 13200 13065
<< properties >>
string FIXED_BBOX 0 13097 15000 70000
<< end >>
