# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_ocd_io__dvss
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_ocd_io__dvss 0 0 ;
  SIZE 75 BY 350 ;
  SYMMETRY X Y R90 ;
  SITE GF_IO_Site ;
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 74 102 75 117 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74 86 75 101 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74 70 75 85 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74 126 75 133 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74 198 75 205 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74 230 75 245 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74 246 75 253 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74 286 75 293 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74 302 75 309 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74 318 75 325 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74 326 75 333 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74 342 75 348.39 ;
    END
    PORT
        CLASS CORE ;
      LAYER Metal2 ;
        RECT 1.36 349 10.86 350 ;
    END
    PORT
        CLASS CORE ;
      LAYER Metal2 ;
        RECT 13.76 349 24.01 350 ;
    END
    PORT
        CLASS CORE ;
      LAYER Metal2 ;
        RECT 25.61 349 35.86 350 ;
    END
    PORT
        CLASS CORE ;
      LAYER Metal2 ;
        RECT 39.14 349 49.39 350 ;
    END
    PORT
        CLASS CORE ;
      LAYER Metal2 ;
        RECT 50.99 349 61.24 350 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 342 1 348.39 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 326 1 333 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 318 1 325 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 302 1 309 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 286 1 293 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 246 1 253 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 230 1 245 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 198 1 205 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 126 1 133 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 70 1 85 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 86 1 101 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 102 1 117 ;
    END
    PORT
        CLASS CORE ;
      LAYER Metal2 ;
        RECT 64.14 349 73.64 350 ;
    END
  END DVSS
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 74 118 75 125 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74 182 75 197 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74 166 75 181 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74 150 75 165 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74 134 75 149 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74 214 75 229 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74 206 75 213 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74 278 75 285 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74 270 75 277 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74 262 75 269 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74 294 75 301 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74 334 75 341 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 334 1 341 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 294 1 301 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 262 1 269 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 270 1 277 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 278 1 285 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 206 1 213 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 214 1 229 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 134 1 149 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 150 1 165 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 166 1 181 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 182 1 197 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 118 1 125 ;
    END
  END DVDD
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 74 254 75 261 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74 310 75 317 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 310 1 317 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 254 1 261 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      RECT 0 0 75 350 ;
    LAYER Metal2 ;
      POLYGON 75 350 73.92 350 73.92 348.72 63.86 348.72 63.86 350 61.52 350 61.52 348.72 50.71 348.72 50.71 350 49.67 350 49.67 348.72 38.86 348.72 38.86 350 36.14 350 36.14 348.72 25.33 348.72 25.33 350 24.29 350 24.29 348.72 13.48 348.72 13.48 350 11.14 350 11.14 348.72 1.08 348.72 1.08 350 0 350 0 0 75 0 ;
    LAYER Metal3 ;
      POLYGON 75 69.72 73.72 69.72 73.72 85.28 75 85.28 75 85.72 73.72 85.72 73.72 101.28 75 101.28 75 101.72 73.72 101.72 73.72 117.28 75 117.28 75 117.72 73.72 117.72 73.72 125.28 75 125.28 75 125.72 73.72 125.72 73.72 133.28 75 133.28 75 133.72 73.72 133.72 73.72 149.28 75 149.28 75 149.72 73.72 149.72 73.72 165.28 75 165.28 75 165.72 73.72 165.72 73.72 181.28 75 181.28 75 181.72 73.72 181.72 73.72 197.28 75 197.28 75 197.72 73.72 197.72 73.72 205.28 75 205.28 75 205.72 73.72 205.72 73.72 213.28 75 213.28 75 213.72 73.72 213.72 73.72 229.28 75 229.28 75 229.72 73.72 229.72 73.72 245.28 75 245.28 75 245.72 73.72 245.72 73.72 253.28 75 253.28 75 253.72 73.72 253.72 73.72 261.28 75 261.28 75 261.72 73.72 261.72 73.72 269.28 75 269.28 75 269.72 73.72 269.72 73.72 277.28 75 277.28 75 277.72 73.72 277.72 73.72 285.28 75 285.28 75 285.72 73.72 285.72 73.72 293.28 75 293.28 75 293.72 73.72 293.72 73.72 301.28 75 301.28 75 301.72 73.72 301.72 73.72 309.28 75 309.28 75 309.72 73.72 309.72 73.72 317.28 75 317.28 75 317.72 73.72 317.72 73.72 325.28 75 325.28 75 325.72 73.72 325.72 73.72 333.28 75 333.28 75 333.72 73.72 333.72 73.72 341.28 75 341.28 75 341.72 73.72 341.72 73.72 348.67 75 348.67 75 350 0 350 0 348.67 1.28 348.67 1.28 341.72 0 341.72 0 341.28 1.28 341.28 1.28 333.72 0 333.72 0 333.28 1.28 333.28 1.28 325.72 0 325.72 0 325.28 1.28 325.28 1.28 317.72 0 317.72 0 317.28 1.28 317.28 1.28 309.72 0 309.72 0 309.28 1.28 309.28 1.28 301.72 0 301.72 0 301.28 1.28 301.28 1.28 293.72 0 293.72 0 293.28 1.28 293.28 1.28 285.72 0 285.72 0 285.28 1.28 285.28 1.28 277.72 0 277.72 0 277.28 1.28 277.28 1.28 269.72 0 269.72 0 269.28 1.28 269.28 1.28 261.72 0 261.72 0 261.28 1.28 261.28 1.28 253.72 0 253.72 0 253.28 1.28 253.28 1.28 245.72 0 245.72 0 245.28 1.28 245.28 1.28 229.72 0 229.72 0 229.28 1.28 229.28 1.28 213.72 0 213.72 0 213.28 1.28 213.28 1.28 205.72 0 205.72 0 205.28 1.28 205.28 1.28 197.72 0 197.72 0 197.28 1.28 197.28 1.28 181.72 0 181.72 0 181.28 1.28 181.28 1.28 165.72 0 165.72 0 165.28 1.28 165.28 1.28 149.72 0 149.72 0 149.28 1.28 149.28 1.28 133.72 0 133.72 0 133.28 1.28 133.28 1.28 125.72 0 125.72 0 125.28 1.28 125.28 1.28 117.72 0 117.72 0 117.28 1.28 117.28 1.28 101.72 0 101.72 0 101.28 1.28 101.28 1.28 85.72 0 85.72 0 85.28 1.28 85.28 1.28 69.72 0 69.72 0 0 75 0 ;
    LAYER Via1 ;
      RECT 0 0 75 350 ;
    LAYER Via2 ;
      RECT 0 0 75 350 ;
  END

END gf180mcu_ocd_io__dvss
