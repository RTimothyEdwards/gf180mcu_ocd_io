magic
tech gf180mcuD
magscale 1 10
timestamp 1484609607
<< pwell >>
rect 597 223 1973 3135
<< mvndiff >>
rect 597 3098 685 3135
rect 597 1772 610 3098
rect 656 1772 685 3098
rect 597 1735 685 1772
rect 1885 3098 1973 3135
rect 1885 1772 1914 3098
rect 1960 1772 1973 3098
rect 1885 1735 1973 1772
rect 597 1586 685 1623
rect 597 260 610 1586
rect 656 260 685 1586
rect 597 223 685 260
rect 1885 1586 1973 1623
rect 1885 260 1914 1586
rect 1960 260 1973 1586
rect 1885 223 1973 260
<< mvndiffc >>
rect 610 1772 656 3098
rect 1914 1772 1960 3098
rect 610 260 656 1586
rect 1914 260 1960 1586
<< mvnmoscap >>
rect 685 1735 1885 3135
rect 685 223 1885 1623
<< polysilicon >>
rect 685 3214 1885 3227
rect 685 3168 738 3214
rect 1832 3168 1885 3214
rect 685 3135 1885 3168
rect 685 1702 1885 1735
rect 685 1656 738 1702
rect 1832 1656 1885 1702
rect 685 1623 1885 1656
rect 685 190 1885 223
rect 685 144 738 190
rect 1832 144 1885 190
rect 685 131 1885 144
<< polycontact >>
rect 738 3168 1832 3214
rect 738 1656 1832 1702
rect 738 144 1832 190
<< metal1 >>
rect 310 3285 2260 3485
rect 310 3098 667 3285
rect 727 3214 1843 3225
rect 727 3168 738 3214
rect 1832 3168 1843 3214
rect 727 3161 1088 3168
rect 1140 3161 1220 3168
rect 1272 3161 1352 3168
rect 1404 3161 1843 3168
rect 727 3157 1843 3161
rect 310 1772 610 3098
rect 656 1772 667 3098
rect 310 1586 667 1772
rect 785 1713 1785 3157
rect 1903 3098 2260 3285
rect 1903 1772 1914 3098
rect 1960 1772 2260 3098
rect 727 1702 1843 1713
rect 727 1656 738 1702
rect 1832 1656 1843 1702
rect 727 1645 1843 1656
rect 310 260 610 1586
rect 656 260 667 1586
rect 310 73 667 260
rect 785 201 1785 1645
rect 1903 1586 2260 1772
rect 1903 260 1914 1586
rect 1960 260 2260 1586
rect 727 197 1843 201
rect 727 190 1088 197
rect 1140 190 1220 197
rect 1272 190 1352 197
rect 1404 190 1843 197
rect 727 144 738 190
rect 1832 144 1843 190
rect 727 133 1843 144
rect 1903 73 2260 260
rect 310 -127 2260 73
<< via1 >>
rect 1088 3168 1140 3213
rect 1220 3168 1272 3213
rect 1352 3168 1404 3213
rect 1088 3161 1140 3168
rect 1220 3161 1272 3168
rect 1352 3161 1404 3168
rect 1088 190 1140 197
rect 1220 190 1272 197
rect 1352 190 1404 197
rect 1088 145 1140 190
rect 1220 145 1272 190
rect 1352 145 1404 190
<< metal2 >>
rect 1076 3213 1427 3485
rect 1076 3161 1088 3213
rect 1140 3161 1220 3213
rect 1272 3161 1352 3213
rect 1404 3161 1427 3213
rect 1076 197 1427 3161
rect 1076 145 1088 197
rect 1140 145 1220 197
rect 1272 145 1352 197
rect 1404 145 1427 197
rect 1076 -127 1427 145
<< end >>
