* NGSPICE file created from gf180mcu_ocd_io__fill10.ext - technology: gf180mcuD

.subckt POLY_SUB_FILL_1 a_597_223# a_685_131#
X0 a_685_131# a_597_223# cap_nmos_06v0 c_width=7u c_length=6u
X1 a_685_131# a_597_223# cap_nmos_06v0 c_width=7u c_length=6u
.ends

.subckt GF_NI_FILL10_1 VSS VDD DVSS DVDD
XPOLY_SUB_FILL_1_0[0] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[1] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[2] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[3] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[4] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[5] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[6] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[7] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[8] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[9] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[10] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[11] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[12] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[13] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[14] VSS VDD POLY_SUB_FILL_1
XPOLY_SUB_FILL_1_0[15] VSS VDD POLY_SUB_FILL_1
.ends

.subckt GF_NI_FILL10_0 DVSS DVDD VDD VSS
XGF_NI_FILL10_1_0 VSS VDD DVSS DVDD GF_NI_FILL10_1
.ends

.subckt gf180mcu_ocd_io__fill10 DVSS DVDD VDD VSS
XGF_NI_FILL10_0_0 DVSS DVDD VDD VSS GF_NI_FILL10_0
.ends

