magic
tech gf180mcuD
magscale 1 10
timestamp 1758744525
<< error_s >>
rect 44700 49809 46320 49817
rect 44824 49685 46444 49693
rect 44948 49561 46568 49569
rect 45072 49437 46692 49445
rect 45196 49313 46816 49321
rect 45320 49189 46940 49197
rect 45444 49065 47064 49073
rect 39075 48629 40695 48637
rect 41310 48629 42930 48637
rect 43609 48629 45229 48637
rect 39199 48505 40819 48513
rect 41434 48505 43054 48513
rect 43733 48505 45353 48513
rect 39323 48381 40943 48389
rect 41558 48381 43178 48389
rect 43857 48381 45477 48389
rect 39447 48257 41067 48265
rect 41682 48257 43302 48265
rect 43981 48257 45601 48265
rect 39571 48133 41191 48141
rect 41806 48133 43426 48141
rect 44105 48133 45725 48141
rect 39695 48009 41315 48017
rect 41930 48009 43550 48017
rect 44229 48009 45849 48017
rect 39819 47885 41439 47893
rect 42054 47885 43674 47893
rect 44353 47885 45973 47893
rect 39943 47761 41563 47769
rect 42178 47761 43798 47769
rect 44477 47761 46097 47769
rect 40067 47637 41687 47645
rect 42302 47637 43922 47645
rect 44601 47637 46221 47645
rect 40191 47513 41811 47521
rect 42426 47513 44046 47521
rect 44725 47513 46345 47521
rect 40315 47389 41935 47397
rect 42550 47389 44170 47397
rect 44849 47389 46469 47397
rect 40439 47265 42059 47273
rect 42674 47265 44294 47273
rect 44973 47265 46593 47273
rect 40563 47141 42183 47149
rect 42798 47141 44418 47149
rect 45097 47141 46717 47149
rect 32511 46686 35935 46694
rect 32520 46562 36053 46570
rect 32576 46438 36124 46446
rect 32556 46314 36228 46322
rect 32535 46190 36331 46198
rect 32550 46066 36464 46074
rect 32674 45942 36650 45950
rect 32798 45818 36774 45826
rect 32922 45694 36898 45702
rect 33046 45570 37022 45578
rect 33170 45446 37146 45454
rect 33294 45322 37270 45330
rect 33418 45198 37394 45206
rect 29440 44570 33416 44578
rect 27739 44542 29055 44550
rect 43161 44519 44905 44527
rect 29564 44446 33540 44454
rect 27741 44418 29057 44426
rect 43285 44395 45029 44403
rect 29688 44322 33664 44330
rect 27731 44294 29171 44302
rect 43409 44271 45153 44279
rect 29812 44198 33788 44206
rect 27762 44170 29326 44178
rect 43533 44147 45277 44155
rect 29936 44074 33912 44082
rect 27752 44046 29440 44054
rect 43657 44023 45401 44031
rect 30060 43950 34036 43958
rect 27833 43922 29577 43930
rect 43781 43899 45525 43907
rect 30184 43826 34160 43834
rect 27957 43798 29701 43806
rect 43905 43775 45649 43783
rect 43718 43284 43726 43340
rect 43774 41720 43782 43284
rect 43842 43160 43850 43216
rect 43898 41596 43906 43160
rect 43966 43036 43974 43092
rect 44022 41472 44030 43036
rect 44090 42912 44098 42968
rect 44146 41348 44154 42912
rect 44214 42788 44222 42844
rect 44270 41224 44278 42788
rect 44338 42664 44346 42720
rect 44394 41100 44402 42664
rect 44462 42540 44470 42596
rect 44518 40976 44526 42540
rect 47084 39918 47092 39974
rect 45141 39599 45149 39655
rect 45197 38035 45205 39599
rect 45265 39475 45273 39531
rect 45321 37911 45329 39475
rect 45389 39351 45397 39407
rect 45445 37787 45453 39351
rect 45513 39227 45521 39283
rect 45569 37663 45577 39227
rect 45637 39103 45645 39159
rect 45693 37539 45701 39103
rect 45761 38979 45769 39035
rect 45817 37415 45825 38979
rect 45885 38855 45893 38911
rect 45941 37291 45949 38855
rect 46009 38731 46017 38787
rect 46065 37167 46073 38731
rect 46133 38607 46141 38663
rect 46189 37043 46197 38607
rect 46257 38483 46265 38539
rect 46313 36919 46321 38483
rect 46381 38359 46389 38415
rect 46437 36795 46445 38359
rect 47140 38354 47148 39918
rect 47208 39794 47216 39850
rect 46505 38235 46513 38291
rect 46561 36671 46569 38235
rect 47264 38230 47272 39794
rect 47332 39670 47340 39726
rect 46629 38111 46637 38167
rect 46685 36547 46693 38111
rect 47388 38106 47396 39670
rect 47456 39546 47464 39602
rect 47512 37982 47520 39546
rect 47580 39422 47588 39478
rect 47636 37858 47644 39422
rect 47704 39298 47712 39354
rect 47760 37734 47768 39298
rect 47828 39174 47836 39230
rect 47884 37610 47892 39174
rect 47952 39050 47960 39106
rect 48008 37486 48016 39050
rect 48076 38920 48084 38976
rect 48132 37362 48140 38920
rect 48200 38791 48208 38847
rect 48256 37356 48264 38791
rect 48324 38680 48332 38725
rect 48380 37364 48388 38680
rect 48448 38659 48456 38680
rect 48504 37364 48512 38659
rect 48572 38658 48580 38659
rect 48628 37343 48636 38658
use comp018green_esd_clamp_v5p0_1  comp018green_esd_clamp_v5p0_1_0
timestamp 1758726819
transform 1 0 43564 0 1 51
box -4188 -51 13013 56967
use comp018green_esd_clamp_v5p0_2  comp018green_esd_clamp_v5p0_2_0
timestamp 1758726819
transform 0 1 51 1 0 43565
box -407 -51 13369 47415
use power_via_cor_3  power_via_cor_3_0
timestamp 1758726819
transform 1 0 42556 0 1 508
box 1094 35210 14833 56443
use power_via_cor_5  power_via_cor_5_0
timestamp 1758726819
transform 0 1 508 1 0 42557
box 1068 32 14833 50982
<< end >>
