magic
tech gf180mcuD
magscale 1 10
timestamp 1758750476
<< metal5 >>
rect 14000 70000 17000 71000
rect 17200 70000 20200 71000
rect 20400 70000 23400 71000
rect 23600 70000 25000 71000
rect 25200 70000 26600 71000
rect 26800 70000 29800 71000
rect 30000 70000 33000 71000
rect 33200 70000 36200 71000
rect 36400 70000 39400 71000
rect 39600 70000 41000 71000
rect 41200 70000 42600 71000
rect 42800 70000 45800 71000
rect 46000 70000 49000 71000
rect 49200 70000 50600 71000
rect 50800 70000 52200 71000
rect 52400 70000 53800 71000
rect 54000 70000 55400 71000
rect 55600 70000 57000 71000
rect 57200 70000 58600 71000
rect 58800 70000 60200 71000
rect 60400 70000 61800 71000
rect 62000 70000 63400 71000
rect 63600 70000 65000 71000
rect 65200 70000 66600 71000
rect 66800 70000 68200 71000
rect 68400 70000 69678 71000
rect 70000 68400 71000 69678
rect 70000 66800 71000 68200
rect 70000 65200 71000 66600
rect 70000 63600 71000 65000
rect 70000 62000 71000 63400
rect 70000 60400 71000 61800
rect 70000 58800 71000 60200
rect 70000 57200 71000 58600
rect 70000 55600 71000 57000
rect 70000 54000 71000 55400
rect 70000 52400 71000 53800
rect 70000 50800 71000 52200
rect 70000 49200 71000 50600
rect 70000 46000 71000 49000
rect 70000 42800 71000 45799
rect 70000 41200 71000 42600
rect 70000 39600 71000 41000
rect 70000 36400 71000 39400
rect 70000 33200 71000 36200
rect 70000 30000 71000 33000
rect 70000 26800 71000 29800
rect 70000 25200 71000 26600
rect 70000 23600 71000 25000
rect 70000 20400 71000 23400
rect 70000 17200 71000 20200
rect 70000 14000 71000 17000
use GF_NI_COR_BASE  GF_NI_COR_BASE_0
timestamp 1758750476
transform 1 0 12 0 1 0
box 13436 13361 70889 70890
use POWER_RAIL_COR  POWER_RAIL_COR_0
timestamp 1758726819
transform 1 0 0 0 1 0
box 13097 13097 71000 71000
<< labels >>
rlabel metal3 s 53064 70220 53064 70220 4 DVDD
port 1 nsew
rlabel metal3 s 49849 70219 49849 70219 4 VSS
port 4 nsew
rlabel metal3 s 44292 70220 44292 70220 4 DVDD
port 1 nsew
rlabel metal3 s 41877 70220 41877 70220 4 DVDD
port 1 nsew
rlabel metal3 s 40319 70220 40319 70220 4 DVSS
port 2 nsew
rlabel metal3 s 37671 70220 37671 70220 4 DVDD
port 1 nsew
rlabel metal3 s 34449 70220 34449 70220 4 DVDD
port 1 nsew
rlabel metal3 s 31313 70220 31313 70220 4 DVDD
port 1 nsew
rlabel metal3 s 28097 70220 28097 70220 4 DVDD
port 1 nsew
rlabel metal3 s 64328 70220 64328 70220 4 VSS
port 4 nsew
rlabel metal3 s 62716 70220 62716 70220 4 VDD
port 3 nsew
rlabel metal3 s 57931 70220 57931 70220 4 DVSS
port 2 nsew
rlabel metal3 s 70444 59576 70444 59576 4 DVDD
port 1 nsew
rlabel metal3 s 70444 56376 70444 56376 4 DVDD
port 1 nsew
rlabel metal3 s 70444 54611 70444 54611 4 DVDD
port 1 nsew
rlabel metal3 s 70444 53176 70444 53176 4 DVDD
port 1 nsew
rlabel metal3 s 70444 44321 70444 44321 4 DVDD
port 1 nsew
rlabel metal3 s 70444 41930 70444 41930 4 DVDD
port 1 nsew
rlabel metal3 s 70444 37912 70444 37912 4 DVDD
port 1 nsew
rlabel metal3 s 70444 34676 70444 34676 4 DVDD
port 1 nsew
rlabel metal3 s 70444 31562 70444 31562 4 DVDD
port 1 nsew
rlabel metal3 s 70444 28347 70444 28347 4 DVDD
port 1 nsew
rlabel metal3 s 70444 24237 70444 24237 4 DVDD
port 1 nsew
rlabel metal3 s 70444 64211 70444 64211 4 VSS
port 4 nsew
rlabel metal3 s 70444 69002 70444 69002 4 DVSS
port 2 nsew
rlabel metal3 s 56327 70220 56327 70220 4 DVDD
port 1 nsew
rlabel metal3 s 51498 70220 51498 70220 4 VDD
port 3 nsew
rlabel metal3 s 47523 70220 47523 70220 4 DVSS
port 2 nsew
rlabel metal3 s 70443 62776 70443 62776 4 VDD
port 3 nsew
rlabel metal3 s 70444 67411 70444 67411 4 DVDD
port 1 nsew
rlabel metal3 s 15448 70196 15448 70196 4 DVSS
port 2 nsew
rlabel metal3 s 18634 70150 18634 70150 4 DVSS
port 2 nsew
rlabel metal3 s 21613 70220 21613 70220 4 DVSS
port 2 nsew
rlabel metal3 s 23985 70220 23985 70220 4 DVDD
port 1 nsew
rlabel metal3 s 25800 70220 25800 70220 4 DVSS
port 2 nsew
rlabel metal3 s 59509 70220 59509 70220 4 DVDD
port 1 nsew
rlabel metal3 s 61124 70220 61124 70220 4 DVSS
port 2 nsew
rlabel metal3 s 65891 70220 65891 70220 4 DVSS
port 2 nsew
rlabel metal3 s 70547 49976 70547 49976 4 VSS
port 4 nsew
rlabel metal3 s 70548 51411 70548 51411 4 VDD
port 3 nsew
rlabel metal3 s 67482 70220 67482 70220 4 DVDD
port 1 nsew
rlabel metal3 s 69026 70220 69026 70220 4 DVSS
port 2 nsew
rlabel metal3 s 70375 18874 70375 18874 4 DVSS
port 2 nsew
rlabel metal3 s 70422 15703 70422 15703 4 DVSS
port 2 nsew
rlabel metal3 s 70444 21860 70444 21860 4 DVSS
port 2 nsew
rlabel metal3 s 70444 26053 70444 26053 4 DVSS
port 2 nsew
rlabel metal3 s 70444 40295 70444 40295 4 DVSS
port 2 nsew
rlabel metal3 s 70444 47548 70444 47548 4 DVSS
port 2 nsew
rlabel metal3 s 70444 57811 70444 57811 4 DVSS
port 2 nsew
rlabel metal3 s 70444 61011 70444 61011 4 DVSS
port 2 nsew
rlabel metal3 s 70444 65976 70444 65976 4 DVSS
port 2 nsew
rlabel metal3 s 54690 70220 54690 70220 4 DVDD
port 1 nsew
rlabel metal4 s 69026 70220 69026 70220 4 DVSS
port 2 nsew
rlabel metal4 s 70548 51411 70548 51411 4 VDD
port 3 nsew
rlabel metal4 s 65891 70220 65891 70220 4 DVSS
port 2 nsew
rlabel metal4 s 62716 70220 62716 70220 4 VDD
port 3 nsew
rlabel metal4 s 59509 70220 59509 70220 4 DVDD
port 1 nsew
rlabel metal4 s 56327 70220 56327 70220 4 DVDD
port 1 nsew
rlabel metal4 s 53064 70220 53064 70220 4 DVDD
port 1 nsew
rlabel metal4 s 49849 70219 49849 70219 4 VSS
port 4 nsew
rlabel metal4 s 44292 70220 44292 70220 4 DVDD
port 1 nsew
rlabel metal4 s 40319 70220 40319 70220 4 DVSS
port 2 nsew
rlabel metal4 s 34449 70220 34449 70220 4 DVDD
port 1 nsew
rlabel metal4 s 28097 70220 28097 70220 4 DVDD
port 1 nsew
rlabel metal4 s 23985 70220 23985 70220 4 DVDD
port 1 nsew
rlabel metal4 s 18634 70150 18634 70150 4 DVSS
port 2 nsew
rlabel metal4 s 70444 67411 70444 67411 4 DVDD
port 1 nsew
rlabel metal4 s 70444 59576 70444 59576 4 DVDD
port 1 nsew
rlabel metal4 s 70444 54611 70444 54611 4 DVDD
port 1 nsew
rlabel metal4 s 70444 44321 70444 44321 4 DVDD
port 1 nsew
rlabel metal4 s 70444 37912 70444 37912 4 DVDD
port 1 nsew
rlabel metal4 s 70444 31562 70444 31562 4 DVDD
port 1 nsew
rlabel metal4 s 70444 24237 70444 24237 4 DVDD
port 1 nsew
rlabel metal4 s 70444 69002 70444 69002 4 DVSS
port 2 nsew
rlabel metal4 s 70444 61011 70444 61011 4 DVSS
port 2 nsew
rlabel metal4 s 70444 47548 70444 47548 4 DVSS
port 2 nsew
rlabel metal4 s 70444 26053 70444 26053 4 DVSS
port 2 nsew
rlabel metal4 s 70422 15703 70422 15703 4 DVSS
port 2 nsew
rlabel metal4 s 67482 70220 67482 70220 4 DVDD
port 1 nsew
rlabel metal4 s 70547 49976 70547 49976 4 VSS
port 4 nsew
rlabel metal4 s 64328 70220 64328 70220 4 VSS
port 4 nsew
rlabel metal4 s 61124 70220 61124 70220 4 DVSS
port 2 nsew
rlabel metal4 s 57931 70220 57931 70220 4 DVSS
port 2 nsew
rlabel metal4 s 54690 70220 54690 70220 4 DVDD
port 1 nsew
rlabel metal4 s 51498 70220 51498 70220 4 VDD
port 3 nsew
rlabel metal4 s 47523 70220 47523 70220 4 DVSS
port 2 nsew
rlabel metal4 s 41877 70220 41877 70220 4 DVDD
port 1 nsew
rlabel metal4 s 37671 70220 37671 70220 4 DVDD
port 1 nsew
rlabel metal4 s 31313 70220 31313 70220 4 DVDD
port 1 nsew
rlabel metal4 s 25800 70220 25800 70220 4 DVSS
port 2 nsew
rlabel metal4 s 21613 70220 21613 70220 4 DVSS
port 2 nsew
rlabel metal4 s 15448 70196 15448 70196 4 DVSS
port 2 nsew
rlabel metal4 s 70444 62776 70444 62776 4 VDD
port 3 nsew
rlabel metal4 s 70444 56376 70444 56376 4 DVDD
port 1 nsew
rlabel metal4 s 70444 53176 70444 53176 4 DVDD
port 1 nsew
rlabel metal4 s 70444 41930 70444 41930 4 DVDD
port 1 nsew
rlabel metal4 s 70444 34676 70444 34676 4 DVDD
port 1 nsew
rlabel metal4 s 70444 28347 70444 28347 4 DVDD
port 1 nsew
rlabel metal4 s 70444 64211 70444 64211 4 VSS
port 4 nsew
rlabel metal4 s 70444 65976 70444 65976 4 DVSS
port 2 nsew
rlabel metal4 s 70444 57811 70444 57811 4 DVSS
port 2 nsew
rlabel metal4 s 70444 40295 70444 40295 4 DVSS
port 2 nsew
rlabel metal4 s 70444 21860 70444 21860 4 DVSS
port 2 nsew
rlabel metal4 s 70375 18874 70375 18874 4 DVSS
port 2 nsew
rlabel metal5 s 67482 70220 67482 70220 4 DVDD
port 1 nsew
rlabel metal5 s 69026 70220 69026 70220 4 DVSS
port 2 nsew
rlabel metal5 s 70547 49976 70547 49976 4 VSS
port 4 nsew
rlabel metal5 s 70444 47548 70444 47548 4 DVSS
port 2 nsew
rlabel metal5 s 70444 57811 70444 57811 4 DVSS
port 2 nsew
rlabel metal5 s 70444 61011 70444 61011 4 DVSS
port 2 nsew
rlabel metal5 s 70444 65976 70444 65976 4 DVSS
port 2 nsew
rlabel metal5 s 70444 69002 70444 69002 4 DVSS
port 2 nsew
rlabel metal5 s 70444 64211 70444 64211 4 VSS
port 4 nsew
rlabel metal5 s 70548 51411 70548 51411 4 VDD
port 3 nsew
rlabel metal5 s 70444 44321 70444 44321 4 DVDD
port 1 nsew
rlabel metal5 s 70444 53176 70444 53176 4 DVDD
port 1 nsew
rlabel metal5 s 70444 54611 70444 54611 4 DVDD
port 1 nsew
rlabel metal5 s 70444 56376 70444 56376 4 DVDD
port 1 nsew
rlabel metal5 s 70444 59576 70444 59576 4 DVDD
port 1 nsew
rlabel metal5 s 70444 62776 70444 62776 4 VDD
port 3 nsew
rlabel metal5 s 70444 67411 70444 67411 4 DVDD
port 1 nsew
rlabel metal5 s 44292 70220 44292 70220 4 DVDD
port 1 nsew
rlabel metal5 s 47523 70220 47523 70220 4 DVSS
port 2 nsew
rlabel metal5 s 49849 70219 49849 70219 4 VSS
port 4 nsew
rlabel metal5 s 51498 70220 51498 70220 4 VDD
port 3 nsew
rlabel metal5 s 53064 70220 53064 70220 4 DVDD
port 1 nsew
rlabel metal5 s 54690 70220 54690 70220 4 DVDD
port 1 nsew
rlabel metal5 s 56327 70220 56327 70220 4 DVDD
port 1 nsew
rlabel metal5 s 57931 70220 57931 70220 4 DVSS
port 2 nsew
rlabel metal5 s 59509 70220 59509 70220 4 DVDD
port 1 nsew
rlabel metal5 s 61124 70220 61124 70220 4 DVSS
port 2 nsew
rlabel metal5 s 62716 70220 62716 70220 4 VDD
port 3 nsew
rlabel metal5 s 64328 70220 64328 70220 4 VSS
port 4 nsew
rlabel metal5 s 65891 70220 65891 70220 4 DVSS
port 2 nsew
rlabel metal5 s 67482 70220 67482 70220 4 DVDD
port 1 nsew
rlabel metal5 s 69026 70220 69026 70220 4 DVSS
port 2 nsew
rlabel metal5 s 70547 49976 70547 49976 4 VSS
port 4 nsew
rlabel metal5 s 70444 47548 70444 47548 4 DVSS
port 2 nsew
rlabel metal5 s 70444 57811 70444 57811 4 DVSS
port 2 nsew
rlabel metal5 s 70444 61011 70444 61011 4 DVSS
port 2 nsew
rlabel metal5 s 70444 65976 70444 65976 4 DVSS
port 2 nsew
rlabel metal5 s 70444 69002 70444 69002 4 DVSS
port 2 nsew
rlabel metal5 s 70444 64211 70444 64211 4 VSS
port 4 nsew
rlabel metal5 s 70548 51411 70548 51411 4 VDD
port 3 nsew
rlabel metal5 s 70444 44321 70444 44321 4 DVDD
port 1 nsew
rlabel metal5 s 70444 53176 70444 53176 4 DVDD
port 1 nsew
rlabel metal5 s 70444 54611 70444 54611 4 DVDD
port 1 nsew
rlabel metal5 s 70444 56376 70444 56376 4 DVDD
port 1 nsew
rlabel metal5 s 70444 59576 70444 59576 4 DVDD
port 1 nsew
rlabel metal5 s 70444 62776 70444 62776 4 VDD
port 3 nsew
rlabel metal5 s 70444 67411 70444 67411 4 DVDD
port 1 nsew
rlabel metal5 s 44292 70220 44292 70220 4 DVDD
port 1 nsew
rlabel metal5 s 47523 70220 47523 70220 4 DVSS
port 2 nsew
rlabel metal5 s 49849 70219 49849 70219 4 VSS
port 4 nsew
rlabel metal5 s 51498 70220 51498 70220 4 VDD
port 3 nsew
rlabel metal5 s 53064 70220 53064 70220 4 DVDD
port 1 nsew
rlabel metal5 s 54690 70220 54690 70220 4 DVDD
port 1 nsew
rlabel metal5 s 56327 70220 56327 70220 4 DVDD
port 1 nsew
rlabel metal5 s 57931 70220 57931 70220 4 DVSS
port 2 nsew
rlabel metal5 s 59509 70220 59509 70220 4 DVDD
port 1 nsew
rlabel metal5 s 61124 70220 61124 70220 4 DVSS
port 2 nsew
rlabel metal5 s 62716 70220 62716 70220 4 VDD
port 3 nsew
rlabel metal5 s 64328 70220 64328 70220 4 VSS
port 4 nsew
rlabel metal5 s 65891 70220 65891 70220 4 DVSS
port 2 nsew
rlabel metal5 s 70547 49976 70547 49976 4 VSS
port 4 nsew
rlabel metal5 s 70548 51411 70548 51411 4 VDD
port 3 nsew
rlabel metal5 s 67482 70220 67482 70220 4 DVDD
port 1 nsew
rlabel metal5 s 69026 70220 69026 70220 4 DVSS
port 2 nsew
rlabel metal5 s 70444 47548 70444 47548 4 DVSS
port 2 nsew
rlabel metal5 s 70444 57811 70444 57811 4 DVSS
port 2 nsew
rlabel metal5 s 70444 61011 70444 61011 4 DVSS
port 2 nsew
rlabel metal5 s 70444 65976 70444 65976 4 DVSS
port 2 nsew
rlabel metal5 s 70444 69002 70444 69002 4 DVSS
port 2 nsew
rlabel metal5 s 70444 44321 70444 44321 4 DVDD
port 1 nsew
rlabel metal5 s 70444 53176 70444 53176 4 DVDD
port 1 nsew
rlabel metal5 s 70444 54611 70444 54611 4 DVDD
port 1 nsew
rlabel metal5 s 70444 56376 70444 56376 4 DVDD
port 1 nsew
rlabel metal5 s 70444 59576 70444 59576 4 DVDD
port 1 nsew
rlabel metal5 s 70444 62776 70444 62776 4 VDD
port 3 nsew
rlabel metal5 s 70444 67411 70444 67411 4 DVDD
port 1 nsew
rlabel metal5 s 44292 70220 44292 70220 4 DVDD
port 1 nsew
rlabel metal5 s 47523 70220 47523 70220 4 DVSS
port 2 nsew
rlabel metal5 s 49849 70219 49849 70219 4 VSS
port 4 nsew
rlabel metal5 s 51498 70220 51498 70220 4 VDD
port 3 nsew
rlabel metal5 s 53064 70220 53064 70220 4 DVDD
port 1 nsew
rlabel metal5 s 54690 70220 54690 70220 4 DVDD
port 1 nsew
rlabel metal5 s 56327 70220 56327 70220 4 DVDD
port 1 nsew
rlabel metal5 s 57931 70220 57931 70220 4 DVSS
port 2 nsew
rlabel metal5 s 59509 70220 59509 70220 4 DVDD
port 1 nsew
rlabel metal5 s 61124 70220 61124 70220 4 DVSS
port 2 nsew
rlabel metal5 s 62716 70220 62716 70220 4 VDD
port 3 nsew
rlabel metal5 s 64328 70220 64328 70220 4 VSS
port 4 nsew
rlabel metal5 s 65891 70220 65891 70220 4 DVSS
port 2 nsew
rlabel metal5 s 40319 70220 40319 70220 4 DVSS
port 2 nsew
rlabel metal5 s 41877 70220 41877 70220 4 DVDD
port 1 nsew
rlabel metal5 s 37671 70220 37671 70220 4 DVDD
port 1 nsew
rlabel metal5 s 40319 70220 40319 70220 4 DVSS
port 2 nsew
rlabel metal5 s 41877 70220 41877 70220 4 DVDD
port 1 nsew
rlabel metal5 s 15448 70196 15448 70196 4 DVSS
port 2 nsew
rlabel metal5 s 18634 70150 18634 70150 4 DVSS
port 2 nsew
rlabel metal5 s 21613 70220 21613 70220 4 DVSS
port 2 nsew
rlabel metal5 s 23985 70220 23985 70220 4 DVDD
port 1 nsew
rlabel metal5 s 15448 70196 15448 70196 4 DVSS
port 2 nsew
rlabel metal5 s 18634 70150 18634 70150 4 DVSS
port 2 nsew
rlabel metal5 s 21613 70220 21613 70220 4 DVSS
port 2 nsew
rlabel metal5 s 23985 70220 23985 70220 4 DVDD
port 1 nsew
rlabel metal5 s 25800 70220 25800 70220 4 DVSS
port 2 nsew
rlabel metal5 s 28097 70220 28097 70220 4 DVDD
port 1 nsew
rlabel metal5 s 31313 70220 31313 70220 4 DVDD
port 1 nsew
rlabel metal5 s 34449 70220 34449 70220 4 DVDD
port 1 nsew
rlabel metal5 s 37671 70220 37671 70220 4 DVDD
port 1 nsew
rlabel metal5 s 40319 70220 40319 70220 4 DVSS
port 2 nsew
rlabel metal5 s 41877 70220 41877 70220 4 DVDD
port 1 nsew
rlabel metal5 s 25800 70220 25800 70220 4 DVSS
port 2 nsew
rlabel metal5 s 28097 70220 28097 70220 4 DVDD
port 1 nsew
rlabel metal5 s 31313 70220 31313 70220 4 DVDD
port 1 nsew
rlabel metal5 s 34449 70220 34449 70220 4 DVDD
port 1 nsew
rlabel metal5 s 15448 70196 15448 70196 4 DVSS
port 2 nsew
rlabel metal5 s 18634 70150 18634 70150 4 DVSS
port 2 nsew
rlabel metal5 s 21613 70220 21613 70220 4 DVSS
port 2 nsew
rlabel metal5 s 23985 70220 23985 70220 4 DVDD
port 1 nsew
rlabel metal5 s 25800 70220 25800 70220 4 DVSS
port 2 nsew
rlabel metal5 s 28097 70220 28097 70220 4 DVDD
port 1 nsew
rlabel metal5 s 31313 70220 31313 70220 4 DVDD
port 1 nsew
rlabel metal5 s 34449 70220 34449 70220 4 DVDD
port 1 nsew
rlabel metal5 s 37671 70220 37671 70220 4 DVDD
port 1 nsew
rlabel metal5 s 70444 37912 70444 37912 4 DVDD
port 1 nsew
rlabel metal5 s 70444 41930 70444 41930 4 DVDD
port 1 nsew
rlabel metal5 s 70444 31562 70444 31562 4 DVDD
port 1 nsew
rlabel metal5 s 70444 34676 70444 34676 4 DVDD
port 1 nsew
rlabel metal5 s 70444 37912 70444 37912 4 DVDD
port 1 nsew
rlabel metal5 s 70444 41930 70444 41930 4 DVDD
port 1 nsew
rlabel metal5 s 70444 34676 70444 34676 4 DVDD
port 1 nsew
rlabel metal5 s 70444 37912 70444 37912 4 DVDD
port 1 nsew
rlabel metal5 s 70444 41930 70444 41930 4 DVDD
port 1 nsew
rlabel metal5 s 70375 18874 70375 18874 4 DVSS
port 2 nsew
rlabel metal5 s 70422 15703 70422 15703 4 DVSS
port 2 nsew
rlabel metal5 s 70444 21860 70444 21860 4 DVSS
port 2 nsew
rlabel metal5 s 70444 21860 70444 21860 4 DVSS
port 2 nsew
rlabel metal5 s 70444 26053 70444 26053 4 DVSS
port 2 nsew
rlabel metal5 s 70444 40295 70444 40295 4 DVSS
port 2 nsew
rlabel metal5 s 70444 26053 70444 26053 4 DVSS
port 2 nsew
rlabel metal5 s 70444 40295 70444 40295 4 DVSS
port 2 nsew
rlabel metal5 s 70422 15703 70422 15703 4 DVSS
port 2 nsew
rlabel metal5 s 70375 18874 70375 18874 4 DVSS
port 2 nsew
rlabel metal5 s 70375 18874 70375 18874 4 DVSS
port 2 nsew
rlabel metal5 s 70422 15703 70422 15703 4 DVSS
port 2 nsew
rlabel metal5 s 70444 21860 70444 21860 4 DVSS
port 2 nsew
rlabel metal5 s 70444 26053 70444 26053 4 DVSS
port 2 nsew
rlabel metal5 s 70444 40295 70444 40295 4 DVSS
port 2 nsew
rlabel metal5 s 70444 24237 70444 24237 4 DVDD
port 1 nsew
rlabel metal5 s 70444 28347 70444 28347 4 DVDD
port 1 nsew
rlabel metal5 s 70444 31562 70444 31562 4 DVDD
port 1 nsew
rlabel metal5 s 70444 24237 70444 24237 4 DVDD
port 1 nsew
rlabel metal5 s 70444 28347 70444 28347 4 DVDD
port 1 nsew
rlabel metal5 s 70444 24237 70444 24237 4 DVDD
port 1 nsew
rlabel metal5 s 70444 28347 70444 28347 4 DVDD
port 1 nsew
rlabel metal5 s 70444 31562 70444 31562 4 DVDD
port 1 nsew
rlabel metal5 s 70444 34676 70444 34676 4 DVDD
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 71000 71000
<< end >>
