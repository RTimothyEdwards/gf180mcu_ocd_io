# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_ocd_io__brk5
    CLASS PAD ;
  ORIGIN 0 0 ;
    FOREIGN gf180mcu_ocd_io__brk5 0 0 ;
  SIZE 5 BY 350 ;
  SYMMETRY X Y R90 ;
  SITE GF_IO_Site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 4 246 5 253 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 4 318 5 325 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 318 1 325 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 246 1 253 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 0 0 5 350 ;
    LAYER Metal2 ;
      RECT 0 0 5 350 ;
    LAYER Metal3 ;
      POLYGON 5 69.72 3.72 69.72 3.72 85.28 5 85.28 5 85.72 3.72 85.72 3.72 101.28 5 101.28 5 101.72 3.72 101.72 3.72 117.28 5 117.28 5 117.72 3.72 117.72 3.72 125.28 5 125.28 5 125.72 3.72 125.72 3.72 133.28 5 133.28 5 133.72 3.72 133.72 3.72 149.28 5 149.28 5 149.72 3.72 149.72 3.72 165.28 5 165.28 5 165.72 3.72 165.72 3.72 181.28 5 181.28 5 181.72 3.72 181.72 3.72 197.28 5 197.28 5 197.72 3.72 197.72 3.72 205.28 5 205.28 5 205.72 3.72 205.72 3.72 213.28 5 213.28 5 213.72 3.72 213.72 3.72 229.28 5 229.28 5 229.72 3.72 229.72 3.72 245.28 5 245.28 5 245.72 3.72 245.72 3.72 253.28 5 253.28 5 253.72 3.72 253.72 3.72 261.28 5 261.28 5 261.72 3.72 261.72 3.72 269.28 5 269.28 5 269.72 3.72 269.72 3.72 277.28 5 277.28 5 277.72 3.72 277.72 3.72 285.28 5 285.28 5 285.72 3.72 285.72 3.72 293.28 5 293.28 5 293.72 3.72 293.72 3.72 301.28 5 301.28 5 301.72 3.72 301.72 3.72 309.28 5 309.28 5 309.72 3.72 309.72 3.72 317.28 5 317.28 5 317.72 3.72 317.72 3.72 325.28 5 325.28 5 325.72 3.72 325.72 3.72 333.28 5 333.28 5 333.72 3.72 333.72 3.72 341.28 5 341.28 5 341.72 3.72 341.72 3.72 348.67 5 348.67 5 350 0 350 0 348.67 1.28 348.67 1.28 341.72 0 341.72 0 341.28 1.28 341.28 1.28 333.72 0 333.72 0 333.28 1.28 333.28 1.28 325.72 0 325.72 0 325.28 1.28 325.28 1.28 317.72 0 317.72 0 317.28 1.28 317.28 1.28 309.72 0 309.72 0 309.28 1.28 309.28 1.28 301.72 0 301.72 0 301.28 1.28 301.28 1.28 293.72 0 293.72 0 293.28 1.28 293.28 1.28 285.72 0 285.72 0 285.28 1.28 285.28 1.28 277.72 0 277.72 0 277.28 1.28 277.28 1.28 269.72 0 269.72 0 269.28 1.28 269.28 1.28 261.72 0 261.72 0 261.28 1.28 261.28 1.28 253.72 0 253.72 0 253.28 1.28 253.28 1.28 245.72 0 245.72 0 245.28 1.28 245.28 1.28 229.72 0 229.72 0 229.28 1.28 229.28 1.28 213.72 0 213.72 0 213.28 1.28 213.28 1.28 205.72 0 205.72 0 205.28 1.28 205.28 1.28 197.72 0 197.72 0 197.28 1.28 197.28 1.28 181.72 0 181.72 0 181.28 1.28 181.28 1.28 165.72 0 165.72 0 165.28 1.28 165.28 1.28 149.72 0 149.72 0 149.28 1.28 149.28 1.28 133.72 0 133.72 0 133.28 1.28 133.28 1.28 125.72 0 125.72 0 125.28 1.28 125.28 1.28 117.72 0 117.72 0 117.28 1.28 117.28 1.28 101.72 0 101.72 0 101.28 1.28 101.28 1.28 85.72 0 85.72 0 85.28 1.28 85.28 1.28 69.72 0 69.72 0 0 5 0 ;
    LAYER Via1 ;
      RECT 0 0 5 350 ;
    LAYER Via2 ;
      RECT 0 0 5 350 ;
  END

END gf180mcu_ocd_io__brk5
