magic
tech gf180mcuD
magscale 1 5
timestamp 1758724778
use pmos_6p0_esd  pmos_6p0_esd_0
timestamp 1758724778
transform 1 0 0 0 1 0
box 0 6 598 6126
<< end >>
