VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_ocd_io__bi_24t
  CLASS PAD INOUT ;
  FOREIGN gf180mcu_ocd_io__bi_24t ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 350.000 ;
  SYMMETRY X Y R90 ;
  SITE GF_IO_Site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.504000 ;
    ANTENNADIFFAREA 1.000000 ;
    PORT
      LAYER Metal2 ;
        RECT 69.400 266.830 69.780 349.760 ;
    END
  END A
  PIN CS
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.504000 ;
    ANTENNADIFFAREA 1.000000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.360 328.305 3.740 349.760 ;
    END
  END CS
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 0.000 118.000 5.000 125.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 134.000 5.000 149.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 150.000 5.000 165.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 166.000 5.000 181.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 182.000 5.000 197.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 206.000 5.000 213.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 214.000 5.000 229.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 262.000 5.000 269.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 270.000 5.000 277.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 278.000 5.000 285.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 294.000 5.000 301.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 334.000 5.000 341.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 70.000 118.000 75.000 125.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 70.000 134.000 75.000 149.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 70.000 150.000 75.000 165.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 70.000 166.000 75.000 181.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 70.000 182.000 75.000 197.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 70.000 206.000 75.000 213.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 70.000 214.000 75.000 229.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 70.000 262.000 75.000 269.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 70.000 270.000 75.000 277.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 70.000 278.000 75.000 285.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 70.000 294.000 75.000 301.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 70.000 334.000 75.000 341.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 0.000 70.000 5.000 85.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 86.000 5.000 101.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 102.000 5.000 117.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 126.000 5.000 133.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 198.000 5.000 205.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 230.000 5.000 245.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 286.000 5.000 293.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 302.000 5.000 309.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 326.000 5.000 333.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 342.000 5.000 348.390 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 70.000 70.000 75.000 85.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 70.000 86.000 75.000 101.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 70.000 102.000 75.000 117.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 70.000 126.000 75.000 133.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 70.000 198.000 75.000 205.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 70.000 230.000 75.000 245.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 70.000 286.000 75.000 293.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 70.000 302.000 75.000 309.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 70.000 326.000 75.000 333.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 70.000 342.000 75.000 348.390 ;
    END
  END DVSS
  PIN IE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.504000 ;
    ANTENNADIFFAREA 1.000000 ;
    PORT
      LAYER Metal2 ;
        RECT 11.385 334.680 11.765 349.760 ;
    END
  END IE
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.016000 ;
    ANTENNADIFFAREA 7.776000 ;
    PORT
      LAYER Metal2 ;
        RECT 70.130 283.205 70.510 349.760 ;
    END
  END OE
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 335.279999 ;
    PORT
      LAYER Metal4 ;
        RECT 7.500 2.000 67.500 62.000 ;
    END
  END PAD
  PIN PD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.512000 ;
    ANTENNADIFFAREA 1.000000 ;
    PORT
      LAYER Metal2 ;
        RECT 10.330 329.860 10.710 349.760 ;
    END
  END PD
  PIN PU
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.008000 ;
    ANTENNADIFFAREA 1.795000 ;
    PORT
      LAYER Metal2 ;
        RECT 5.965 330.180 6.345 349.760 ;
    END
  END PU
  PIN SL
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.504000 ;
    ANTENNADIFFAREA 1.000000 ;
    PORT
      LAYER Metal2 ;
        RECT 68.670 266.100 69.050 349.760 ;
    END
  END SL
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 0.000 254.000 5.000 261.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 310.000 5.000 317.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 70.000 254.000 75.000 261.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 70.000 310.000 75.000 317.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 0.000 246.000 5.000 253.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 318.000 5.000 325.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 70.000 246.000 75.000 253.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 70.000 318.000 75.000 325.000 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.240000 ;
    PORT
      LAYER Metal2 ;
        RECT 70.860 319.660 71.240 349.760 ;
    END
  END Y
  OBS
      LAYER Nwell ;
        RECT 1.820 67.400 73.180 346.295 ;
      LAYER Metal1 ;
        RECT -0.160 65.450 75.160 349.785 ;
      LAYER Metal2 ;
        RECT 0.000 328.005 3.060 348.135 ;
        RECT 4.040 329.880 5.665 348.135 ;
        RECT 6.645 329.880 10.030 348.135 ;
        RECT 4.040 329.560 10.030 329.880 ;
        RECT 11.010 334.380 11.085 348.135 ;
        RECT 12.065 334.380 68.370 348.135 ;
        RECT 11.010 329.560 68.370 334.380 ;
        RECT 4.040 328.005 68.370 329.560 ;
        RECT 0.000 265.800 68.370 328.005 ;
        RECT 71.540 319.360 75.000 348.135 ;
        RECT 70.810 282.905 75.000 319.360 ;
        RECT 70.080 266.530 75.000 282.905 ;
        RECT 69.350 265.800 75.000 266.530 ;
        RECT 0.000 0.000 75.000 265.800 ;
      LAYER Metal3 ;
        RECT 0.000 0.000 75.000 348.390 ;
      LAYER Metal4 ;
        RECT 5.600 69.400 69.400 348.390 ;
        RECT 3.500 62.600 71.500 69.400 ;
        RECT 3.500 1.400 6.900 62.600 ;
        RECT 68.100 1.400 71.500 62.600 ;
        RECT 3.500 0.000 71.500 1.400 ;
  END
END gf180mcu_ocd_io__bi_24t
END LIBRARY

