magic
tech gf180mcuD
magscale 1 10
timestamp 1586916644
<< metal3 >>
rect 151 69637 14853 69647
rect 151 69581 161 69637
rect 217 69581 303 69637
rect 359 69581 445 69637
rect 501 69581 587 69637
rect 643 69581 729 69637
rect 785 69581 871 69637
rect 927 69581 1013 69637
rect 1069 69581 1155 69637
rect 1211 69581 1297 69637
rect 1353 69581 1439 69637
rect 1495 69581 1581 69637
rect 1637 69581 1723 69637
rect 1779 69581 1865 69637
rect 1921 69581 2007 69637
rect 2063 69581 2149 69637
rect 2205 69581 2291 69637
rect 2347 69581 2433 69637
rect 2489 69581 2575 69637
rect 2631 69581 2717 69637
rect 2773 69581 2859 69637
rect 2915 69581 3001 69637
rect 3057 69581 3143 69637
rect 3199 69581 3285 69637
rect 3341 69581 3427 69637
rect 3483 69581 3569 69637
rect 3625 69581 3711 69637
rect 3767 69581 3853 69637
rect 3909 69581 3995 69637
rect 4051 69581 4137 69637
rect 4193 69581 4279 69637
rect 4335 69581 4421 69637
rect 4477 69581 4563 69637
rect 4619 69581 4705 69637
rect 4761 69581 4847 69637
rect 4903 69581 4989 69637
rect 5045 69581 5131 69637
rect 5187 69581 5273 69637
rect 5329 69581 5415 69637
rect 5471 69581 5557 69637
rect 5613 69581 5699 69637
rect 5755 69581 5841 69637
rect 5897 69581 5983 69637
rect 6039 69581 6125 69637
rect 6181 69581 6267 69637
rect 6323 69581 6409 69637
rect 6465 69581 6551 69637
rect 6607 69581 6693 69637
rect 6749 69581 6835 69637
rect 6891 69581 6977 69637
rect 7033 69581 7119 69637
rect 7175 69581 7261 69637
rect 7317 69581 7403 69637
rect 7459 69581 7545 69637
rect 7601 69581 7687 69637
rect 7743 69581 7829 69637
rect 7885 69581 7971 69637
rect 8027 69581 8113 69637
rect 8169 69581 8255 69637
rect 8311 69581 8397 69637
rect 8453 69581 8539 69637
rect 8595 69581 8681 69637
rect 8737 69581 8823 69637
rect 8879 69581 8965 69637
rect 9021 69581 9107 69637
rect 9163 69581 9249 69637
rect 9305 69581 9391 69637
rect 9447 69581 9533 69637
rect 9589 69581 9675 69637
rect 9731 69581 9817 69637
rect 9873 69581 9959 69637
rect 10015 69581 10101 69637
rect 10157 69581 10243 69637
rect 10299 69581 10385 69637
rect 10441 69581 10527 69637
rect 10583 69581 10669 69637
rect 10725 69581 10811 69637
rect 10867 69581 10953 69637
rect 11009 69581 11095 69637
rect 11151 69581 11237 69637
rect 11293 69581 11379 69637
rect 11435 69581 11521 69637
rect 11577 69581 11663 69637
rect 11719 69581 11805 69637
rect 11861 69581 11947 69637
rect 12003 69581 12089 69637
rect 12145 69581 12231 69637
rect 12287 69581 12373 69637
rect 12429 69581 12515 69637
rect 12571 69581 12657 69637
rect 12713 69581 12799 69637
rect 12855 69581 12941 69637
rect 12997 69581 13083 69637
rect 13139 69581 13225 69637
rect 13281 69581 13367 69637
rect 13423 69581 13509 69637
rect 13565 69581 13651 69637
rect 13707 69581 13793 69637
rect 13849 69581 13935 69637
rect 13991 69581 14077 69637
rect 14133 69581 14219 69637
rect 14275 69581 14361 69637
rect 14417 69581 14503 69637
rect 14559 69581 14645 69637
rect 14701 69581 14787 69637
rect 14843 69581 14853 69637
rect 151 69495 14853 69581
rect 151 69439 161 69495
rect 217 69439 303 69495
rect 359 69439 445 69495
rect 501 69439 587 69495
rect 643 69439 729 69495
rect 785 69439 871 69495
rect 927 69439 1013 69495
rect 1069 69439 1155 69495
rect 1211 69439 1297 69495
rect 1353 69439 1439 69495
rect 1495 69439 1581 69495
rect 1637 69439 1723 69495
rect 1779 69439 1865 69495
rect 1921 69439 2007 69495
rect 2063 69439 2149 69495
rect 2205 69439 2291 69495
rect 2347 69439 2433 69495
rect 2489 69439 2575 69495
rect 2631 69439 2717 69495
rect 2773 69439 2859 69495
rect 2915 69439 3001 69495
rect 3057 69439 3143 69495
rect 3199 69439 3285 69495
rect 3341 69439 3427 69495
rect 3483 69439 3569 69495
rect 3625 69439 3711 69495
rect 3767 69439 3853 69495
rect 3909 69439 3995 69495
rect 4051 69439 4137 69495
rect 4193 69439 4279 69495
rect 4335 69439 4421 69495
rect 4477 69439 4563 69495
rect 4619 69439 4705 69495
rect 4761 69439 4847 69495
rect 4903 69439 4989 69495
rect 5045 69439 5131 69495
rect 5187 69439 5273 69495
rect 5329 69439 5415 69495
rect 5471 69439 5557 69495
rect 5613 69439 5699 69495
rect 5755 69439 5841 69495
rect 5897 69439 5983 69495
rect 6039 69439 6125 69495
rect 6181 69439 6267 69495
rect 6323 69439 6409 69495
rect 6465 69439 6551 69495
rect 6607 69439 6693 69495
rect 6749 69439 6835 69495
rect 6891 69439 6977 69495
rect 7033 69439 7119 69495
rect 7175 69439 7261 69495
rect 7317 69439 7403 69495
rect 7459 69439 7545 69495
rect 7601 69439 7687 69495
rect 7743 69439 7829 69495
rect 7885 69439 7971 69495
rect 8027 69439 8113 69495
rect 8169 69439 8255 69495
rect 8311 69439 8397 69495
rect 8453 69439 8539 69495
rect 8595 69439 8681 69495
rect 8737 69439 8823 69495
rect 8879 69439 8965 69495
rect 9021 69439 9107 69495
rect 9163 69439 9249 69495
rect 9305 69439 9391 69495
rect 9447 69439 9533 69495
rect 9589 69439 9675 69495
rect 9731 69439 9817 69495
rect 9873 69439 9959 69495
rect 10015 69439 10101 69495
rect 10157 69439 10243 69495
rect 10299 69439 10385 69495
rect 10441 69439 10527 69495
rect 10583 69439 10669 69495
rect 10725 69439 10811 69495
rect 10867 69439 10953 69495
rect 11009 69439 11095 69495
rect 11151 69439 11237 69495
rect 11293 69439 11379 69495
rect 11435 69439 11521 69495
rect 11577 69439 11663 69495
rect 11719 69439 11805 69495
rect 11861 69439 11947 69495
rect 12003 69439 12089 69495
rect 12145 69439 12231 69495
rect 12287 69439 12373 69495
rect 12429 69439 12515 69495
rect 12571 69439 12657 69495
rect 12713 69439 12799 69495
rect 12855 69439 12941 69495
rect 12997 69439 13083 69495
rect 13139 69439 13225 69495
rect 13281 69439 13367 69495
rect 13423 69439 13509 69495
rect 13565 69439 13651 69495
rect 13707 69439 13793 69495
rect 13849 69439 13935 69495
rect 13991 69439 14077 69495
rect 14133 69439 14219 69495
rect 14275 69439 14361 69495
rect 14417 69439 14503 69495
rect 14559 69439 14645 69495
rect 14701 69439 14787 69495
rect 14843 69439 14853 69495
rect 151 69353 14853 69439
rect 151 69297 161 69353
rect 217 69297 303 69353
rect 359 69297 445 69353
rect 501 69297 587 69353
rect 643 69297 729 69353
rect 785 69297 871 69353
rect 927 69297 1013 69353
rect 1069 69297 1155 69353
rect 1211 69297 1297 69353
rect 1353 69297 1439 69353
rect 1495 69297 1581 69353
rect 1637 69297 1723 69353
rect 1779 69297 1865 69353
rect 1921 69297 2007 69353
rect 2063 69297 2149 69353
rect 2205 69297 2291 69353
rect 2347 69297 2433 69353
rect 2489 69297 2575 69353
rect 2631 69297 2717 69353
rect 2773 69297 2859 69353
rect 2915 69297 3001 69353
rect 3057 69297 3143 69353
rect 3199 69297 3285 69353
rect 3341 69297 3427 69353
rect 3483 69297 3569 69353
rect 3625 69297 3711 69353
rect 3767 69297 3853 69353
rect 3909 69297 3995 69353
rect 4051 69297 4137 69353
rect 4193 69297 4279 69353
rect 4335 69297 4421 69353
rect 4477 69297 4563 69353
rect 4619 69297 4705 69353
rect 4761 69297 4847 69353
rect 4903 69297 4989 69353
rect 5045 69297 5131 69353
rect 5187 69297 5273 69353
rect 5329 69297 5415 69353
rect 5471 69297 5557 69353
rect 5613 69297 5699 69353
rect 5755 69297 5841 69353
rect 5897 69297 5983 69353
rect 6039 69297 6125 69353
rect 6181 69297 6267 69353
rect 6323 69297 6409 69353
rect 6465 69297 6551 69353
rect 6607 69297 6693 69353
rect 6749 69297 6835 69353
rect 6891 69297 6977 69353
rect 7033 69297 7119 69353
rect 7175 69297 7261 69353
rect 7317 69297 7403 69353
rect 7459 69297 7545 69353
rect 7601 69297 7687 69353
rect 7743 69297 7829 69353
rect 7885 69297 7971 69353
rect 8027 69297 8113 69353
rect 8169 69297 8255 69353
rect 8311 69297 8397 69353
rect 8453 69297 8539 69353
rect 8595 69297 8681 69353
rect 8737 69297 8823 69353
rect 8879 69297 8965 69353
rect 9021 69297 9107 69353
rect 9163 69297 9249 69353
rect 9305 69297 9391 69353
rect 9447 69297 9533 69353
rect 9589 69297 9675 69353
rect 9731 69297 9817 69353
rect 9873 69297 9959 69353
rect 10015 69297 10101 69353
rect 10157 69297 10243 69353
rect 10299 69297 10385 69353
rect 10441 69297 10527 69353
rect 10583 69297 10669 69353
rect 10725 69297 10811 69353
rect 10867 69297 10953 69353
rect 11009 69297 11095 69353
rect 11151 69297 11237 69353
rect 11293 69297 11379 69353
rect 11435 69297 11521 69353
rect 11577 69297 11663 69353
rect 11719 69297 11805 69353
rect 11861 69297 11947 69353
rect 12003 69297 12089 69353
rect 12145 69297 12231 69353
rect 12287 69297 12373 69353
rect 12429 69297 12515 69353
rect 12571 69297 12657 69353
rect 12713 69297 12799 69353
rect 12855 69297 12941 69353
rect 12997 69297 13083 69353
rect 13139 69297 13225 69353
rect 13281 69297 13367 69353
rect 13423 69297 13509 69353
rect 13565 69297 13651 69353
rect 13707 69297 13793 69353
rect 13849 69297 13935 69353
rect 13991 69297 14077 69353
rect 14133 69297 14219 69353
rect 14275 69297 14361 69353
rect 14417 69297 14503 69353
rect 14559 69297 14645 69353
rect 14701 69297 14787 69353
rect 14843 69297 14853 69353
rect 151 69211 14853 69297
rect 151 69155 161 69211
rect 217 69155 303 69211
rect 359 69155 445 69211
rect 501 69155 587 69211
rect 643 69155 729 69211
rect 785 69155 871 69211
rect 927 69155 1013 69211
rect 1069 69155 1155 69211
rect 1211 69155 1297 69211
rect 1353 69155 1439 69211
rect 1495 69155 1581 69211
rect 1637 69155 1723 69211
rect 1779 69155 1865 69211
rect 1921 69155 2007 69211
rect 2063 69155 2149 69211
rect 2205 69155 2291 69211
rect 2347 69155 2433 69211
rect 2489 69155 2575 69211
rect 2631 69155 2717 69211
rect 2773 69155 2859 69211
rect 2915 69155 3001 69211
rect 3057 69155 3143 69211
rect 3199 69155 3285 69211
rect 3341 69155 3427 69211
rect 3483 69155 3569 69211
rect 3625 69155 3711 69211
rect 3767 69155 3853 69211
rect 3909 69155 3995 69211
rect 4051 69155 4137 69211
rect 4193 69155 4279 69211
rect 4335 69155 4421 69211
rect 4477 69155 4563 69211
rect 4619 69155 4705 69211
rect 4761 69155 4847 69211
rect 4903 69155 4989 69211
rect 5045 69155 5131 69211
rect 5187 69155 5273 69211
rect 5329 69155 5415 69211
rect 5471 69155 5557 69211
rect 5613 69155 5699 69211
rect 5755 69155 5841 69211
rect 5897 69155 5983 69211
rect 6039 69155 6125 69211
rect 6181 69155 6267 69211
rect 6323 69155 6409 69211
rect 6465 69155 6551 69211
rect 6607 69155 6693 69211
rect 6749 69155 6835 69211
rect 6891 69155 6977 69211
rect 7033 69155 7119 69211
rect 7175 69155 7261 69211
rect 7317 69155 7403 69211
rect 7459 69155 7545 69211
rect 7601 69155 7687 69211
rect 7743 69155 7829 69211
rect 7885 69155 7971 69211
rect 8027 69155 8113 69211
rect 8169 69155 8255 69211
rect 8311 69155 8397 69211
rect 8453 69155 8539 69211
rect 8595 69155 8681 69211
rect 8737 69155 8823 69211
rect 8879 69155 8965 69211
rect 9021 69155 9107 69211
rect 9163 69155 9249 69211
rect 9305 69155 9391 69211
rect 9447 69155 9533 69211
rect 9589 69155 9675 69211
rect 9731 69155 9817 69211
rect 9873 69155 9959 69211
rect 10015 69155 10101 69211
rect 10157 69155 10243 69211
rect 10299 69155 10385 69211
rect 10441 69155 10527 69211
rect 10583 69155 10669 69211
rect 10725 69155 10811 69211
rect 10867 69155 10953 69211
rect 11009 69155 11095 69211
rect 11151 69155 11237 69211
rect 11293 69155 11379 69211
rect 11435 69155 11521 69211
rect 11577 69155 11663 69211
rect 11719 69155 11805 69211
rect 11861 69155 11947 69211
rect 12003 69155 12089 69211
rect 12145 69155 12231 69211
rect 12287 69155 12373 69211
rect 12429 69155 12515 69211
rect 12571 69155 12657 69211
rect 12713 69155 12799 69211
rect 12855 69155 12941 69211
rect 12997 69155 13083 69211
rect 13139 69155 13225 69211
rect 13281 69155 13367 69211
rect 13423 69155 13509 69211
rect 13565 69155 13651 69211
rect 13707 69155 13793 69211
rect 13849 69155 13935 69211
rect 13991 69155 14077 69211
rect 14133 69155 14219 69211
rect 14275 69155 14361 69211
rect 14417 69155 14503 69211
rect 14559 69155 14645 69211
rect 14701 69155 14787 69211
rect 14843 69155 14853 69211
rect 151 69069 14853 69155
rect 151 69013 161 69069
rect 217 69013 303 69069
rect 359 69013 445 69069
rect 501 69013 587 69069
rect 643 69013 729 69069
rect 785 69013 871 69069
rect 927 69013 1013 69069
rect 1069 69013 1155 69069
rect 1211 69013 1297 69069
rect 1353 69013 1439 69069
rect 1495 69013 1581 69069
rect 1637 69013 1723 69069
rect 1779 69013 1865 69069
rect 1921 69013 2007 69069
rect 2063 69013 2149 69069
rect 2205 69013 2291 69069
rect 2347 69013 2433 69069
rect 2489 69013 2575 69069
rect 2631 69013 2717 69069
rect 2773 69013 2859 69069
rect 2915 69013 3001 69069
rect 3057 69013 3143 69069
rect 3199 69013 3285 69069
rect 3341 69013 3427 69069
rect 3483 69013 3569 69069
rect 3625 69013 3711 69069
rect 3767 69013 3853 69069
rect 3909 69013 3995 69069
rect 4051 69013 4137 69069
rect 4193 69013 4279 69069
rect 4335 69013 4421 69069
rect 4477 69013 4563 69069
rect 4619 69013 4705 69069
rect 4761 69013 4847 69069
rect 4903 69013 4989 69069
rect 5045 69013 5131 69069
rect 5187 69013 5273 69069
rect 5329 69013 5415 69069
rect 5471 69013 5557 69069
rect 5613 69013 5699 69069
rect 5755 69013 5841 69069
rect 5897 69013 5983 69069
rect 6039 69013 6125 69069
rect 6181 69013 6267 69069
rect 6323 69013 6409 69069
rect 6465 69013 6551 69069
rect 6607 69013 6693 69069
rect 6749 69013 6835 69069
rect 6891 69013 6977 69069
rect 7033 69013 7119 69069
rect 7175 69013 7261 69069
rect 7317 69013 7403 69069
rect 7459 69013 7545 69069
rect 7601 69013 7687 69069
rect 7743 69013 7829 69069
rect 7885 69013 7971 69069
rect 8027 69013 8113 69069
rect 8169 69013 8255 69069
rect 8311 69013 8397 69069
rect 8453 69013 8539 69069
rect 8595 69013 8681 69069
rect 8737 69013 8823 69069
rect 8879 69013 8965 69069
rect 9021 69013 9107 69069
rect 9163 69013 9249 69069
rect 9305 69013 9391 69069
rect 9447 69013 9533 69069
rect 9589 69013 9675 69069
rect 9731 69013 9817 69069
rect 9873 69013 9959 69069
rect 10015 69013 10101 69069
rect 10157 69013 10243 69069
rect 10299 69013 10385 69069
rect 10441 69013 10527 69069
rect 10583 69013 10669 69069
rect 10725 69013 10811 69069
rect 10867 69013 10953 69069
rect 11009 69013 11095 69069
rect 11151 69013 11237 69069
rect 11293 69013 11379 69069
rect 11435 69013 11521 69069
rect 11577 69013 11663 69069
rect 11719 69013 11805 69069
rect 11861 69013 11947 69069
rect 12003 69013 12089 69069
rect 12145 69013 12231 69069
rect 12287 69013 12373 69069
rect 12429 69013 12515 69069
rect 12571 69013 12657 69069
rect 12713 69013 12799 69069
rect 12855 69013 12941 69069
rect 12997 69013 13083 69069
rect 13139 69013 13225 69069
rect 13281 69013 13367 69069
rect 13423 69013 13509 69069
rect 13565 69013 13651 69069
rect 13707 69013 13793 69069
rect 13849 69013 13935 69069
rect 13991 69013 14077 69069
rect 14133 69013 14219 69069
rect 14275 69013 14361 69069
rect 14417 69013 14503 69069
rect 14559 69013 14645 69069
rect 14701 69013 14787 69069
rect 14843 69013 14853 69069
rect 151 68927 14853 69013
rect 151 68871 161 68927
rect 217 68871 303 68927
rect 359 68871 445 68927
rect 501 68871 587 68927
rect 643 68871 729 68927
rect 785 68871 871 68927
rect 927 68871 1013 68927
rect 1069 68871 1155 68927
rect 1211 68871 1297 68927
rect 1353 68871 1439 68927
rect 1495 68871 1581 68927
rect 1637 68871 1723 68927
rect 1779 68871 1865 68927
rect 1921 68871 2007 68927
rect 2063 68871 2149 68927
rect 2205 68871 2291 68927
rect 2347 68871 2433 68927
rect 2489 68871 2575 68927
rect 2631 68871 2717 68927
rect 2773 68871 2859 68927
rect 2915 68871 3001 68927
rect 3057 68871 3143 68927
rect 3199 68871 3285 68927
rect 3341 68871 3427 68927
rect 3483 68871 3569 68927
rect 3625 68871 3711 68927
rect 3767 68871 3853 68927
rect 3909 68871 3995 68927
rect 4051 68871 4137 68927
rect 4193 68871 4279 68927
rect 4335 68871 4421 68927
rect 4477 68871 4563 68927
rect 4619 68871 4705 68927
rect 4761 68871 4847 68927
rect 4903 68871 4989 68927
rect 5045 68871 5131 68927
rect 5187 68871 5273 68927
rect 5329 68871 5415 68927
rect 5471 68871 5557 68927
rect 5613 68871 5699 68927
rect 5755 68871 5841 68927
rect 5897 68871 5983 68927
rect 6039 68871 6125 68927
rect 6181 68871 6267 68927
rect 6323 68871 6409 68927
rect 6465 68871 6551 68927
rect 6607 68871 6693 68927
rect 6749 68871 6835 68927
rect 6891 68871 6977 68927
rect 7033 68871 7119 68927
rect 7175 68871 7261 68927
rect 7317 68871 7403 68927
rect 7459 68871 7545 68927
rect 7601 68871 7687 68927
rect 7743 68871 7829 68927
rect 7885 68871 7971 68927
rect 8027 68871 8113 68927
rect 8169 68871 8255 68927
rect 8311 68871 8397 68927
rect 8453 68871 8539 68927
rect 8595 68871 8681 68927
rect 8737 68871 8823 68927
rect 8879 68871 8965 68927
rect 9021 68871 9107 68927
rect 9163 68871 9249 68927
rect 9305 68871 9391 68927
rect 9447 68871 9533 68927
rect 9589 68871 9675 68927
rect 9731 68871 9817 68927
rect 9873 68871 9959 68927
rect 10015 68871 10101 68927
rect 10157 68871 10243 68927
rect 10299 68871 10385 68927
rect 10441 68871 10527 68927
rect 10583 68871 10669 68927
rect 10725 68871 10811 68927
rect 10867 68871 10953 68927
rect 11009 68871 11095 68927
rect 11151 68871 11237 68927
rect 11293 68871 11379 68927
rect 11435 68871 11521 68927
rect 11577 68871 11663 68927
rect 11719 68871 11805 68927
rect 11861 68871 11947 68927
rect 12003 68871 12089 68927
rect 12145 68871 12231 68927
rect 12287 68871 12373 68927
rect 12429 68871 12515 68927
rect 12571 68871 12657 68927
rect 12713 68871 12799 68927
rect 12855 68871 12941 68927
rect 12997 68871 13083 68927
rect 13139 68871 13225 68927
rect 13281 68871 13367 68927
rect 13423 68871 13509 68927
rect 13565 68871 13651 68927
rect 13707 68871 13793 68927
rect 13849 68871 13935 68927
rect 13991 68871 14077 68927
rect 14133 68871 14219 68927
rect 14275 68871 14361 68927
rect 14417 68871 14503 68927
rect 14559 68871 14645 68927
rect 14701 68871 14787 68927
rect 14843 68871 14853 68927
rect 151 68785 14853 68871
rect 151 68729 161 68785
rect 217 68729 303 68785
rect 359 68729 445 68785
rect 501 68729 587 68785
rect 643 68729 729 68785
rect 785 68729 871 68785
rect 927 68729 1013 68785
rect 1069 68729 1155 68785
rect 1211 68729 1297 68785
rect 1353 68729 1439 68785
rect 1495 68729 1581 68785
rect 1637 68729 1723 68785
rect 1779 68729 1865 68785
rect 1921 68729 2007 68785
rect 2063 68729 2149 68785
rect 2205 68729 2291 68785
rect 2347 68729 2433 68785
rect 2489 68729 2575 68785
rect 2631 68729 2717 68785
rect 2773 68729 2859 68785
rect 2915 68729 3001 68785
rect 3057 68729 3143 68785
rect 3199 68729 3285 68785
rect 3341 68729 3427 68785
rect 3483 68729 3569 68785
rect 3625 68729 3711 68785
rect 3767 68729 3853 68785
rect 3909 68729 3995 68785
rect 4051 68729 4137 68785
rect 4193 68729 4279 68785
rect 4335 68729 4421 68785
rect 4477 68729 4563 68785
rect 4619 68729 4705 68785
rect 4761 68729 4847 68785
rect 4903 68729 4989 68785
rect 5045 68729 5131 68785
rect 5187 68729 5273 68785
rect 5329 68729 5415 68785
rect 5471 68729 5557 68785
rect 5613 68729 5699 68785
rect 5755 68729 5841 68785
rect 5897 68729 5983 68785
rect 6039 68729 6125 68785
rect 6181 68729 6267 68785
rect 6323 68729 6409 68785
rect 6465 68729 6551 68785
rect 6607 68729 6693 68785
rect 6749 68729 6835 68785
rect 6891 68729 6977 68785
rect 7033 68729 7119 68785
rect 7175 68729 7261 68785
rect 7317 68729 7403 68785
rect 7459 68729 7545 68785
rect 7601 68729 7687 68785
rect 7743 68729 7829 68785
rect 7885 68729 7971 68785
rect 8027 68729 8113 68785
rect 8169 68729 8255 68785
rect 8311 68729 8397 68785
rect 8453 68729 8539 68785
rect 8595 68729 8681 68785
rect 8737 68729 8823 68785
rect 8879 68729 8965 68785
rect 9021 68729 9107 68785
rect 9163 68729 9249 68785
rect 9305 68729 9391 68785
rect 9447 68729 9533 68785
rect 9589 68729 9675 68785
rect 9731 68729 9817 68785
rect 9873 68729 9959 68785
rect 10015 68729 10101 68785
rect 10157 68729 10243 68785
rect 10299 68729 10385 68785
rect 10441 68729 10527 68785
rect 10583 68729 10669 68785
rect 10725 68729 10811 68785
rect 10867 68729 10953 68785
rect 11009 68729 11095 68785
rect 11151 68729 11237 68785
rect 11293 68729 11379 68785
rect 11435 68729 11521 68785
rect 11577 68729 11663 68785
rect 11719 68729 11805 68785
rect 11861 68729 11947 68785
rect 12003 68729 12089 68785
rect 12145 68729 12231 68785
rect 12287 68729 12373 68785
rect 12429 68729 12515 68785
rect 12571 68729 12657 68785
rect 12713 68729 12799 68785
rect 12855 68729 12941 68785
rect 12997 68729 13083 68785
rect 13139 68729 13225 68785
rect 13281 68729 13367 68785
rect 13423 68729 13509 68785
rect 13565 68729 13651 68785
rect 13707 68729 13793 68785
rect 13849 68729 13935 68785
rect 13991 68729 14077 68785
rect 14133 68729 14219 68785
rect 14275 68729 14361 68785
rect 14417 68729 14503 68785
rect 14559 68729 14645 68785
rect 14701 68729 14787 68785
rect 14843 68729 14853 68785
rect 151 68643 14853 68729
rect 151 68587 161 68643
rect 217 68587 303 68643
rect 359 68587 445 68643
rect 501 68587 587 68643
rect 643 68587 729 68643
rect 785 68587 871 68643
rect 927 68587 1013 68643
rect 1069 68587 1155 68643
rect 1211 68587 1297 68643
rect 1353 68587 1439 68643
rect 1495 68587 1581 68643
rect 1637 68587 1723 68643
rect 1779 68587 1865 68643
rect 1921 68587 2007 68643
rect 2063 68587 2149 68643
rect 2205 68587 2291 68643
rect 2347 68587 2433 68643
rect 2489 68587 2575 68643
rect 2631 68587 2717 68643
rect 2773 68587 2859 68643
rect 2915 68587 3001 68643
rect 3057 68587 3143 68643
rect 3199 68587 3285 68643
rect 3341 68587 3427 68643
rect 3483 68587 3569 68643
rect 3625 68587 3711 68643
rect 3767 68587 3853 68643
rect 3909 68587 3995 68643
rect 4051 68587 4137 68643
rect 4193 68587 4279 68643
rect 4335 68587 4421 68643
rect 4477 68587 4563 68643
rect 4619 68587 4705 68643
rect 4761 68587 4847 68643
rect 4903 68587 4989 68643
rect 5045 68587 5131 68643
rect 5187 68587 5273 68643
rect 5329 68587 5415 68643
rect 5471 68587 5557 68643
rect 5613 68587 5699 68643
rect 5755 68587 5841 68643
rect 5897 68587 5983 68643
rect 6039 68587 6125 68643
rect 6181 68587 6267 68643
rect 6323 68587 6409 68643
rect 6465 68587 6551 68643
rect 6607 68587 6693 68643
rect 6749 68587 6835 68643
rect 6891 68587 6977 68643
rect 7033 68587 7119 68643
rect 7175 68587 7261 68643
rect 7317 68587 7403 68643
rect 7459 68587 7545 68643
rect 7601 68587 7687 68643
rect 7743 68587 7829 68643
rect 7885 68587 7971 68643
rect 8027 68587 8113 68643
rect 8169 68587 8255 68643
rect 8311 68587 8397 68643
rect 8453 68587 8539 68643
rect 8595 68587 8681 68643
rect 8737 68587 8823 68643
rect 8879 68587 8965 68643
rect 9021 68587 9107 68643
rect 9163 68587 9249 68643
rect 9305 68587 9391 68643
rect 9447 68587 9533 68643
rect 9589 68587 9675 68643
rect 9731 68587 9817 68643
rect 9873 68587 9959 68643
rect 10015 68587 10101 68643
rect 10157 68587 10243 68643
rect 10299 68587 10385 68643
rect 10441 68587 10527 68643
rect 10583 68587 10669 68643
rect 10725 68587 10811 68643
rect 10867 68587 10953 68643
rect 11009 68587 11095 68643
rect 11151 68587 11237 68643
rect 11293 68587 11379 68643
rect 11435 68587 11521 68643
rect 11577 68587 11663 68643
rect 11719 68587 11805 68643
rect 11861 68587 11947 68643
rect 12003 68587 12089 68643
rect 12145 68587 12231 68643
rect 12287 68587 12373 68643
rect 12429 68587 12515 68643
rect 12571 68587 12657 68643
rect 12713 68587 12799 68643
rect 12855 68587 12941 68643
rect 12997 68587 13083 68643
rect 13139 68587 13225 68643
rect 13281 68587 13367 68643
rect 13423 68587 13509 68643
rect 13565 68587 13651 68643
rect 13707 68587 13793 68643
rect 13849 68587 13935 68643
rect 13991 68587 14077 68643
rect 14133 68587 14219 68643
rect 14275 68587 14361 68643
rect 14417 68587 14503 68643
rect 14559 68587 14645 68643
rect 14701 68587 14787 68643
rect 14843 68587 14853 68643
rect 151 68501 14853 68587
rect 151 68445 161 68501
rect 217 68445 303 68501
rect 359 68445 445 68501
rect 501 68445 587 68501
rect 643 68445 729 68501
rect 785 68445 871 68501
rect 927 68445 1013 68501
rect 1069 68445 1155 68501
rect 1211 68445 1297 68501
rect 1353 68445 1439 68501
rect 1495 68445 1581 68501
rect 1637 68445 1723 68501
rect 1779 68445 1865 68501
rect 1921 68445 2007 68501
rect 2063 68445 2149 68501
rect 2205 68445 2291 68501
rect 2347 68445 2433 68501
rect 2489 68445 2575 68501
rect 2631 68445 2717 68501
rect 2773 68445 2859 68501
rect 2915 68445 3001 68501
rect 3057 68445 3143 68501
rect 3199 68445 3285 68501
rect 3341 68445 3427 68501
rect 3483 68445 3569 68501
rect 3625 68445 3711 68501
rect 3767 68445 3853 68501
rect 3909 68445 3995 68501
rect 4051 68445 4137 68501
rect 4193 68445 4279 68501
rect 4335 68445 4421 68501
rect 4477 68445 4563 68501
rect 4619 68445 4705 68501
rect 4761 68445 4847 68501
rect 4903 68445 4989 68501
rect 5045 68445 5131 68501
rect 5187 68445 5273 68501
rect 5329 68445 5415 68501
rect 5471 68445 5557 68501
rect 5613 68445 5699 68501
rect 5755 68445 5841 68501
rect 5897 68445 5983 68501
rect 6039 68445 6125 68501
rect 6181 68445 6267 68501
rect 6323 68445 6409 68501
rect 6465 68445 6551 68501
rect 6607 68445 6693 68501
rect 6749 68445 6835 68501
rect 6891 68445 6977 68501
rect 7033 68445 7119 68501
rect 7175 68445 7261 68501
rect 7317 68445 7403 68501
rect 7459 68445 7545 68501
rect 7601 68445 7687 68501
rect 7743 68445 7829 68501
rect 7885 68445 7971 68501
rect 8027 68445 8113 68501
rect 8169 68445 8255 68501
rect 8311 68445 8397 68501
rect 8453 68445 8539 68501
rect 8595 68445 8681 68501
rect 8737 68445 8823 68501
rect 8879 68445 8965 68501
rect 9021 68445 9107 68501
rect 9163 68445 9249 68501
rect 9305 68445 9391 68501
rect 9447 68445 9533 68501
rect 9589 68445 9675 68501
rect 9731 68445 9817 68501
rect 9873 68445 9959 68501
rect 10015 68445 10101 68501
rect 10157 68445 10243 68501
rect 10299 68445 10385 68501
rect 10441 68445 10527 68501
rect 10583 68445 10669 68501
rect 10725 68445 10811 68501
rect 10867 68445 10953 68501
rect 11009 68445 11095 68501
rect 11151 68445 11237 68501
rect 11293 68445 11379 68501
rect 11435 68445 11521 68501
rect 11577 68445 11663 68501
rect 11719 68445 11805 68501
rect 11861 68445 11947 68501
rect 12003 68445 12089 68501
rect 12145 68445 12231 68501
rect 12287 68445 12373 68501
rect 12429 68445 12515 68501
rect 12571 68445 12657 68501
rect 12713 68445 12799 68501
rect 12855 68445 12941 68501
rect 12997 68445 13083 68501
rect 13139 68445 13225 68501
rect 13281 68445 13367 68501
rect 13423 68445 13509 68501
rect 13565 68445 13651 68501
rect 13707 68445 13793 68501
rect 13849 68445 13935 68501
rect 13991 68445 14077 68501
rect 14133 68445 14219 68501
rect 14275 68445 14361 68501
rect 14417 68445 14503 68501
rect 14559 68445 14645 68501
rect 14701 68445 14787 68501
rect 14843 68445 14853 68501
rect 151 68435 14853 68445
rect 151 68171 14853 68181
rect 151 68115 161 68171
rect 217 68115 303 68171
rect 359 68115 445 68171
rect 501 68115 587 68171
rect 643 68115 729 68171
rect 785 68115 871 68171
rect 927 68115 1013 68171
rect 1069 68115 1155 68171
rect 1211 68115 1297 68171
rect 1353 68115 1439 68171
rect 1495 68115 1581 68171
rect 1637 68115 1723 68171
rect 1779 68115 1865 68171
rect 1921 68115 2007 68171
rect 2063 68115 2149 68171
rect 2205 68115 2291 68171
rect 2347 68115 2433 68171
rect 2489 68115 2575 68171
rect 2631 68115 2717 68171
rect 2773 68115 2859 68171
rect 2915 68115 3001 68171
rect 3057 68115 3143 68171
rect 3199 68115 3285 68171
rect 3341 68115 3427 68171
rect 3483 68115 3569 68171
rect 3625 68115 3711 68171
rect 3767 68115 3853 68171
rect 3909 68115 3995 68171
rect 4051 68115 4137 68171
rect 4193 68115 4279 68171
rect 4335 68115 4421 68171
rect 4477 68115 4563 68171
rect 4619 68115 4705 68171
rect 4761 68115 4847 68171
rect 4903 68115 4989 68171
rect 5045 68115 5131 68171
rect 5187 68115 5273 68171
rect 5329 68115 5415 68171
rect 5471 68115 5557 68171
rect 5613 68115 5699 68171
rect 5755 68115 5841 68171
rect 5897 68115 5983 68171
rect 6039 68115 6125 68171
rect 6181 68115 6267 68171
rect 6323 68115 6409 68171
rect 6465 68115 6551 68171
rect 6607 68115 6693 68171
rect 6749 68115 6835 68171
rect 6891 68115 6977 68171
rect 7033 68115 7119 68171
rect 7175 68115 7261 68171
rect 7317 68115 7403 68171
rect 7459 68115 7545 68171
rect 7601 68115 7687 68171
rect 7743 68115 7829 68171
rect 7885 68115 7971 68171
rect 8027 68115 8113 68171
rect 8169 68115 8255 68171
rect 8311 68115 8397 68171
rect 8453 68115 8539 68171
rect 8595 68115 8681 68171
rect 8737 68115 8823 68171
rect 8879 68115 8965 68171
rect 9021 68115 9107 68171
rect 9163 68115 9249 68171
rect 9305 68115 9391 68171
rect 9447 68115 9533 68171
rect 9589 68115 9675 68171
rect 9731 68115 9817 68171
rect 9873 68115 9959 68171
rect 10015 68115 10101 68171
rect 10157 68115 10243 68171
rect 10299 68115 10385 68171
rect 10441 68115 10527 68171
rect 10583 68115 10669 68171
rect 10725 68115 10811 68171
rect 10867 68115 10953 68171
rect 11009 68115 11095 68171
rect 11151 68115 11237 68171
rect 11293 68115 11379 68171
rect 11435 68115 11521 68171
rect 11577 68115 11663 68171
rect 11719 68115 11805 68171
rect 11861 68115 11947 68171
rect 12003 68115 12089 68171
rect 12145 68115 12231 68171
rect 12287 68115 12373 68171
rect 12429 68115 12515 68171
rect 12571 68115 12657 68171
rect 12713 68115 12799 68171
rect 12855 68115 12941 68171
rect 12997 68115 13083 68171
rect 13139 68115 13225 68171
rect 13281 68115 13367 68171
rect 13423 68115 13509 68171
rect 13565 68115 13651 68171
rect 13707 68115 13793 68171
rect 13849 68115 13935 68171
rect 13991 68115 14077 68171
rect 14133 68115 14219 68171
rect 14275 68115 14361 68171
rect 14417 68115 14503 68171
rect 14559 68115 14645 68171
rect 14701 68115 14787 68171
rect 14843 68115 14853 68171
rect 151 68029 14853 68115
rect 151 67973 161 68029
rect 217 67973 303 68029
rect 359 67973 445 68029
rect 501 67973 587 68029
rect 643 67973 729 68029
rect 785 67973 871 68029
rect 927 67973 1013 68029
rect 1069 67973 1155 68029
rect 1211 67973 1297 68029
rect 1353 67973 1439 68029
rect 1495 67973 1581 68029
rect 1637 67973 1723 68029
rect 1779 67973 1865 68029
rect 1921 67973 2007 68029
rect 2063 67973 2149 68029
rect 2205 67973 2291 68029
rect 2347 67973 2433 68029
rect 2489 67973 2575 68029
rect 2631 67973 2717 68029
rect 2773 67973 2859 68029
rect 2915 67973 3001 68029
rect 3057 67973 3143 68029
rect 3199 67973 3285 68029
rect 3341 67973 3427 68029
rect 3483 67973 3569 68029
rect 3625 67973 3711 68029
rect 3767 67973 3853 68029
rect 3909 67973 3995 68029
rect 4051 67973 4137 68029
rect 4193 67973 4279 68029
rect 4335 67973 4421 68029
rect 4477 67973 4563 68029
rect 4619 67973 4705 68029
rect 4761 67973 4847 68029
rect 4903 67973 4989 68029
rect 5045 67973 5131 68029
rect 5187 67973 5273 68029
rect 5329 67973 5415 68029
rect 5471 67973 5557 68029
rect 5613 67973 5699 68029
rect 5755 67973 5841 68029
rect 5897 67973 5983 68029
rect 6039 67973 6125 68029
rect 6181 67973 6267 68029
rect 6323 67973 6409 68029
rect 6465 67973 6551 68029
rect 6607 67973 6693 68029
rect 6749 67973 6835 68029
rect 6891 67973 6977 68029
rect 7033 67973 7119 68029
rect 7175 67973 7261 68029
rect 7317 67973 7403 68029
rect 7459 67973 7545 68029
rect 7601 67973 7687 68029
rect 7743 67973 7829 68029
rect 7885 67973 7971 68029
rect 8027 67973 8113 68029
rect 8169 67973 8255 68029
rect 8311 67973 8397 68029
rect 8453 67973 8539 68029
rect 8595 67973 8681 68029
rect 8737 67973 8823 68029
rect 8879 67973 8965 68029
rect 9021 67973 9107 68029
rect 9163 67973 9249 68029
rect 9305 67973 9391 68029
rect 9447 67973 9533 68029
rect 9589 67973 9675 68029
rect 9731 67973 9817 68029
rect 9873 67973 9959 68029
rect 10015 67973 10101 68029
rect 10157 67973 10243 68029
rect 10299 67973 10385 68029
rect 10441 67973 10527 68029
rect 10583 67973 10669 68029
rect 10725 67973 10811 68029
rect 10867 67973 10953 68029
rect 11009 67973 11095 68029
rect 11151 67973 11237 68029
rect 11293 67973 11379 68029
rect 11435 67973 11521 68029
rect 11577 67973 11663 68029
rect 11719 67973 11805 68029
rect 11861 67973 11947 68029
rect 12003 67973 12089 68029
rect 12145 67973 12231 68029
rect 12287 67973 12373 68029
rect 12429 67973 12515 68029
rect 12571 67973 12657 68029
rect 12713 67973 12799 68029
rect 12855 67973 12941 68029
rect 12997 67973 13083 68029
rect 13139 67973 13225 68029
rect 13281 67973 13367 68029
rect 13423 67973 13509 68029
rect 13565 67973 13651 68029
rect 13707 67973 13793 68029
rect 13849 67973 13935 68029
rect 13991 67973 14077 68029
rect 14133 67973 14219 68029
rect 14275 67973 14361 68029
rect 14417 67973 14503 68029
rect 14559 67973 14645 68029
rect 14701 67973 14787 68029
rect 14843 67973 14853 68029
rect 151 67887 14853 67973
rect 151 67831 161 67887
rect 217 67831 303 67887
rect 359 67831 445 67887
rect 501 67831 587 67887
rect 643 67831 729 67887
rect 785 67831 871 67887
rect 927 67831 1013 67887
rect 1069 67831 1155 67887
rect 1211 67831 1297 67887
rect 1353 67831 1439 67887
rect 1495 67831 1581 67887
rect 1637 67831 1723 67887
rect 1779 67831 1865 67887
rect 1921 67831 2007 67887
rect 2063 67831 2149 67887
rect 2205 67831 2291 67887
rect 2347 67831 2433 67887
rect 2489 67831 2575 67887
rect 2631 67831 2717 67887
rect 2773 67831 2859 67887
rect 2915 67831 3001 67887
rect 3057 67831 3143 67887
rect 3199 67831 3285 67887
rect 3341 67831 3427 67887
rect 3483 67831 3569 67887
rect 3625 67831 3711 67887
rect 3767 67831 3853 67887
rect 3909 67831 3995 67887
rect 4051 67831 4137 67887
rect 4193 67831 4279 67887
rect 4335 67831 4421 67887
rect 4477 67831 4563 67887
rect 4619 67831 4705 67887
rect 4761 67831 4847 67887
rect 4903 67831 4989 67887
rect 5045 67831 5131 67887
rect 5187 67831 5273 67887
rect 5329 67831 5415 67887
rect 5471 67831 5557 67887
rect 5613 67831 5699 67887
rect 5755 67831 5841 67887
rect 5897 67831 5983 67887
rect 6039 67831 6125 67887
rect 6181 67831 6267 67887
rect 6323 67831 6409 67887
rect 6465 67831 6551 67887
rect 6607 67831 6693 67887
rect 6749 67831 6835 67887
rect 6891 67831 6977 67887
rect 7033 67831 7119 67887
rect 7175 67831 7261 67887
rect 7317 67831 7403 67887
rect 7459 67831 7545 67887
rect 7601 67831 7687 67887
rect 7743 67831 7829 67887
rect 7885 67831 7971 67887
rect 8027 67831 8113 67887
rect 8169 67831 8255 67887
rect 8311 67831 8397 67887
rect 8453 67831 8539 67887
rect 8595 67831 8681 67887
rect 8737 67831 8823 67887
rect 8879 67831 8965 67887
rect 9021 67831 9107 67887
rect 9163 67831 9249 67887
rect 9305 67831 9391 67887
rect 9447 67831 9533 67887
rect 9589 67831 9675 67887
rect 9731 67831 9817 67887
rect 9873 67831 9959 67887
rect 10015 67831 10101 67887
rect 10157 67831 10243 67887
rect 10299 67831 10385 67887
rect 10441 67831 10527 67887
rect 10583 67831 10669 67887
rect 10725 67831 10811 67887
rect 10867 67831 10953 67887
rect 11009 67831 11095 67887
rect 11151 67831 11237 67887
rect 11293 67831 11379 67887
rect 11435 67831 11521 67887
rect 11577 67831 11663 67887
rect 11719 67831 11805 67887
rect 11861 67831 11947 67887
rect 12003 67831 12089 67887
rect 12145 67831 12231 67887
rect 12287 67831 12373 67887
rect 12429 67831 12515 67887
rect 12571 67831 12657 67887
rect 12713 67831 12799 67887
rect 12855 67831 12941 67887
rect 12997 67831 13083 67887
rect 13139 67831 13225 67887
rect 13281 67831 13367 67887
rect 13423 67831 13509 67887
rect 13565 67831 13651 67887
rect 13707 67831 13793 67887
rect 13849 67831 13935 67887
rect 13991 67831 14077 67887
rect 14133 67831 14219 67887
rect 14275 67831 14361 67887
rect 14417 67831 14503 67887
rect 14559 67831 14645 67887
rect 14701 67831 14787 67887
rect 14843 67831 14853 67887
rect 151 67745 14853 67831
rect 151 67689 161 67745
rect 217 67689 303 67745
rect 359 67689 445 67745
rect 501 67689 587 67745
rect 643 67689 729 67745
rect 785 67689 871 67745
rect 927 67689 1013 67745
rect 1069 67689 1155 67745
rect 1211 67689 1297 67745
rect 1353 67689 1439 67745
rect 1495 67689 1581 67745
rect 1637 67689 1723 67745
rect 1779 67689 1865 67745
rect 1921 67689 2007 67745
rect 2063 67689 2149 67745
rect 2205 67689 2291 67745
rect 2347 67689 2433 67745
rect 2489 67689 2575 67745
rect 2631 67689 2717 67745
rect 2773 67689 2859 67745
rect 2915 67689 3001 67745
rect 3057 67689 3143 67745
rect 3199 67689 3285 67745
rect 3341 67689 3427 67745
rect 3483 67689 3569 67745
rect 3625 67689 3711 67745
rect 3767 67689 3853 67745
rect 3909 67689 3995 67745
rect 4051 67689 4137 67745
rect 4193 67689 4279 67745
rect 4335 67689 4421 67745
rect 4477 67689 4563 67745
rect 4619 67689 4705 67745
rect 4761 67689 4847 67745
rect 4903 67689 4989 67745
rect 5045 67689 5131 67745
rect 5187 67689 5273 67745
rect 5329 67689 5415 67745
rect 5471 67689 5557 67745
rect 5613 67689 5699 67745
rect 5755 67689 5841 67745
rect 5897 67689 5983 67745
rect 6039 67689 6125 67745
rect 6181 67689 6267 67745
rect 6323 67689 6409 67745
rect 6465 67689 6551 67745
rect 6607 67689 6693 67745
rect 6749 67689 6835 67745
rect 6891 67689 6977 67745
rect 7033 67689 7119 67745
rect 7175 67689 7261 67745
rect 7317 67689 7403 67745
rect 7459 67689 7545 67745
rect 7601 67689 7687 67745
rect 7743 67689 7829 67745
rect 7885 67689 7971 67745
rect 8027 67689 8113 67745
rect 8169 67689 8255 67745
rect 8311 67689 8397 67745
rect 8453 67689 8539 67745
rect 8595 67689 8681 67745
rect 8737 67689 8823 67745
rect 8879 67689 8965 67745
rect 9021 67689 9107 67745
rect 9163 67689 9249 67745
rect 9305 67689 9391 67745
rect 9447 67689 9533 67745
rect 9589 67689 9675 67745
rect 9731 67689 9817 67745
rect 9873 67689 9959 67745
rect 10015 67689 10101 67745
rect 10157 67689 10243 67745
rect 10299 67689 10385 67745
rect 10441 67689 10527 67745
rect 10583 67689 10669 67745
rect 10725 67689 10811 67745
rect 10867 67689 10953 67745
rect 11009 67689 11095 67745
rect 11151 67689 11237 67745
rect 11293 67689 11379 67745
rect 11435 67689 11521 67745
rect 11577 67689 11663 67745
rect 11719 67689 11805 67745
rect 11861 67689 11947 67745
rect 12003 67689 12089 67745
rect 12145 67689 12231 67745
rect 12287 67689 12373 67745
rect 12429 67689 12515 67745
rect 12571 67689 12657 67745
rect 12713 67689 12799 67745
rect 12855 67689 12941 67745
rect 12997 67689 13083 67745
rect 13139 67689 13225 67745
rect 13281 67689 13367 67745
rect 13423 67689 13509 67745
rect 13565 67689 13651 67745
rect 13707 67689 13793 67745
rect 13849 67689 13935 67745
rect 13991 67689 14077 67745
rect 14133 67689 14219 67745
rect 14275 67689 14361 67745
rect 14417 67689 14503 67745
rect 14559 67689 14645 67745
rect 14701 67689 14787 67745
rect 14843 67689 14853 67745
rect 151 67603 14853 67689
rect 151 67547 161 67603
rect 217 67547 303 67603
rect 359 67547 445 67603
rect 501 67547 587 67603
rect 643 67547 729 67603
rect 785 67547 871 67603
rect 927 67547 1013 67603
rect 1069 67547 1155 67603
rect 1211 67547 1297 67603
rect 1353 67547 1439 67603
rect 1495 67547 1581 67603
rect 1637 67547 1723 67603
rect 1779 67547 1865 67603
rect 1921 67547 2007 67603
rect 2063 67547 2149 67603
rect 2205 67547 2291 67603
rect 2347 67547 2433 67603
rect 2489 67547 2575 67603
rect 2631 67547 2717 67603
rect 2773 67547 2859 67603
rect 2915 67547 3001 67603
rect 3057 67547 3143 67603
rect 3199 67547 3285 67603
rect 3341 67547 3427 67603
rect 3483 67547 3569 67603
rect 3625 67547 3711 67603
rect 3767 67547 3853 67603
rect 3909 67547 3995 67603
rect 4051 67547 4137 67603
rect 4193 67547 4279 67603
rect 4335 67547 4421 67603
rect 4477 67547 4563 67603
rect 4619 67547 4705 67603
rect 4761 67547 4847 67603
rect 4903 67547 4989 67603
rect 5045 67547 5131 67603
rect 5187 67547 5273 67603
rect 5329 67547 5415 67603
rect 5471 67547 5557 67603
rect 5613 67547 5699 67603
rect 5755 67547 5841 67603
rect 5897 67547 5983 67603
rect 6039 67547 6125 67603
rect 6181 67547 6267 67603
rect 6323 67547 6409 67603
rect 6465 67547 6551 67603
rect 6607 67547 6693 67603
rect 6749 67547 6835 67603
rect 6891 67547 6977 67603
rect 7033 67547 7119 67603
rect 7175 67547 7261 67603
rect 7317 67547 7403 67603
rect 7459 67547 7545 67603
rect 7601 67547 7687 67603
rect 7743 67547 7829 67603
rect 7885 67547 7971 67603
rect 8027 67547 8113 67603
rect 8169 67547 8255 67603
rect 8311 67547 8397 67603
rect 8453 67547 8539 67603
rect 8595 67547 8681 67603
rect 8737 67547 8823 67603
rect 8879 67547 8965 67603
rect 9021 67547 9107 67603
rect 9163 67547 9249 67603
rect 9305 67547 9391 67603
rect 9447 67547 9533 67603
rect 9589 67547 9675 67603
rect 9731 67547 9817 67603
rect 9873 67547 9959 67603
rect 10015 67547 10101 67603
rect 10157 67547 10243 67603
rect 10299 67547 10385 67603
rect 10441 67547 10527 67603
rect 10583 67547 10669 67603
rect 10725 67547 10811 67603
rect 10867 67547 10953 67603
rect 11009 67547 11095 67603
rect 11151 67547 11237 67603
rect 11293 67547 11379 67603
rect 11435 67547 11521 67603
rect 11577 67547 11663 67603
rect 11719 67547 11805 67603
rect 11861 67547 11947 67603
rect 12003 67547 12089 67603
rect 12145 67547 12231 67603
rect 12287 67547 12373 67603
rect 12429 67547 12515 67603
rect 12571 67547 12657 67603
rect 12713 67547 12799 67603
rect 12855 67547 12941 67603
rect 12997 67547 13083 67603
rect 13139 67547 13225 67603
rect 13281 67547 13367 67603
rect 13423 67547 13509 67603
rect 13565 67547 13651 67603
rect 13707 67547 13793 67603
rect 13849 67547 13935 67603
rect 13991 67547 14077 67603
rect 14133 67547 14219 67603
rect 14275 67547 14361 67603
rect 14417 67547 14503 67603
rect 14559 67547 14645 67603
rect 14701 67547 14787 67603
rect 14843 67547 14853 67603
rect 151 67461 14853 67547
rect 151 67405 161 67461
rect 217 67405 303 67461
rect 359 67405 445 67461
rect 501 67405 587 67461
rect 643 67405 729 67461
rect 785 67405 871 67461
rect 927 67405 1013 67461
rect 1069 67405 1155 67461
rect 1211 67405 1297 67461
rect 1353 67405 1439 67461
rect 1495 67405 1581 67461
rect 1637 67405 1723 67461
rect 1779 67405 1865 67461
rect 1921 67405 2007 67461
rect 2063 67405 2149 67461
rect 2205 67405 2291 67461
rect 2347 67405 2433 67461
rect 2489 67405 2575 67461
rect 2631 67405 2717 67461
rect 2773 67405 2859 67461
rect 2915 67405 3001 67461
rect 3057 67405 3143 67461
rect 3199 67405 3285 67461
rect 3341 67405 3427 67461
rect 3483 67405 3569 67461
rect 3625 67405 3711 67461
rect 3767 67405 3853 67461
rect 3909 67405 3995 67461
rect 4051 67405 4137 67461
rect 4193 67405 4279 67461
rect 4335 67405 4421 67461
rect 4477 67405 4563 67461
rect 4619 67405 4705 67461
rect 4761 67405 4847 67461
rect 4903 67405 4989 67461
rect 5045 67405 5131 67461
rect 5187 67405 5273 67461
rect 5329 67405 5415 67461
rect 5471 67405 5557 67461
rect 5613 67405 5699 67461
rect 5755 67405 5841 67461
rect 5897 67405 5983 67461
rect 6039 67405 6125 67461
rect 6181 67405 6267 67461
rect 6323 67405 6409 67461
rect 6465 67405 6551 67461
rect 6607 67405 6693 67461
rect 6749 67405 6835 67461
rect 6891 67405 6977 67461
rect 7033 67405 7119 67461
rect 7175 67405 7261 67461
rect 7317 67405 7403 67461
rect 7459 67405 7545 67461
rect 7601 67405 7687 67461
rect 7743 67405 7829 67461
rect 7885 67405 7971 67461
rect 8027 67405 8113 67461
rect 8169 67405 8255 67461
rect 8311 67405 8397 67461
rect 8453 67405 8539 67461
rect 8595 67405 8681 67461
rect 8737 67405 8823 67461
rect 8879 67405 8965 67461
rect 9021 67405 9107 67461
rect 9163 67405 9249 67461
rect 9305 67405 9391 67461
rect 9447 67405 9533 67461
rect 9589 67405 9675 67461
rect 9731 67405 9817 67461
rect 9873 67405 9959 67461
rect 10015 67405 10101 67461
rect 10157 67405 10243 67461
rect 10299 67405 10385 67461
rect 10441 67405 10527 67461
rect 10583 67405 10669 67461
rect 10725 67405 10811 67461
rect 10867 67405 10953 67461
rect 11009 67405 11095 67461
rect 11151 67405 11237 67461
rect 11293 67405 11379 67461
rect 11435 67405 11521 67461
rect 11577 67405 11663 67461
rect 11719 67405 11805 67461
rect 11861 67405 11947 67461
rect 12003 67405 12089 67461
rect 12145 67405 12231 67461
rect 12287 67405 12373 67461
rect 12429 67405 12515 67461
rect 12571 67405 12657 67461
rect 12713 67405 12799 67461
rect 12855 67405 12941 67461
rect 12997 67405 13083 67461
rect 13139 67405 13225 67461
rect 13281 67405 13367 67461
rect 13423 67405 13509 67461
rect 13565 67405 13651 67461
rect 13707 67405 13793 67461
rect 13849 67405 13935 67461
rect 13991 67405 14077 67461
rect 14133 67405 14219 67461
rect 14275 67405 14361 67461
rect 14417 67405 14503 67461
rect 14559 67405 14645 67461
rect 14701 67405 14787 67461
rect 14843 67405 14853 67461
rect 151 67319 14853 67405
rect 151 67263 161 67319
rect 217 67263 303 67319
rect 359 67263 445 67319
rect 501 67263 587 67319
rect 643 67263 729 67319
rect 785 67263 871 67319
rect 927 67263 1013 67319
rect 1069 67263 1155 67319
rect 1211 67263 1297 67319
rect 1353 67263 1439 67319
rect 1495 67263 1581 67319
rect 1637 67263 1723 67319
rect 1779 67263 1865 67319
rect 1921 67263 2007 67319
rect 2063 67263 2149 67319
rect 2205 67263 2291 67319
rect 2347 67263 2433 67319
rect 2489 67263 2575 67319
rect 2631 67263 2717 67319
rect 2773 67263 2859 67319
rect 2915 67263 3001 67319
rect 3057 67263 3143 67319
rect 3199 67263 3285 67319
rect 3341 67263 3427 67319
rect 3483 67263 3569 67319
rect 3625 67263 3711 67319
rect 3767 67263 3853 67319
rect 3909 67263 3995 67319
rect 4051 67263 4137 67319
rect 4193 67263 4279 67319
rect 4335 67263 4421 67319
rect 4477 67263 4563 67319
rect 4619 67263 4705 67319
rect 4761 67263 4847 67319
rect 4903 67263 4989 67319
rect 5045 67263 5131 67319
rect 5187 67263 5273 67319
rect 5329 67263 5415 67319
rect 5471 67263 5557 67319
rect 5613 67263 5699 67319
rect 5755 67263 5841 67319
rect 5897 67263 5983 67319
rect 6039 67263 6125 67319
rect 6181 67263 6267 67319
rect 6323 67263 6409 67319
rect 6465 67263 6551 67319
rect 6607 67263 6693 67319
rect 6749 67263 6835 67319
rect 6891 67263 6977 67319
rect 7033 67263 7119 67319
rect 7175 67263 7261 67319
rect 7317 67263 7403 67319
rect 7459 67263 7545 67319
rect 7601 67263 7687 67319
rect 7743 67263 7829 67319
rect 7885 67263 7971 67319
rect 8027 67263 8113 67319
rect 8169 67263 8255 67319
rect 8311 67263 8397 67319
rect 8453 67263 8539 67319
rect 8595 67263 8681 67319
rect 8737 67263 8823 67319
rect 8879 67263 8965 67319
rect 9021 67263 9107 67319
rect 9163 67263 9249 67319
rect 9305 67263 9391 67319
rect 9447 67263 9533 67319
rect 9589 67263 9675 67319
rect 9731 67263 9817 67319
rect 9873 67263 9959 67319
rect 10015 67263 10101 67319
rect 10157 67263 10243 67319
rect 10299 67263 10385 67319
rect 10441 67263 10527 67319
rect 10583 67263 10669 67319
rect 10725 67263 10811 67319
rect 10867 67263 10953 67319
rect 11009 67263 11095 67319
rect 11151 67263 11237 67319
rect 11293 67263 11379 67319
rect 11435 67263 11521 67319
rect 11577 67263 11663 67319
rect 11719 67263 11805 67319
rect 11861 67263 11947 67319
rect 12003 67263 12089 67319
rect 12145 67263 12231 67319
rect 12287 67263 12373 67319
rect 12429 67263 12515 67319
rect 12571 67263 12657 67319
rect 12713 67263 12799 67319
rect 12855 67263 12941 67319
rect 12997 67263 13083 67319
rect 13139 67263 13225 67319
rect 13281 67263 13367 67319
rect 13423 67263 13509 67319
rect 13565 67263 13651 67319
rect 13707 67263 13793 67319
rect 13849 67263 13935 67319
rect 13991 67263 14077 67319
rect 14133 67263 14219 67319
rect 14275 67263 14361 67319
rect 14417 67263 14503 67319
rect 14559 67263 14645 67319
rect 14701 67263 14787 67319
rect 14843 67263 14853 67319
rect 151 67177 14853 67263
rect 151 67121 161 67177
rect 217 67121 303 67177
rect 359 67121 445 67177
rect 501 67121 587 67177
rect 643 67121 729 67177
rect 785 67121 871 67177
rect 927 67121 1013 67177
rect 1069 67121 1155 67177
rect 1211 67121 1297 67177
rect 1353 67121 1439 67177
rect 1495 67121 1581 67177
rect 1637 67121 1723 67177
rect 1779 67121 1865 67177
rect 1921 67121 2007 67177
rect 2063 67121 2149 67177
rect 2205 67121 2291 67177
rect 2347 67121 2433 67177
rect 2489 67121 2575 67177
rect 2631 67121 2717 67177
rect 2773 67121 2859 67177
rect 2915 67121 3001 67177
rect 3057 67121 3143 67177
rect 3199 67121 3285 67177
rect 3341 67121 3427 67177
rect 3483 67121 3569 67177
rect 3625 67121 3711 67177
rect 3767 67121 3853 67177
rect 3909 67121 3995 67177
rect 4051 67121 4137 67177
rect 4193 67121 4279 67177
rect 4335 67121 4421 67177
rect 4477 67121 4563 67177
rect 4619 67121 4705 67177
rect 4761 67121 4847 67177
rect 4903 67121 4989 67177
rect 5045 67121 5131 67177
rect 5187 67121 5273 67177
rect 5329 67121 5415 67177
rect 5471 67121 5557 67177
rect 5613 67121 5699 67177
rect 5755 67121 5841 67177
rect 5897 67121 5983 67177
rect 6039 67121 6125 67177
rect 6181 67121 6267 67177
rect 6323 67121 6409 67177
rect 6465 67121 6551 67177
rect 6607 67121 6693 67177
rect 6749 67121 6835 67177
rect 6891 67121 6977 67177
rect 7033 67121 7119 67177
rect 7175 67121 7261 67177
rect 7317 67121 7403 67177
rect 7459 67121 7545 67177
rect 7601 67121 7687 67177
rect 7743 67121 7829 67177
rect 7885 67121 7971 67177
rect 8027 67121 8113 67177
rect 8169 67121 8255 67177
rect 8311 67121 8397 67177
rect 8453 67121 8539 67177
rect 8595 67121 8681 67177
rect 8737 67121 8823 67177
rect 8879 67121 8965 67177
rect 9021 67121 9107 67177
rect 9163 67121 9249 67177
rect 9305 67121 9391 67177
rect 9447 67121 9533 67177
rect 9589 67121 9675 67177
rect 9731 67121 9817 67177
rect 9873 67121 9959 67177
rect 10015 67121 10101 67177
rect 10157 67121 10243 67177
rect 10299 67121 10385 67177
rect 10441 67121 10527 67177
rect 10583 67121 10669 67177
rect 10725 67121 10811 67177
rect 10867 67121 10953 67177
rect 11009 67121 11095 67177
rect 11151 67121 11237 67177
rect 11293 67121 11379 67177
rect 11435 67121 11521 67177
rect 11577 67121 11663 67177
rect 11719 67121 11805 67177
rect 11861 67121 11947 67177
rect 12003 67121 12089 67177
rect 12145 67121 12231 67177
rect 12287 67121 12373 67177
rect 12429 67121 12515 67177
rect 12571 67121 12657 67177
rect 12713 67121 12799 67177
rect 12855 67121 12941 67177
rect 12997 67121 13083 67177
rect 13139 67121 13225 67177
rect 13281 67121 13367 67177
rect 13423 67121 13509 67177
rect 13565 67121 13651 67177
rect 13707 67121 13793 67177
rect 13849 67121 13935 67177
rect 13991 67121 14077 67177
rect 14133 67121 14219 67177
rect 14275 67121 14361 67177
rect 14417 67121 14503 67177
rect 14559 67121 14645 67177
rect 14701 67121 14787 67177
rect 14843 67121 14853 67177
rect 151 67035 14853 67121
rect 151 66979 161 67035
rect 217 66979 303 67035
rect 359 66979 445 67035
rect 501 66979 587 67035
rect 643 66979 729 67035
rect 785 66979 871 67035
rect 927 66979 1013 67035
rect 1069 66979 1155 67035
rect 1211 66979 1297 67035
rect 1353 66979 1439 67035
rect 1495 66979 1581 67035
rect 1637 66979 1723 67035
rect 1779 66979 1865 67035
rect 1921 66979 2007 67035
rect 2063 66979 2149 67035
rect 2205 66979 2291 67035
rect 2347 66979 2433 67035
rect 2489 66979 2575 67035
rect 2631 66979 2717 67035
rect 2773 66979 2859 67035
rect 2915 66979 3001 67035
rect 3057 66979 3143 67035
rect 3199 66979 3285 67035
rect 3341 66979 3427 67035
rect 3483 66979 3569 67035
rect 3625 66979 3711 67035
rect 3767 66979 3853 67035
rect 3909 66979 3995 67035
rect 4051 66979 4137 67035
rect 4193 66979 4279 67035
rect 4335 66979 4421 67035
rect 4477 66979 4563 67035
rect 4619 66979 4705 67035
rect 4761 66979 4847 67035
rect 4903 66979 4989 67035
rect 5045 66979 5131 67035
rect 5187 66979 5273 67035
rect 5329 66979 5415 67035
rect 5471 66979 5557 67035
rect 5613 66979 5699 67035
rect 5755 66979 5841 67035
rect 5897 66979 5983 67035
rect 6039 66979 6125 67035
rect 6181 66979 6267 67035
rect 6323 66979 6409 67035
rect 6465 66979 6551 67035
rect 6607 66979 6693 67035
rect 6749 66979 6835 67035
rect 6891 66979 6977 67035
rect 7033 66979 7119 67035
rect 7175 66979 7261 67035
rect 7317 66979 7403 67035
rect 7459 66979 7545 67035
rect 7601 66979 7687 67035
rect 7743 66979 7829 67035
rect 7885 66979 7971 67035
rect 8027 66979 8113 67035
rect 8169 66979 8255 67035
rect 8311 66979 8397 67035
rect 8453 66979 8539 67035
rect 8595 66979 8681 67035
rect 8737 66979 8823 67035
rect 8879 66979 8965 67035
rect 9021 66979 9107 67035
rect 9163 66979 9249 67035
rect 9305 66979 9391 67035
rect 9447 66979 9533 67035
rect 9589 66979 9675 67035
rect 9731 66979 9817 67035
rect 9873 66979 9959 67035
rect 10015 66979 10101 67035
rect 10157 66979 10243 67035
rect 10299 66979 10385 67035
rect 10441 66979 10527 67035
rect 10583 66979 10669 67035
rect 10725 66979 10811 67035
rect 10867 66979 10953 67035
rect 11009 66979 11095 67035
rect 11151 66979 11237 67035
rect 11293 66979 11379 67035
rect 11435 66979 11521 67035
rect 11577 66979 11663 67035
rect 11719 66979 11805 67035
rect 11861 66979 11947 67035
rect 12003 66979 12089 67035
rect 12145 66979 12231 67035
rect 12287 66979 12373 67035
rect 12429 66979 12515 67035
rect 12571 66979 12657 67035
rect 12713 66979 12799 67035
rect 12855 66979 12941 67035
rect 12997 66979 13083 67035
rect 13139 66979 13225 67035
rect 13281 66979 13367 67035
rect 13423 66979 13509 67035
rect 13565 66979 13651 67035
rect 13707 66979 13793 67035
rect 13849 66979 13935 67035
rect 13991 66979 14077 67035
rect 14133 66979 14219 67035
rect 14275 66979 14361 67035
rect 14417 66979 14503 67035
rect 14559 66979 14645 67035
rect 14701 66979 14787 67035
rect 14843 66979 14853 67035
rect 151 66893 14853 66979
rect 151 66837 161 66893
rect 217 66837 303 66893
rect 359 66837 445 66893
rect 501 66837 587 66893
rect 643 66837 729 66893
rect 785 66837 871 66893
rect 927 66837 1013 66893
rect 1069 66837 1155 66893
rect 1211 66837 1297 66893
rect 1353 66837 1439 66893
rect 1495 66837 1581 66893
rect 1637 66837 1723 66893
rect 1779 66837 1865 66893
rect 1921 66837 2007 66893
rect 2063 66837 2149 66893
rect 2205 66837 2291 66893
rect 2347 66837 2433 66893
rect 2489 66837 2575 66893
rect 2631 66837 2717 66893
rect 2773 66837 2859 66893
rect 2915 66837 3001 66893
rect 3057 66837 3143 66893
rect 3199 66837 3285 66893
rect 3341 66837 3427 66893
rect 3483 66837 3569 66893
rect 3625 66837 3711 66893
rect 3767 66837 3853 66893
rect 3909 66837 3995 66893
rect 4051 66837 4137 66893
rect 4193 66837 4279 66893
rect 4335 66837 4421 66893
rect 4477 66837 4563 66893
rect 4619 66837 4705 66893
rect 4761 66837 4847 66893
rect 4903 66837 4989 66893
rect 5045 66837 5131 66893
rect 5187 66837 5273 66893
rect 5329 66837 5415 66893
rect 5471 66837 5557 66893
rect 5613 66837 5699 66893
rect 5755 66837 5841 66893
rect 5897 66837 5983 66893
rect 6039 66837 6125 66893
rect 6181 66837 6267 66893
rect 6323 66837 6409 66893
rect 6465 66837 6551 66893
rect 6607 66837 6693 66893
rect 6749 66837 6835 66893
rect 6891 66837 6977 66893
rect 7033 66837 7119 66893
rect 7175 66837 7261 66893
rect 7317 66837 7403 66893
rect 7459 66837 7545 66893
rect 7601 66837 7687 66893
rect 7743 66837 7829 66893
rect 7885 66837 7971 66893
rect 8027 66837 8113 66893
rect 8169 66837 8255 66893
rect 8311 66837 8397 66893
rect 8453 66837 8539 66893
rect 8595 66837 8681 66893
rect 8737 66837 8823 66893
rect 8879 66837 8965 66893
rect 9021 66837 9107 66893
rect 9163 66837 9249 66893
rect 9305 66837 9391 66893
rect 9447 66837 9533 66893
rect 9589 66837 9675 66893
rect 9731 66837 9817 66893
rect 9873 66837 9959 66893
rect 10015 66837 10101 66893
rect 10157 66837 10243 66893
rect 10299 66837 10385 66893
rect 10441 66837 10527 66893
rect 10583 66837 10669 66893
rect 10725 66837 10811 66893
rect 10867 66837 10953 66893
rect 11009 66837 11095 66893
rect 11151 66837 11237 66893
rect 11293 66837 11379 66893
rect 11435 66837 11521 66893
rect 11577 66837 11663 66893
rect 11719 66837 11805 66893
rect 11861 66837 11947 66893
rect 12003 66837 12089 66893
rect 12145 66837 12231 66893
rect 12287 66837 12373 66893
rect 12429 66837 12515 66893
rect 12571 66837 12657 66893
rect 12713 66837 12799 66893
rect 12855 66837 12941 66893
rect 12997 66837 13083 66893
rect 13139 66837 13225 66893
rect 13281 66837 13367 66893
rect 13423 66837 13509 66893
rect 13565 66837 13651 66893
rect 13707 66837 13793 66893
rect 13849 66837 13935 66893
rect 13991 66837 14077 66893
rect 14133 66837 14219 66893
rect 14275 66837 14361 66893
rect 14417 66837 14503 66893
rect 14559 66837 14645 66893
rect 14701 66837 14787 66893
rect 14843 66837 14853 66893
rect 151 66827 14853 66837
rect 151 66571 14853 66581
rect 151 66515 161 66571
rect 217 66515 303 66571
rect 359 66515 445 66571
rect 501 66515 587 66571
rect 643 66515 729 66571
rect 785 66515 871 66571
rect 927 66515 1013 66571
rect 1069 66515 1155 66571
rect 1211 66515 1297 66571
rect 1353 66515 1439 66571
rect 1495 66515 1581 66571
rect 1637 66515 1723 66571
rect 1779 66515 1865 66571
rect 1921 66515 2007 66571
rect 2063 66515 2149 66571
rect 2205 66515 2291 66571
rect 2347 66515 2433 66571
rect 2489 66515 2575 66571
rect 2631 66515 2717 66571
rect 2773 66515 2859 66571
rect 2915 66515 3001 66571
rect 3057 66515 3143 66571
rect 3199 66515 3285 66571
rect 3341 66515 3427 66571
rect 3483 66515 3569 66571
rect 3625 66515 3711 66571
rect 3767 66515 3853 66571
rect 3909 66515 3995 66571
rect 4051 66515 4137 66571
rect 4193 66515 4279 66571
rect 4335 66515 4421 66571
rect 4477 66515 4563 66571
rect 4619 66515 4705 66571
rect 4761 66515 4847 66571
rect 4903 66515 4989 66571
rect 5045 66515 5131 66571
rect 5187 66515 5273 66571
rect 5329 66515 5415 66571
rect 5471 66515 5557 66571
rect 5613 66515 5699 66571
rect 5755 66515 5841 66571
rect 5897 66515 5983 66571
rect 6039 66515 6125 66571
rect 6181 66515 6267 66571
rect 6323 66515 6409 66571
rect 6465 66515 6551 66571
rect 6607 66515 6693 66571
rect 6749 66515 6835 66571
rect 6891 66515 6977 66571
rect 7033 66515 7119 66571
rect 7175 66515 7261 66571
rect 7317 66515 7403 66571
rect 7459 66515 7545 66571
rect 7601 66515 7687 66571
rect 7743 66515 7829 66571
rect 7885 66515 7971 66571
rect 8027 66515 8113 66571
rect 8169 66515 8255 66571
rect 8311 66515 8397 66571
rect 8453 66515 8539 66571
rect 8595 66515 8681 66571
rect 8737 66515 8823 66571
rect 8879 66515 8965 66571
rect 9021 66515 9107 66571
rect 9163 66515 9249 66571
rect 9305 66515 9391 66571
rect 9447 66515 9533 66571
rect 9589 66515 9675 66571
rect 9731 66515 9817 66571
rect 9873 66515 9959 66571
rect 10015 66515 10101 66571
rect 10157 66515 10243 66571
rect 10299 66515 10385 66571
rect 10441 66515 10527 66571
rect 10583 66515 10669 66571
rect 10725 66515 10811 66571
rect 10867 66515 10953 66571
rect 11009 66515 11095 66571
rect 11151 66515 11237 66571
rect 11293 66515 11379 66571
rect 11435 66515 11521 66571
rect 11577 66515 11663 66571
rect 11719 66515 11805 66571
rect 11861 66515 11947 66571
rect 12003 66515 12089 66571
rect 12145 66515 12231 66571
rect 12287 66515 12373 66571
rect 12429 66515 12515 66571
rect 12571 66515 12657 66571
rect 12713 66515 12799 66571
rect 12855 66515 12941 66571
rect 12997 66515 13083 66571
rect 13139 66515 13225 66571
rect 13281 66515 13367 66571
rect 13423 66515 13509 66571
rect 13565 66515 13651 66571
rect 13707 66515 13793 66571
rect 13849 66515 13935 66571
rect 13991 66515 14077 66571
rect 14133 66515 14219 66571
rect 14275 66515 14361 66571
rect 14417 66515 14503 66571
rect 14559 66515 14645 66571
rect 14701 66515 14787 66571
rect 14843 66515 14853 66571
rect 151 66429 14853 66515
rect 151 66373 161 66429
rect 217 66373 303 66429
rect 359 66373 445 66429
rect 501 66373 587 66429
rect 643 66373 729 66429
rect 785 66373 871 66429
rect 927 66373 1013 66429
rect 1069 66373 1155 66429
rect 1211 66373 1297 66429
rect 1353 66373 1439 66429
rect 1495 66373 1581 66429
rect 1637 66373 1723 66429
rect 1779 66373 1865 66429
rect 1921 66373 2007 66429
rect 2063 66373 2149 66429
rect 2205 66373 2291 66429
rect 2347 66373 2433 66429
rect 2489 66373 2575 66429
rect 2631 66373 2717 66429
rect 2773 66373 2859 66429
rect 2915 66373 3001 66429
rect 3057 66373 3143 66429
rect 3199 66373 3285 66429
rect 3341 66373 3427 66429
rect 3483 66373 3569 66429
rect 3625 66373 3711 66429
rect 3767 66373 3853 66429
rect 3909 66373 3995 66429
rect 4051 66373 4137 66429
rect 4193 66373 4279 66429
rect 4335 66373 4421 66429
rect 4477 66373 4563 66429
rect 4619 66373 4705 66429
rect 4761 66373 4847 66429
rect 4903 66373 4989 66429
rect 5045 66373 5131 66429
rect 5187 66373 5273 66429
rect 5329 66373 5415 66429
rect 5471 66373 5557 66429
rect 5613 66373 5699 66429
rect 5755 66373 5841 66429
rect 5897 66373 5983 66429
rect 6039 66373 6125 66429
rect 6181 66373 6267 66429
rect 6323 66373 6409 66429
rect 6465 66373 6551 66429
rect 6607 66373 6693 66429
rect 6749 66373 6835 66429
rect 6891 66373 6977 66429
rect 7033 66373 7119 66429
rect 7175 66373 7261 66429
rect 7317 66373 7403 66429
rect 7459 66373 7545 66429
rect 7601 66373 7687 66429
rect 7743 66373 7829 66429
rect 7885 66373 7971 66429
rect 8027 66373 8113 66429
rect 8169 66373 8255 66429
rect 8311 66373 8397 66429
rect 8453 66373 8539 66429
rect 8595 66373 8681 66429
rect 8737 66373 8823 66429
rect 8879 66373 8965 66429
rect 9021 66373 9107 66429
rect 9163 66373 9249 66429
rect 9305 66373 9391 66429
rect 9447 66373 9533 66429
rect 9589 66373 9675 66429
rect 9731 66373 9817 66429
rect 9873 66373 9959 66429
rect 10015 66373 10101 66429
rect 10157 66373 10243 66429
rect 10299 66373 10385 66429
rect 10441 66373 10527 66429
rect 10583 66373 10669 66429
rect 10725 66373 10811 66429
rect 10867 66373 10953 66429
rect 11009 66373 11095 66429
rect 11151 66373 11237 66429
rect 11293 66373 11379 66429
rect 11435 66373 11521 66429
rect 11577 66373 11663 66429
rect 11719 66373 11805 66429
rect 11861 66373 11947 66429
rect 12003 66373 12089 66429
rect 12145 66373 12231 66429
rect 12287 66373 12373 66429
rect 12429 66373 12515 66429
rect 12571 66373 12657 66429
rect 12713 66373 12799 66429
rect 12855 66373 12941 66429
rect 12997 66373 13083 66429
rect 13139 66373 13225 66429
rect 13281 66373 13367 66429
rect 13423 66373 13509 66429
rect 13565 66373 13651 66429
rect 13707 66373 13793 66429
rect 13849 66373 13935 66429
rect 13991 66373 14077 66429
rect 14133 66373 14219 66429
rect 14275 66373 14361 66429
rect 14417 66373 14503 66429
rect 14559 66373 14645 66429
rect 14701 66373 14787 66429
rect 14843 66373 14853 66429
rect 151 66287 14853 66373
rect 151 66231 161 66287
rect 217 66231 303 66287
rect 359 66231 445 66287
rect 501 66231 587 66287
rect 643 66231 729 66287
rect 785 66231 871 66287
rect 927 66231 1013 66287
rect 1069 66231 1155 66287
rect 1211 66231 1297 66287
rect 1353 66231 1439 66287
rect 1495 66231 1581 66287
rect 1637 66231 1723 66287
rect 1779 66231 1865 66287
rect 1921 66231 2007 66287
rect 2063 66231 2149 66287
rect 2205 66231 2291 66287
rect 2347 66231 2433 66287
rect 2489 66231 2575 66287
rect 2631 66231 2717 66287
rect 2773 66231 2859 66287
rect 2915 66231 3001 66287
rect 3057 66231 3143 66287
rect 3199 66231 3285 66287
rect 3341 66231 3427 66287
rect 3483 66231 3569 66287
rect 3625 66231 3711 66287
rect 3767 66231 3853 66287
rect 3909 66231 3995 66287
rect 4051 66231 4137 66287
rect 4193 66231 4279 66287
rect 4335 66231 4421 66287
rect 4477 66231 4563 66287
rect 4619 66231 4705 66287
rect 4761 66231 4847 66287
rect 4903 66231 4989 66287
rect 5045 66231 5131 66287
rect 5187 66231 5273 66287
rect 5329 66231 5415 66287
rect 5471 66231 5557 66287
rect 5613 66231 5699 66287
rect 5755 66231 5841 66287
rect 5897 66231 5983 66287
rect 6039 66231 6125 66287
rect 6181 66231 6267 66287
rect 6323 66231 6409 66287
rect 6465 66231 6551 66287
rect 6607 66231 6693 66287
rect 6749 66231 6835 66287
rect 6891 66231 6977 66287
rect 7033 66231 7119 66287
rect 7175 66231 7261 66287
rect 7317 66231 7403 66287
rect 7459 66231 7545 66287
rect 7601 66231 7687 66287
rect 7743 66231 7829 66287
rect 7885 66231 7971 66287
rect 8027 66231 8113 66287
rect 8169 66231 8255 66287
rect 8311 66231 8397 66287
rect 8453 66231 8539 66287
rect 8595 66231 8681 66287
rect 8737 66231 8823 66287
rect 8879 66231 8965 66287
rect 9021 66231 9107 66287
rect 9163 66231 9249 66287
rect 9305 66231 9391 66287
rect 9447 66231 9533 66287
rect 9589 66231 9675 66287
rect 9731 66231 9817 66287
rect 9873 66231 9959 66287
rect 10015 66231 10101 66287
rect 10157 66231 10243 66287
rect 10299 66231 10385 66287
rect 10441 66231 10527 66287
rect 10583 66231 10669 66287
rect 10725 66231 10811 66287
rect 10867 66231 10953 66287
rect 11009 66231 11095 66287
rect 11151 66231 11237 66287
rect 11293 66231 11379 66287
rect 11435 66231 11521 66287
rect 11577 66231 11663 66287
rect 11719 66231 11805 66287
rect 11861 66231 11947 66287
rect 12003 66231 12089 66287
rect 12145 66231 12231 66287
rect 12287 66231 12373 66287
rect 12429 66231 12515 66287
rect 12571 66231 12657 66287
rect 12713 66231 12799 66287
rect 12855 66231 12941 66287
rect 12997 66231 13083 66287
rect 13139 66231 13225 66287
rect 13281 66231 13367 66287
rect 13423 66231 13509 66287
rect 13565 66231 13651 66287
rect 13707 66231 13793 66287
rect 13849 66231 13935 66287
rect 13991 66231 14077 66287
rect 14133 66231 14219 66287
rect 14275 66231 14361 66287
rect 14417 66231 14503 66287
rect 14559 66231 14645 66287
rect 14701 66231 14787 66287
rect 14843 66231 14853 66287
rect 151 66145 14853 66231
rect 151 66089 161 66145
rect 217 66089 303 66145
rect 359 66089 445 66145
rect 501 66089 587 66145
rect 643 66089 729 66145
rect 785 66089 871 66145
rect 927 66089 1013 66145
rect 1069 66089 1155 66145
rect 1211 66089 1297 66145
rect 1353 66089 1439 66145
rect 1495 66089 1581 66145
rect 1637 66089 1723 66145
rect 1779 66089 1865 66145
rect 1921 66089 2007 66145
rect 2063 66089 2149 66145
rect 2205 66089 2291 66145
rect 2347 66089 2433 66145
rect 2489 66089 2575 66145
rect 2631 66089 2717 66145
rect 2773 66089 2859 66145
rect 2915 66089 3001 66145
rect 3057 66089 3143 66145
rect 3199 66089 3285 66145
rect 3341 66089 3427 66145
rect 3483 66089 3569 66145
rect 3625 66089 3711 66145
rect 3767 66089 3853 66145
rect 3909 66089 3995 66145
rect 4051 66089 4137 66145
rect 4193 66089 4279 66145
rect 4335 66089 4421 66145
rect 4477 66089 4563 66145
rect 4619 66089 4705 66145
rect 4761 66089 4847 66145
rect 4903 66089 4989 66145
rect 5045 66089 5131 66145
rect 5187 66089 5273 66145
rect 5329 66089 5415 66145
rect 5471 66089 5557 66145
rect 5613 66089 5699 66145
rect 5755 66089 5841 66145
rect 5897 66089 5983 66145
rect 6039 66089 6125 66145
rect 6181 66089 6267 66145
rect 6323 66089 6409 66145
rect 6465 66089 6551 66145
rect 6607 66089 6693 66145
rect 6749 66089 6835 66145
rect 6891 66089 6977 66145
rect 7033 66089 7119 66145
rect 7175 66089 7261 66145
rect 7317 66089 7403 66145
rect 7459 66089 7545 66145
rect 7601 66089 7687 66145
rect 7743 66089 7829 66145
rect 7885 66089 7971 66145
rect 8027 66089 8113 66145
rect 8169 66089 8255 66145
rect 8311 66089 8397 66145
rect 8453 66089 8539 66145
rect 8595 66089 8681 66145
rect 8737 66089 8823 66145
rect 8879 66089 8965 66145
rect 9021 66089 9107 66145
rect 9163 66089 9249 66145
rect 9305 66089 9391 66145
rect 9447 66089 9533 66145
rect 9589 66089 9675 66145
rect 9731 66089 9817 66145
rect 9873 66089 9959 66145
rect 10015 66089 10101 66145
rect 10157 66089 10243 66145
rect 10299 66089 10385 66145
rect 10441 66089 10527 66145
rect 10583 66089 10669 66145
rect 10725 66089 10811 66145
rect 10867 66089 10953 66145
rect 11009 66089 11095 66145
rect 11151 66089 11237 66145
rect 11293 66089 11379 66145
rect 11435 66089 11521 66145
rect 11577 66089 11663 66145
rect 11719 66089 11805 66145
rect 11861 66089 11947 66145
rect 12003 66089 12089 66145
rect 12145 66089 12231 66145
rect 12287 66089 12373 66145
rect 12429 66089 12515 66145
rect 12571 66089 12657 66145
rect 12713 66089 12799 66145
rect 12855 66089 12941 66145
rect 12997 66089 13083 66145
rect 13139 66089 13225 66145
rect 13281 66089 13367 66145
rect 13423 66089 13509 66145
rect 13565 66089 13651 66145
rect 13707 66089 13793 66145
rect 13849 66089 13935 66145
rect 13991 66089 14077 66145
rect 14133 66089 14219 66145
rect 14275 66089 14361 66145
rect 14417 66089 14503 66145
rect 14559 66089 14645 66145
rect 14701 66089 14787 66145
rect 14843 66089 14853 66145
rect 151 66003 14853 66089
rect 151 65947 161 66003
rect 217 65947 303 66003
rect 359 65947 445 66003
rect 501 65947 587 66003
rect 643 65947 729 66003
rect 785 65947 871 66003
rect 927 65947 1013 66003
rect 1069 65947 1155 66003
rect 1211 65947 1297 66003
rect 1353 65947 1439 66003
rect 1495 65947 1581 66003
rect 1637 65947 1723 66003
rect 1779 65947 1865 66003
rect 1921 65947 2007 66003
rect 2063 65947 2149 66003
rect 2205 65947 2291 66003
rect 2347 65947 2433 66003
rect 2489 65947 2575 66003
rect 2631 65947 2717 66003
rect 2773 65947 2859 66003
rect 2915 65947 3001 66003
rect 3057 65947 3143 66003
rect 3199 65947 3285 66003
rect 3341 65947 3427 66003
rect 3483 65947 3569 66003
rect 3625 65947 3711 66003
rect 3767 65947 3853 66003
rect 3909 65947 3995 66003
rect 4051 65947 4137 66003
rect 4193 65947 4279 66003
rect 4335 65947 4421 66003
rect 4477 65947 4563 66003
rect 4619 65947 4705 66003
rect 4761 65947 4847 66003
rect 4903 65947 4989 66003
rect 5045 65947 5131 66003
rect 5187 65947 5273 66003
rect 5329 65947 5415 66003
rect 5471 65947 5557 66003
rect 5613 65947 5699 66003
rect 5755 65947 5841 66003
rect 5897 65947 5983 66003
rect 6039 65947 6125 66003
rect 6181 65947 6267 66003
rect 6323 65947 6409 66003
rect 6465 65947 6551 66003
rect 6607 65947 6693 66003
rect 6749 65947 6835 66003
rect 6891 65947 6977 66003
rect 7033 65947 7119 66003
rect 7175 65947 7261 66003
rect 7317 65947 7403 66003
rect 7459 65947 7545 66003
rect 7601 65947 7687 66003
rect 7743 65947 7829 66003
rect 7885 65947 7971 66003
rect 8027 65947 8113 66003
rect 8169 65947 8255 66003
rect 8311 65947 8397 66003
rect 8453 65947 8539 66003
rect 8595 65947 8681 66003
rect 8737 65947 8823 66003
rect 8879 65947 8965 66003
rect 9021 65947 9107 66003
rect 9163 65947 9249 66003
rect 9305 65947 9391 66003
rect 9447 65947 9533 66003
rect 9589 65947 9675 66003
rect 9731 65947 9817 66003
rect 9873 65947 9959 66003
rect 10015 65947 10101 66003
rect 10157 65947 10243 66003
rect 10299 65947 10385 66003
rect 10441 65947 10527 66003
rect 10583 65947 10669 66003
rect 10725 65947 10811 66003
rect 10867 65947 10953 66003
rect 11009 65947 11095 66003
rect 11151 65947 11237 66003
rect 11293 65947 11379 66003
rect 11435 65947 11521 66003
rect 11577 65947 11663 66003
rect 11719 65947 11805 66003
rect 11861 65947 11947 66003
rect 12003 65947 12089 66003
rect 12145 65947 12231 66003
rect 12287 65947 12373 66003
rect 12429 65947 12515 66003
rect 12571 65947 12657 66003
rect 12713 65947 12799 66003
rect 12855 65947 12941 66003
rect 12997 65947 13083 66003
rect 13139 65947 13225 66003
rect 13281 65947 13367 66003
rect 13423 65947 13509 66003
rect 13565 65947 13651 66003
rect 13707 65947 13793 66003
rect 13849 65947 13935 66003
rect 13991 65947 14077 66003
rect 14133 65947 14219 66003
rect 14275 65947 14361 66003
rect 14417 65947 14503 66003
rect 14559 65947 14645 66003
rect 14701 65947 14787 66003
rect 14843 65947 14853 66003
rect 151 65861 14853 65947
rect 151 65805 161 65861
rect 217 65805 303 65861
rect 359 65805 445 65861
rect 501 65805 587 65861
rect 643 65805 729 65861
rect 785 65805 871 65861
rect 927 65805 1013 65861
rect 1069 65805 1155 65861
rect 1211 65805 1297 65861
rect 1353 65805 1439 65861
rect 1495 65805 1581 65861
rect 1637 65805 1723 65861
rect 1779 65805 1865 65861
rect 1921 65805 2007 65861
rect 2063 65805 2149 65861
rect 2205 65805 2291 65861
rect 2347 65805 2433 65861
rect 2489 65805 2575 65861
rect 2631 65805 2717 65861
rect 2773 65805 2859 65861
rect 2915 65805 3001 65861
rect 3057 65805 3143 65861
rect 3199 65805 3285 65861
rect 3341 65805 3427 65861
rect 3483 65805 3569 65861
rect 3625 65805 3711 65861
rect 3767 65805 3853 65861
rect 3909 65805 3995 65861
rect 4051 65805 4137 65861
rect 4193 65805 4279 65861
rect 4335 65805 4421 65861
rect 4477 65805 4563 65861
rect 4619 65805 4705 65861
rect 4761 65805 4847 65861
rect 4903 65805 4989 65861
rect 5045 65805 5131 65861
rect 5187 65805 5273 65861
rect 5329 65805 5415 65861
rect 5471 65805 5557 65861
rect 5613 65805 5699 65861
rect 5755 65805 5841 65861
rect 5897 65805 5983 65861
rect 6039 65805 6125 65861
rect 6181 65805 6267 65861
rect 6323 65805 6409 65861
rect 6465 65805 6551 65861
rect 6607 65805 6693 65861
rect 6749 65805 6835 65861
rect 6891 65805 6977 65861
rect 7033 65805 7119 65861
rect 7175 65805 7261 65861
rect 7317 65805 7403 65861
rect 7459 65805 7545 65861
rect 7601 65805 7687 65861
rect 7743 65805 7829 65861
rect 7885 65805 7971 65861
rect 8027 65805 8113 65861
rect 8169 65805 8255 65861
rect 8311 65805 8397 65861
rect 8453 65805 8539 65861
rect 8595 65805 8681 65861
rect 8737 65805 8823 65861
rect 8879 65805 8965 65861
rect 9021 65805 9107 65861
rect 9163 65805 9249 65861
rect 9305 65805 9391 65861
rect 9447 65805 9533 65861
rect 9589 65805 9675 65861
rect 9731 65805 9817 65861
rect 9873 65805 9959 65861
rect 10015 65805 10101 65861
rect 10157 65805 10243 65861
rect 10299 65805 10385 65861
rect 10441 65805 10527 65861
rect 10583 65805 10669 65861
rect 10725 65805 10811 65861
rect 10867 65805 10953 65861
rect 11009 65805 11095 65861
rect 11151 65805 11237 65861
rect 11293 65805 11379 65861
rect 11435 65805 11521 65861
rect 11577 65805 11663 65861
rect 11719 65805 11805 65861
rect 11861 65805 11947 65861
rect 12003 65805 12089 65861
rect 12145 65805 12231 65861
rect 12287 65805 12373 65861
rect 12429 65805 12515 65861
rect 12571 65805 12657 65861
rect 12713 65805 12799 65861
rect 12855 65805 12941 65861
rect 12997 65805 13083 65861
rect 13139 65805 13225 65861
rect 13281 65805 13367 65861
rect 13423 65805 13509 65861
rect 13565 65805 13651 65861
rect 13707 65805 13793 65861
rect 13849 65805 13935 65861
rect 13991 65805 14077 65861
rect 14133 65805 14219 65861
rect 14275 65805 14361 65861
rect 14417 65805 14503 65861
rect 14559 65805 14645 65861
rect 14701 65805 14787 65861
rect 14843 65805 14853 65861
rect 151 65719 14853 65805
rect 151 65663 161 65719
rect 217 65663 303 65719
rect 359 65663 445 65719
rect 501 65663 587 65719
rect 643 65663 729 65719
rect 785 65663 871 65719
rect 927 65663 1013 65719
rect 1069 65663 1155 65719
rect 1211 65663 1297 65719
rect 1353 65663 1439 65719
rect 1495 65663 1581 65719
rect 1637 65663 1723 65719
rect 1779 65663 1865 65719
rect 1921 65663 2007 65719
rect 2063 65663 2149 65719
rect 2205 65663 2291 65719
rect 2347 65663 2433 65719
rect 2489 65663 2575 65719
rect 2631 65663 2717 65719
rect 2773 65663 2859 65719
rect 2915 65663 3001 65719
rect 3057 65663 3143 65719
rect 3199 65663 3285 65719
rect 3341 65663 3427 65719
rect 3483 65663 3569 65719
rect 3625 65663 3711 65719
rect 3767 65663 3853 65719
rect 3909 65663 3995 65719
rect 4051 65663 4137 65719
rect 4193 65663 4279 65719
rect 4335 65663 4421 65719
rect 4477 65663 4563 65719
rect 4619 65663 4705 65719
rect 4761 65663 4847 65719
rect 4903 65663 4989 65719
rect 5045 65663 5131 65719
rect 5187 65663 5273 65719
rect 5329 65663 5415 65719
rect 5471 65663 5557 65719
rect 5613 65663 5699 65719
rect 5755 65663 5841 65719
rect 5897 65663 5983 65719
rect 6039 65663 6125 65719
rect 6181 65663 6267 65719
rect 6323 65663 6409 65719
rect 6465 65663 6551 65719
rect 6607 65663 6693 65719
rect 6749 65663 6835 65719
rect 6891 65663 6977 65719
rect 7033 65663 7119 65719
rect 7175 65663 7261 65719
rect 7317 65663 7403 65719
rect 7459 65663 7545 65719
rect 7601 65663 7687 65719
rect 7743 65663 7829 65719
rect 7885 65663 7971 65719
rect 8027 65663 8113 65719
rect 8169 65663 8255 65719
rect 8311 65663 8397 65719
rect 8453 65663 8539 65719
rect 8595 65663 8681 65719
rect 8737 65663 8823 65719
rect 8879 65663 8965 65719
rect 9021 65663 9107 65719
rect 9163 65663 9249 65719
rect 9305 65663 9391 65719
rect 9447 65663 9533 65719
rect 9589 65663 9675 65719
rect 9731 65663 9817 65719
rect 9873 65663 9959 65719
rect 10015 65663 10101 65719
rect 10157 65663 10243 65719
rect 10299 65663 10385 65719
rect 10441 65663 10527 65719
rect 10583 65663 10669 65719
rect 10725 65663 10811 65719
rect 10867 65663 10953 65719
rect 11009 65663 11095 65719
rect 11151 65663 11237 65719
rect 11293 65663 11379 65719
rect 11435 65663 11521 65719
rect 11577 65663 11663 65719
rect 11719 65663 11805 65719
rect 11861 65663 11947 65719
rect 12003 65663 12089 65719
rect 12145 65663 12231 65719
rect 12287 65663 12373 65719
rect 12429 65663 12515 65719
rect 12571 65663 12657 65719
rect 12713 65663 12799 65719
rect 12855 65663 12941 65719
rect 12997 65663 13083 65719
rect 13139 65663 13225 65719
rect 13281 65663 13367 65719
rect 13423 65663 13509 65719
rect 13565 65663 13651 65719
rect 13707 65663 13793 65719
rect 13849 65663 13935 65719
rect 13991 65663 14077 65719
rect 14133 65663 14219 65719
rect 14275 65663 14361 65719
rect 14417 65663 14503 65719
rect 14559 65663 14645 65719
rect 14701 65663 14787 65719
rect 14843 65663 14853 65719
rect 151 65577 14853 65663
rect 151 65521 161 65577
rect 217 65521 303 65577
rect 359 65521 445 65577
rect 501 65521 587 65577
rect 643 65521 729 65577
rect 785 65521 871 65577
rect 927 65521 1013 65577
rect 1069 65521 1155 65577
rect 1211 65521 1297 65577
rect 1353 65521 1439 65577
rect 1495 65521 1581 65577
rect 1637 65521 1723 65577
rect 1779 65521 1865 65577
rect 1921 65521 2007 65577
rect 2063 65521 2149 65577
rect 2205 65521 2291 65577
rect 2347 65521 2433 65577
rect 2489 65521 2575 65577
rect 2631 65521 2717 65577
rect 2773 65521 2859 65577
rect 2915 65521 3001 65577
rect 3057 65521 3143 65577
rect 3199 65521 3285 65577
rect 3341 65521 3427 65577
rect 3483 65521 3569 65577
rect 3625 65521 3711 65577
rect 3767 65521 3853 65577
rect 3909 65521 3995 65577
rect 4051 65521 4137 65577
rect 4193 65521 4279 65577
rect 4335 65521 4421 65577
rect 4477 65521 4563 65577
rect 4619 65521 4705 65577
rect 4761 65521 4847 65577
rect 4903 65521 4989 65577
rect 5045 65521 5131 65577
rect 5187 65521 5273 65577
rect 5329 65521 5415 65577
rect 5471 65521 5557 65577
rect 5613 65521 5699 65577
rect 5755 65521 5841 65577
rect 5897 65521 5983 65577
rect 6039 65521 6125 65577
rect 6181 65521 6267 65577
rect 6323 65521 6409 65577
rect 6465 65521 6551 65577
rect 6607 65521 6693 65577
rect 6749 65521 6835 65577
rect 6891 65521 6977 65577
rect 7033 65521 7119 65577
rect 7175 65521 7261 65577
rect 7317 65521 7403 65577
rect 7459 65521 7545 65577
rect 7601 65521 7687 65577
rect 7743 65521 7829 65577
rect 7885 65521 7971 65577
rect 8027 65521 8113 65577
rect 8169 65521 8255 65577
rect 8311 65521 8397 65577
rect 8453 65521 8539 65577
rect 8595 65521 8681 65577
rect 8737 65521 8823 65577
rect 8879 65521 8965 65577
rect 9021 65521 9107 65577
rect 9163 65521 9249 65577
rect 9305 65521 9391 65577
rect 9447 65521 9533 65577
rect 9589 65521 9675 65577
rect 9731 65521 9817 65577
rect 9873 65521 9959 65577
rect 10015 65521 10101 65577
rect 10157 65521 10243 65577
rect 10299 65521 10385 65577
rect 10441 65521 10527 65577
rect 10583 65521 10669 65577
rect 10725 65521 10811 65577
rect 10867 65521 10953 65577
rect 11009 65521 11095 65577
rect 11151 65521 11237 65577
rect 11293 65521 11379 65577
rect 11435 65521 11521 65577
rect 11577 65521 11663 65577
rect 11719 65521 11805 65577
rect 11861 65521 11947 65577
rect 12003 65521 12089 65577
rect 12145 65521 12231 65577
rect 12287 65521 12373 65577
rect 12429 65521 12515 65577
rect 12571 65521 12657 65577
rect 12713 65521 12799 65577
rect 12855 65521 12941 65577
rect 12997 65521 13083 65577
rect 13139 65521 13225 65577
rect 13281 65521 13367 65577
rect 13423 65521 13509 65577
rect 13565 65521 13651 65577
rect 13707 65521 13793 65577
rect 13849 65521 13935 65577
rect 13991 65521 14077 65577
rect 14133 65521 14219 65577
rect 14275 65521 14361 65577
rect 14417 65521 14503 65577
rect 14559 65521 14645 65577
rect 14701 65521 14787 65577
rect 14843 65521 14853 65577
rect 151 65435 14853 65521
rect 151 65379 161 65435
rect 217 65379 303 65435
rect 359 65379 445 65435
rect 501 65379 587 65435
rect 643 65379 729 65435
rect 785 65379 871 65435
rect 927 65379 1013 65435
rect 1069 65379 1155 65435
rect 1211 65379 1297 65435
rect 1353 65379 1439 65435
rect 1495 65379 1581 65435
rect 1637 65379 1723 65435
rect 1779 65379 1865 65435
rect 1921 65379 2007 65435
rect 2063 65379 2149 65435
rect 2205 65379 2291 65435
rect 2347 65379 2433 65435
rect 2489 65379 2575 65435
rect 2631 65379 2717 65435
rect 2773 65379 2859 65435
rect 2915 65379 3001 65435
rect 3057 65379 3143 65435
rect 3199 65379 3285 65435
rect 3341 65379 3427 65435
rect 3483 65379 3569 65435
rect 3625 65379 3711 65435
rect 3767 65379 3853 65435
rect 3909 65379 3995 65435
rect 4051 65379 4137 65435
rect 4193 65379 4279 65435
rect 4335 65379 4421 65435
rect 4477 65379 4563 65435
rect 4619 65379 4705 65435
rect 4761 65379 4847 65435
rect 4903 65379 4989 65435
rect 5045 65379 5131 65435
rect 5187 65379 5273 65435
rect 5329 65379 5415 65435
rect 5471 65379 5557 65435
rect 5613 65379 5699 65435
rect 5755 65379 5841 65435
rect 5897 65379 5983 65435
rect 6039 65379 6125 65435
rect 6181 65379 6267 65435
rect 6323 65379 6409 65435
rect 6465 65379 6551 65435
rect 6607 65379 6693 65435
rect 6749 65379 6835 65435
rect 6891 65379 6977 65435
rect 7033 65379 7119 65435
rect 7175 65379 7261 65435
rect 7317 65379 7403 65435
rect 7459 65379 7545 65435
rect 7601 65379 7687 65435
rect 7743 65379 7829 65435
rect 7885 65379 7971 65435
rect 8027 65379 8113 65435
rect 8169 65379 8255 65435
rect 8311 65379 8397 65435
rect 8453 65379 8539 65435
rect 8595 65379 8681 65435
rect 8737 65379 8823 65435
rect 8879 65379 8965 65435
rect 9021 65379 9107 65435
rect 9163 65379 9249 65435
rect 9305 65379 9391 65435
rect 9447 65379 9533 65435
rect 9589 65379 9675 65435
rect 9731 65379 9817 65435
rect 9873 65379 9959 65435
rect 10015 65379 10101 65435
rect 10157 65379 10243 65435
rect 10299 65379 10385 65435
rect 10441 65379 10527 65435
rect 10583 65379 10669 65435
rect 10725 65379 10811 65435
rect 10867 65379 10953 65435
rect 11009 65379 11095 65435
rect 11151 65379 11237 65435
rect 11293 65379 11379 65435
rect 11435 65379 11521 65435
rect 11577 65379 11663 65435
rect 11719 65379 11805 65435
rect 11861 65379 11947 65435
rect 12003 65379 12089 65435
rect 12145 65379 12231 65435
rect 12287 65379 12373 65435
rect 12429 65379 12515 65435
rect 12571 65379 12657 65435
rect 12713 65379 12799 65435
rect 12855 65379 12941 65435
rect 12997 65379 13083 65435
rect 13139 65379 13225 65435
rect 13281 65379 13367 65435
rect 13423 65379 13509 65435
rect 13565 65379 13651 65435
rect 13707 65379 13793 65435
rect 13849 65379 13935 65435
rect 13991 65379 14077 65435
rect 14133 65379 14219 65435
rect 14275 65379 14361 65435
rect 14417 65379 14503 65435
rect 14559 65379 14645 65435
rect 14701 65379 14787 65435
rect 14843 65379 14853 65435
rect 151 65293 14853 65379
rect 151 65237 161 65293
rect 217 65237 303 65293
rect 359 65237 445 65293
rect 501 65237 587 65293
rect 643 65237 729 65293
rect 785 65237 871 65293
rect 927 65237 1013 65293
rect 1069 65237 1155 65293
rect 1211 65237 1297 65293
rect 1353 65237 1439 65293
rect 1495 65237 1581 65293
rect 1637 65237 1723 65293
rect 1779 65237 1865 65293
rect 1921 65237 2007 65293
rect 2063 65237 2149 65293
rect 2205 65237 2291 65293
rect 2347 65237 2433 65293
rect 2489 65237 2575 65293
rect 2631 65237 2717 65293
rect 2773 65237 2859 65293
rect 2915 65237 3001 65293
rect 3057 65237 3143 65293
rect 3199 65237 3285 65293
rect 3341 65237 3427 65293
rect 3483 65237 3569 65293
rect 3625 65237 3711 65293
rect 3767 65237 3853 65293
rect 3909 65237 3995 65293
rect 4051 65237 4137 65293
rect 4193 65237 4279 65293
rect 4335 65237 4421 65293
rect 4477 65237 4563 65293
rect 4619 65237 4705 65293
rect 4761 65237 4847 65293
rect 4903 65237 4989 65293
rect 5045 65237 5131 65293
rect 5187 65237 5273 65293
rect 5329 65237 5415 65293
rect 5471 65237 5557 65293
rect 5613 65237 5699 65293
rect 5755 65237 5841 65293
rect 5897 65237 5983 65293
rect 6039 65237 6125 65293
rect 6181 65237 6267 65293
rect 6323 65237 6409 65293
rect 6465 65237 6551 65293
rect 6607 65237 6693 65293
rect 6749 65237 6835 65293
rect 6891 65237 6977 65293
rect 7033 65237 7119 65293
rect 7175 65237 7261 65293
rect 7317 65237 7403 65293
rect 7459 65237 7545 65293
rect 7601 65237 7687 65293
rect 7743 65237 7829 65293
rect 7885 65237 7971 65293
rect 8027 65237 8113 65293
rect 8169 65237 8255 65293
rect 8311 65237 8397 65293
rect 8453 65237 8539 65293
rect 8595 65237 8681 65293
rect 8737 65237 8823 65293
rect 8879 65237 8965 65293
rect 9021 65237 9107 65293
rect 9163 65237 9249 65293
rect 9305 65237 9391 65293
rect 9447 65237 9533 65293
rect 9589 65237 9675 65293
rect 9731 65237 9817 65293
rect 9873 65237 9959 65293
rect 10015 65237 10101 65293
rect 10157 65237 10243 65293
rect 10299 65237 10385 65293
rect 10441 65237 10527 65293
rect 10583 65237 10669 65293
rect 10725 65237 10811 65293
rect 10867 65237 10953 65293
rect 11009 65237 11095 65293
rect 11151 65237 11237 65293
rect 11293 65237 11379 65293
rect 11435 65237 11521 65293
rect 11577 65237 11663 65293
rect 11719 65237 11805 65293
rect 11861 65237 11947 65293
rect 12003 65237 12089 65293
rect 12145 65237 12231 65293
rect 12287 65237 12373 65293
rect 12429 65237 12515 65293
rect 12571 65237 12657 65293
rect 12713 65237 12799 65293
rect 12855 65237 12941 65293
rect 12997 65237 13083 65293
rect 13139 65237 13225 65293
rect 13281 65237 13367 65293
rect 13423 65237 13509 65293
rect 13565 65237 13651 65293
rect 13707 65237 13793 65293
rect 13849 65237 13935 65293
rect 13991 65237 14077 65293
rect 14133 65237 14219 65293
rect 14275 65237 14361 65293
rect 14417 65237 14503 65293
rect 14559 65237 14645 65293
rect 14701 65237 14787 65293
rect 14843 65237 14853 65293
rect 151 65227 14853 65237
rect 151 64963 14853 64973
rect 151 64907 161 64963
rect 217 64907 303 64963
rect 359 64907 445 64963
rect 501 64907 587 64963
rect 643 64907 729 64963
rect 785 64907 871 64963
rect 927 64907 1013 64963
rect 1069 64907 1155 64963
rect 1211 64907 1297 64963
rect 1353 64907 1439 64963
rect 1495 64907 1581 64963
rect 1637 64907 1723 64963
rect 1779 64907 1865 64963
rect 1921 64907 2007 64963
rect 2063 64907 2149 64963
rect 2205 64907 2291 64963
rect 2347 64907 2433 64963
rect 2489 64907 2575 64963
rect 2631 64907 2717 64963
rect 2773 64907 2859 64963
rect 2915 64907 3001 64963
rect 3057 64907 3143 64963
rect 3199 64907 3285 64963
rect 3341 64907 3427 64963
rect 3483 64907 3569 64963
rect 3625 64907 3711 64963
rect 3767 64907 3853 64963
rect 3909 64907 3995 64963
rect 4051 64907 4137 64963
rect 4193 64907 4279 64963
rect 4335 64907 4421 64963
rect 4477 64907 4563 64963
rect 4619 64907 4705 64963
rect 4761 64907 4847 64963
rect 4903 64907 4989 64963
rect 5045 64907 5131 64963
rect 5187 64907 5273 64963
rect 5329 64907 5415 64963
rect 5471 64907 5557 64963
rect 5613 64907 5699 64963
rect 5755 64907 5841 64963
rect 5897 64907 5983 64963
rect 6039 64907 6125 64963
rect 6181 64907 6267 64963
rect 6323 64907 6409 64963
rect 6465 64907 6551 64963
rect 6607 64907 6693 64963
rect 6749 64907 6835 64963
rect 6891 64907 6977 64963
rect 7033 64907 7119 64963
rect 7175 64907 7261 64963
rect 7317 64907 7403 64963
rect 7459 64907 7545 64963
rect 7601 64907 7687 64963
rect 7743 64907 7829 64963
rect 7885 64907 7971 64963
rect 8027 64907 8113 64963
rect 8169 64907 8255 64963
rect 8311 64907 8397 64963
rect 8453 64907 8539 64963
rect 8595 64907 8681 64963
rect 8737 64907 8823 64963
rect 8879 64907 8965 64963
rect 9021 64907 9107 64963
rect 9163 64907 9249 64963
rect 9305 64907 9391 64963
rect 9447 64907 9533 64963
rect 9589 64907 9675 64963
rect 9731 64907 9817 64963
rect 9873 64907 9959 64963
rect 10015 64907 10101 64963
rect 10157 64907 10243 64963
rect 10299 64907 10385 64963
rect 10441 64907 10527 64963
rect 10583 64907 10669 64963
rect 10725 64907 10811 64963
rect 10867 64907 10953 64963
rect 11009 64907 11095 64963
rect 11151 64907 11237 64963
rect 11293 64907 11379 64963
rect 11435 64907 11521 64963
rect 11577 64907 11663 64963
rect 11719 64907 11805 64963
rect 11861 64907 11947 64963
rect 12003 64907 12089 64963
rect 12145 64907 12231 64963
rect 12287 64907 12373 64963
rect 12429 64907 12515 64963
rect 12571 64907 12657 64963
rect 12713 64907 12799 64963
rect 12855 64907 12941 64963
rect 12997 64907 13083 64963
rect 13139 64907 13225 64963
rect 13281 64907 13367 64963
rect 13423 64907 13509 64963
rect 13565 64907 13651 64963
rect 13707 64907 13793 64963
rect 13849 64907 13935 64963
rect 13991 64907 14077 64963
rect 14133 64907 14219 64963
rect 14275 64907 14361 64963
rect 14417 64907 14503 64963
rect 14559 64907 14645 64963
rect 14701 64907 14787 64963
rect 14843 64907 14853 64963
rect 151 64821 14853 64907
rect 151 64765 161 64821
rect 217 64765 303 64821
rect 359 64765 445 64821
rect 501 64765 587 64821
rect 643 64765 729 64821
rect 785 64765 871 64821
rect 927 64765 1013 64821
rect 1069 64765 1155 64821
rect 1211 64765 1297 64821
rect 1353 64765 1439 64821
rect 1495 64765 1581 64821
rect 1637 64765 1723 64821
rect 1779 64765 1865 64821
rect 1921 64765 2007 64821
rect 2063 64765 2149 64821
rect 2205 64765 2291 64821
rect 2347 64765 2433 64821
rect 2489 64765 2575 64821
rect 2631 64765 2717 64821
rect 2773 64765 2859 64821
rect 2915 64765 3001 64821
rect 3057 64765 3143 64821
rect 3199 64765 3285 64821
rect 3341 64765 3427 64821
rect 3483 64765 3569 64821
rect 3625 64765 3711 64821
rect 3767 64765 3853 64821
rect 3909 64765 3995 64821
rect 4051 64765 4137 64821
rect 4193 64765 4279 64821
rect 4335 64765 4421 64821
rect 4477 64765 4563 64821
rect 4619 64765 4705 64821
rect 4761 64765 4847 64821
rect 4903 64765 4989 64821
rect 5045 64765 5131 64821
rect 5187 64765 5273 64821
rect 5329 64765 5415 64821
rect 5471 64765 5557 64821
rect 5613 64765 5699 64821
rect 5755 64765 5841 64821
rect 5897 64765 5983 64821
rect 6039 64765 6125 64821
rect 6181 64765 6267 64821
rect 6323 64765 6409 64821
rect 6465 64765 6551 64821
rect 6607 64765 6693 64821
rect 6749 64765 6835 64821
rect 6891 64765 6977 64821
rect 7033 64765 7119 64821
rect 7175 64765 7261 64821
rect 7317 64765 7403 64821
rect 7459 64765 7545 64821
rect 7601 64765 7687 64821
rect 7743 64765 7829 64821
rect 7885 64765 7971 64821
rect 8027 64765 8113 64821
rect 8169 64765 8255 64821
rect 8311 64765 8397 64821
rect 8453 64765 8539 64821
rect 8595 64765 8681 64821
rect 8737 64765 8823 64821
rect 8879 64765 8965 64821
rect 9021 64765 9107 64821
rect 9163 64765 9249 64821
rect 9305 64765 9391 64821
rect 9447 64765 9533 64821
rect 9589 64765 9675 64821
rect 9731 64765 9817 64821
rect 9873 64765 9959 64821
rect 10015 64765 10101 64821
rect 10157 64765 10243 64821
rect 10299 64765 10385 64821
rect 10441 64765 10527 64821
rect 10583 64765 10669 64821
rect 10725 64765 10811 64821
rect 10867 64765 10953 64821
rect 11009 64765 11095 64821
rect 11151 64765 11237 64821
rect 11293 64765 11379 64821
rect 11435 64765 11521 64821
rect 11577 64765 11663 64821
rect 11719 64765 11805 64821
rect 11861 64765 11947 64821
rect 12003 64765 12089 64821
rect 12145 64765 12231 64821
rect 12287 64765 12373 64821
rect 12429 64765 12515 64821
rect 12571 64765 12657 64821
rect 12713 64765 12799 64821
rect 12855 64765 12941 64821
rect 12997 64765 13083 64821
rect 13139 64765 13225 64821
rect 13281 64765 13367 64821
rect 13423 64765 13509 64821
rect 13565 64765 13651 64821
rect 13707 64765 13793 64821
rect 13849 64765 13935 64821
rect 13991 64765 14077 64821
rect 14133 64765 14219 64821
rect 14275 64765 14361 64821
rect 14417 64765 14503 64821
rect 14559 64765 14645 64821
rect 14701 64765 14787 64821
rect 14843 64765 14853 64821
rect 151 64679 14853 64765
rect 151 64623 161 64679
rect 217 64623 303 64679
rect 359 64623 445 64679
rect 501 64623 587 64679
rect 643 64623 729 64679
rect 785 64623 871 64679
rect 927 64623 1013 64679
rect 1069 64623 1155 64679
rect 1211 64623 1297 64679
rect 1353 64623 1439 64679
rect 1495 64623 1581 64679
rect 1637 64623 1723 64679
rect 1779 64623 1865 64679
rect 1921 64623 2007 64679
rect 2063 64623 2149 64679
rect 2205 64623 2291 64679
rect 2347 64623 2433 64679
rect 2489 64623 2575 64679
rect 2631 64623 2717 64679
rect 2773 64623 2859 64679
rect 2915 64623 3001 64679
rect 3057 64623 3143 64679
rect 3199 64623 3285 64679
rect 3341 64623 3427 64679
rect 3483 64623 3569 64679
rect 3625 64623 3711 64679
rect 3767 64623 3853 64679
rect 3909 64623 3995 64679
rect 4051 64623 4137 64679
rect 4193 64623 4279 64679
rect 4335 64623 4421 64679
rect 4477 64623 4563 64679
rect 4619 64623 4705 64679
rect 4761 64623 4847 64679
rect 4903 64623 4989 64679
rect 5045 64623 5131 64679
rect 5187 64623 5273 64679
rect 5329 64623 5415 64679
rect 5471 64623 5557 64679
rect 5613 64623 5699 64679
rect 5755 64623 5841 64679
rect 5897 64623 5983 64679
rect 6039 64623 6125 64679
rect 6181 64623 6267 64679
rect 6323 64623 6409 64679
rect 6465 64623 6551 64679
rect 6607 64623 6693 64679
rect 6749 64623 6835 64679
rect 6891 64623 6977 64679
rect 7033 64623 7119 64679
rect 7175 64623 7261 64679
rect 7317 64623 7403 64679
rect 7459 64623 7545 64679
rect 7601 64623 7687 64679
rect 7743 64623 7829 64679
rect 7885 64623 7971 64679
rect 8027 64623 8113 64679
rect 8169 64623 8255 64679
rect 8311 64623 8397 64679
rect 8453 64623 8539 64679
rect 8595 64623 8681 64679
rect 8737 64623 8823 64679
rect 8879 64623 8965 64679
rect 9021 64623 9107 64679
rect 9163 64623 9249 64679
rect 9305 64623 9391 64679
rect 9447 64623 9533 64679
rect 9589 64623 9675 64679
rect 9731 64623 9817 64679
rect 9873 64623 9959 64679
rect 10015 64623 10101 64679
rect 10157 64623 10243 64679
rect 10299 64623 10385 64679
rect 10441 64623 10527 64679
rect 10583 64623 10669 64679
rect 10725 64623 10811 64679
rect 10867 64623 10953 64679
rect 11009 64623 11095 64679
rect 11151 64623 11237 64679
rect 11293 64623 11379 64679
rect 11435 64623 11521 64679
rect 11577 64623 11663 64679
rect 11719 64623 11805 64679
rect 11861 64623 11947 64679
rect 12003 64623 12089 64679
rect 12145 64623 12231 64679
rect 12287 64623 12373 64679
rect 12429 64623 12515 64679
rect 12571 64623 12657 64679
rect 12713 64623 12799 64679
rect 12855 64623 12941 64679
rect 12997 64623 13083 64679
rect 13139 64623 13225 64679
rect 13281 64623 13367 64679
rect 13423 64623 13509 64679
rect 13565 64623 13651 64679
rect 13707 64623 13793 64679
rect 13849 64623 13935 64679
rect 13991 64623 14077 64679
rect 14133 64623 14219 64679
rect 14275 64623 14361 64679
rect 14417 64623 14503 64679
rect 14559 64623 14645 64679
rect 14701 64623 14787 64679
rect 14843 64623 14853 64679
rect 151 64537 14853 64623
rect 151 64481 161 64537
rect 217 64481 303 64537
rect 359 64481 445 64537
rect 501 64481 587 64537
rect 643 64481 729 64537
rect 785 64481 871 64537
rect 927 64481 1013 64537
rect 1069 64481 1155 64537
rect 1211 64481 1297 64537
rect 1353 64481 1439 64537
rect 1495 64481 1581 64537
rect 1637 64481 1723 64537
rect 1779 64481 1865 64537
rect 1921 64481 2007 64537
rect 2063 64481 2149 64537
rect 2205 64481 2291 64537
rect 2347 64481 2433 64537
rect 2489 64481 2575 64537
rect 2631 64481 2717 64537
rect 2773 64481 2859 64537
rect 2915 64481 3001 64537
rect 3057 64481 3143 64537
rect 3199 64481 3285 64537
rect 3341 64481 3427 64537
rect 3483 64481 3569 64537
rect 3625 64481 3711 64537
rect 3767 64481 3853 64537
rect 3909 64481 3995 64537
rect 4051 64481 4137 64537
rect 4193 64481 4279 64537
rect 4335 64481 4421 64537
rect 4477 64481 4563 64537
rect 4619 64481 4705 64537
rect 4761 64481 4847 64537
rect 4903 64481 4989 64537
rect 5045 64481 5131 64537
rect 5187 64481 5273 64537
rect 5329 64481 5415 64537
rect 5471 64481 5557 64537
rect 5613 64481 5699 64537
rect 5755 64481 5841 64537
rect 5897 64481 5983 64537
rect 6039 64481 6125 64537
rect 6181 64481 6267 64537
rect 6323 64481 6409 64537
rect 6465 64481 6551 64537
rect 6607 64481 6693 64537
rect 6749 64481 6835 64537
rect 6891 64481 6977 64537
rect 7033 64481 7119 64537
rect 7175 64481 7261 64537
rect 7317 64481 7403 64537
rect 7459 64481 7545 64537
rect 7601 64481 7687 64537
rect 7743 64481 7829 64537
rect 7885 64481 7971 64537
rect 8027 64481 8113 64537
rect 8169 64481 8255 64537
rect 8311 64481 8397 64537
rect 8453 64481 8539 64537
rect 8595 64481 8681 64537
rect 8737 64481 8823 64537
rect 8879 64481 8965 64537
rect 9021 64481 9107 64537
rect 9163 64481 9249 64537
rect 9305 64481 9391 64537
rect 9447 64481 9533 64537
rect 9589 64481 9675 64537
rect 9731 64481 9817 64537
rect 9873 64481 9959 64537
rect 10015 64481 10101 64537
rect 10157 64481 10243 64537
rect 10299 64481 10385 64537
rect 10441 64481 10527 64537
rect 10583 64481 10669 64537
rect 10725 64481 10811 64537
rect 10867 64481 10953 64537
rect 11009 64481 11095 64537
rect 11151 64481 11237 64537
rect 11293 64481 11379 64537
rect 11435 64481 11521 64537
rect 11577 64481 11663 64537
rect 11719 64481 11805 64537
rect 11861 64481 11947 64537
rect 12003 64481 12089 64537
rect 12145 64481 12231 64537
rect 12287 64481 12373 64537
rect 12429 64481 12515 64537
rect 12571 64481 12657 64537
rect 12713 64481 12799 64537
rect 12855 64481 12941 64537
rect 12997 64481 13083 64537
rect 13139 64481 13225 64537
rect 13281 64481 13367 64537
rect 13423 64481 13509 64537
rect 13565 64481 13651 64537
rect 13707 64481 13793 64537
rect 13849 64481 13935 64537
rect 13991 64481 14077 64537
rect 14133 64481 14219 64537
rect 14275 64481 14361 64537
rect 14417 64481 14503 64537
rect 14559 64481 14645 64537
rect 14701 64481 14787 64537
rect 14843 64481 14853 64537
rect 151 64395 14853 64481
rect 151 64339 161 64395
rect 217 64339 303 64395
rect 359 64339 445 64395
rect 501 64339 587 64395
rect 643 64339 729 64395
rect 785 64339 871 64395
rect 927 64339 1013 64395
rect 1069 64339 1155 64395
rect 1211 64339 1297 64395
rect 1353 64339 1439 64395
rect 1495 64339 1581 64395
rect 1637 64339 1723 64395
rect 1779 64339 1865 64395
rect 1921 64339 2007 64395
rect 2063 64339 2149 64395
rect 2205 64339 2291 64395
rect 2347 64339 2433 64395
rect 2489 64339 2575 64395
rect 2631 64339 2717 64395
rect 2773 64339 2859 64395
rect 2915 64339 3001 64395
rect 3057 64339 3143 64395
rect 3199 64339 3285 64395
rect 3341 64339 3427 64395
rect 3483 64339 3569 64395
rect 3625 64339 3711 64395
rect 3767 64339 3853 64395
rect 3909 64339 3995 64395
rect 4051 64339 4137 64395
rect 4193 64339 4279 64395
rect 4335 64339 4421 64395
rect 4477 64339 4563 64395
rect 4619 64339 4705 64395
rect 4761 64339 4847 64395
rect 4903 64339 4989 64395
rect 5045 64339 5131 64395
rect 5187 64339 5273 64395
rect 5329 64339 5415 64395
rect 5471 64339 5557 64395
rect 5613 64339 5699 64395
rect 5755 64339 5841 64395
rect 5897 64339 5983 64395
rect 6039 64339 6125 64395
rect 6181 64339 6267 64395
rect 6323 64339 6409 64395
rect 6465 64339 6551 64395
rect 6607 64339 6693 64395
rect 6749 64339 6835 64395
rect 6891 64339 6977 64395
rect 7033 64339 7119 64395
rect 7175 64339 7261 64395
rect 7317 64339 7403 64395
rect 7459 64339 7545 64395
rect 7601 64339 7687 64395
rect 7743 64339 7829 64395
rect 7885 64339 7971 64395
rect 8027 64339 8113 64395
rect 8169 64339 8255 64395
rect 8311 64339 8397 64395
rect 8453 64339 8539 64395
rect 8595 64339 8681 64395
rect 8737 64339 8823 64395
rect 8879 64339 8965 64395
rect 9021 64339 9107 64395
rect 9163 64339 9249 64395
rect 9305 64339 9391 64395
rect 9447 64339 9533 64395
rect 9589 64339 9675 64395
rect 9731 64339 9817 64395
rect 9873 64339 9959 64395
rect 10015 64339 10101 64395
rect 10157 64339 10243 64395
rect 10299 64339 10385 64395
rect 10441 64339 10527 64395
rect 10583 64339 10669 64395
rect 10725 64339 10811 64395
rect 10867 64339 10953 64395
rect 11009 64339 11095 64395
rect 11151 64339 11237 64395
rect 11293 64339 11379 64395
rect 11435 64339 11521 64395
rect 11577 64339 11663 64395
rect 11719 64339 11805 64395
rect 11861 64339 11947 64395
rect 12003 64339 12089 64395
rect 12145 64339 12231 64395
rect 12287 64339 12373 64395
rect 12429 64339 12515 64395
rect 12571 64339 12657 64395
rect 12713 64339 12799 64395
rect 12855 64339 12941 64395
rect 12997 64339 13083 64395
rect 13139 64339 13225 64395
rect 13281 64339 13367 64395
rect 13423 64339 13509 64395
rect 13565 64339 13651 64395
rect 13707 64339 13793 64395
rect 13849 64339 13935 64395
rect 13991 64339 14077 64395
rect 14133 64339 14219 64395
rect 14275 64339 14361 64395
rect 14417 64339 14503 64395
rect 14559 64339 14645 64395
rect 14701 64339 14787 64395
rect 14843 64339 14853 64395
rect 151 64253 14853 64339
rect 151 64197 161 64253
rect 217 64197 303 64253
rect 359 64197 445 64253
rect 501 64197 587 64253
rect 643 64197 729 64253
rect 785 64197 871 64253
rect 927 64197 1013 64253
rect 1069 64197 1155 64253
rect 1211 64197 1297 64253
rect 1353 64197 1439 64253
rect 1495 64197 1581 64253
rect 1637 64197 1723 64253
rect 1779 64197 1865 64253
rect 1921 64197 2007 64253
rect 2063 64197 2149 64253
rect 2205 64197 2291 64253
rect 2347 64197 2433 64253
rect 2489 64197 2575 64253
rect 2631 64197 2717 64253
rect 2773 64197 2859 64253
rect 2915 64197 3001 64253
rect 3057 64197 3143 64253
rect 3199 64197 3285 64253
rect 3341 64197 3427 64253
rect 3483 64197 3569 64253
rect 3625 64197 3711 64253
rect 3767 64197 3853 64253
rect 3909 64197 3995 64253
rect 4051 64197 4137 64253
rect 4193 64197 4279 64253
rect 4335 64197 4421 64253
rect 4477 64197 4563 64253
rect 4619 64197 4705 64253
rect 4761 64197 4847 64253
rect 4903 64197 4989 64253
rect 5045 64197 5131 64253
rect 5187 64197 5273 64253
rect 5329 64197 5415 64253
rect 5471 64197 5557 64253
rect 5613 64197 5699 64253
rect 5755 64197 5841 64253
rect 5897 64197 5983 64253
rect 6039 64197 6125 64253
rect 6181 64197 6267 64253
rect 6323 64197 6409 64253
rect 6465 64197 6551 64253
rect 6607 64197 6693 64253
rect 6749 64197 6835 64253
rect 6891 64197 6977 64253
rect 7033 64197 7119 64253
rect 7175 64197 7261 64253
rect 7317 64197 7403 64253
rect 7459 64197 7545 64253
rect 7601 64197 7687 64253
rect 7743 64197 7829 64253
rect 7885 64197 7971 64253
rect 8027 64197 8113 64253
rect 8169 64197 8255 64253
rect 8311 64197 8397 64253
rect 8453 64197 8539 64253
rect 8595 64197 8681 64253
rect 8737 64197 8823 64253
rect 8879 64197 8965 64253
rect 9021 64197 9107 64253
rect 9163 64197 9249 64253
rect 9305 64197 9391 64253
rect 9447 64197 9533 64253
rect 9589 64197 9675 64253
rect 9731 64197 9817 64253
rect 9873 64197 9959 64253
rect 10015 64197 10101 64253
rect 10157 64197 10243 64253
rect 10299 64197 10385 64253
rect 10441 64197 10527 64253
rect 10583 64197 10669 64253
rect 10725 64197 10811 64253
rect 10867 64197 10953 64253
rect 11009 64197 11095 64253
rect 11151 64197 11237 64253
rect 11293 64197 11379 64253
rect 11435 64197 11521 64253
rect 11577 64197 11663 64253
rect 11719 64197 11805 64253
rect 11861 64197 11947 64253
rect 12003 64197 12089 64253
rect 12145 64197 12231 64253
rect 12287 64197 12373 64253
rect 12429 64197 12515 64253
rect 12571 64197 12657 64253
rect 12713 64197 12799 64253
rect 12855 64197 12941 64253
rect 12997 64197 13083 64253
rect 13139 64197 13225 64253
rect 13281 64197 13367 64253
rect 13423 64197 13509 64253
rect 13565 64197 13651 64253
rect 13707 64197 13793 64253
rect 13849 64197 13935 64253
rect 13991 64197 14077 64253
rect 14133 64197 14219 64253
rect 14275 64197 14361 64253
rect 14417 64197 14503 64253
rect 14559 64197 14645 64253
rect 14701 64197 14787 64253
rect 14843 64197 14853 64253
rect 151 64111 14853 64197
rect 151 64055 161 64111
rect 217 64055 303 64111
rect 359 64055 445 64111
rect 501 64055 587 64111
rect 643 64055 729 64111
rect 785 64055 871 64111
rect 927 64055 1013 64111
rect 1069 64055 1155 64111
rect 1211 64055 1297 64111
rect 1353 64055 1439 64111
rect 1495 64055 1581 64111
rect 1637 64055 1723 64111
rect 1779 64055 1865 64111
rect 1921 64055 2007 64111
rect 2063 64055 2149 64111
rect 2205 64055 2291 64111
rect 2347 64055 2433 64111
rect 2489 64055 2575 64111
rect 2631 64055 2717 64111
rect 2773 64055 2859 64111
rect 2915 64055 3001 64111
rect 3057 64055 3143 64111
rect 3199 64055 3285 64111
rect 3341 64055 3427 64111
rect 3483 64055 3569 64111
rect 3625 64055 3711 64111
rect 3767 64055 3853 64111
rect 3909 64055 3995 64111
rect 4051 64055 4137 64111
rect 4193 64055 4279 64111
rect 4335 64055 4421 64111
rect 4477 64055 4563 64111
rect 4619 64055 4705 64111
rect 4761 64055 4847 64111
rect 4903 64055 4989 64111
rect 5045 64055 5131 64111
rect 5187 64055 5273 64111
rect 5329 64055 5415 64111
rect 5471 64055 5557 64111
rect 5613 64055 5699 64111
rect 5755 64055 5841 64111
rect 5897 64055 5983 64111
rect 6039 64055 6125 64111
rect 6181 64055 6267 64111
rect 6323 64055 6409 64111
rect 6465 64055 6551 64111
rect 6607 64055 6693 64111
rect 6749 64055 6835 64111
rect 6891 64055 6977 64111
rect 7033 64055 7119 64111
rect 7175 64055 7261 64111
rect 7317 64055 7403 64111
rect 7459 64055 7545 64111
rect 7601 64055 7687 64111
rect 7743 64055 7829 64111
rect 7885 64055 7971 64111
rect 8027 64055 8113 64111
rect 8169 64055 8255 64111
rect 8311 64055 8397 64111
rect 8453 64055 8539 64111
rect 8595 64055 8681 64111
rect 8737 64055 8823 64111
rect 8879 64055 8965 64111
rect 9021 64055 9107 64111
rect 9163 64055 9249 64111
rect 9305 64055 9391 64111
rect 9447 64055 9533 64111
rect 9589 64055 9675 64111
rect 9731 64055 9817 64111
rect 9873 64055 9959 64111
rect 10015 64055 10101 64111
rect 10157 64055 10243 64111
rect 10299 64055 10385 64111
rect 10441 64055 10527 64111
rect 10583 64055 10669 64111
rect 10725 64055 10811 64111
rect 10867 64055 10953 64111
rect 11009 64055 11095 64111
rect 11151 64055 11237 64111
rect 11293 64055 11379 64111
rect 11435 64055 11521 64111
rect 11577 64055 11663 64111
rect 11719 64055 11805 64111
rect 11861 64055 11947 64111
rect 12003 64055 12089 64111
rect 12145 64055 12231 64111
rect 12287 64055 12373 64111
rect 12429 64055 12515 64111
rect 12571 64055 12657 64111
rect 12713 64055 12799 64111
rect 12855 64055 12941 64111
rect 12997 64055 13083 64111
rect 13139 64055 13225 64111
rect 13281 64055 13367 64111
rect 13423 64055 13509 64111
rect 13565 64055 13651 64111
rect 13707 64055 13793 64111
rect 13849 64055 13935 64111
rect 13991 64055 14077 64111
rect 14133 64055 14219 64111
rect 14275 64055 14361 64111
rect 14417 64055 14503 64111
rect 14559 64055 14645 64111
rect 14701 64055 14787 64111
rect 14843 64055 14853 64111
rect 151 63969 14853 64055
rect 151 63913 161 63969
rect 217 63913 303 63969
rect 359 63913 445 63969
rect 501 63913 587 63969
rect 643 63913 729 63969
rect 785 63913 871 63969
rect 927 63913 1013 63969
rect 1069 63913 1155 63969
rect 1211 63913 1297 63969
rect 1353 63913 1439 63969
rect 1495 63913 1581 63969
rect 1637 63913 1723 63969
rect 1779 63913 1865 63969
rect 1921 63913 2007 63969
rect 2063 63913 2149 63969
rect 2205 63913 2291 63969
rect 2347 63913 2433 63969
rect 2489 63913 2575 63969
rect 2631 63913 2717 63969
rect 2773 63913 2859 63969
rect 2915 63913 3001 63969
rect 3057 63913 3143 63969
rect 3199 63913 3285 63969
rect 3341 63913 3427 63969
rect 3483 63913 3569 63969
rect 3625 63913 3711 63969
rect 3767 63913 3853 63969
rect 3909 63913 3995 63969
rect 4051 63913 4137 63969
rect 4193 63913 4279 63969
rect 4335 63913 4421 63969
rect 4477 63913 4563 63969
rect 4619 63913 4705 63969
rect 4761 63913 4847 63969
rect 4903 63913 4989 63969
rect 5045 63913 5131 63969
rect 5187 63913 5273 63969
rect 5329 63913 5415 63969
rect 5471 63913 5557 63969
rect 5613 63913 5699 63969
rect 5755 63913 5841 63969
rect 5897 63913 5983 63969
rect 6039 63913 6125 63969
rect 6181 63913 6267 63969
rect 6323 63913 6409 63969
rect 6465 63913 6551 63969
rect 6607 63913 6693 63969
rect 6749 63913 6835 63969
rect 6891 63913 6977 63969
rect 7033 63913 7119 63969
rect 7175 63913 7261 63969
rect 7317 63913 7403 63969
rect 7459 63913 7545 63969
rect 7601 63913 7687 63969
rect 7743 63913 7829 63969
rect 7885 63913 7971 63969
rect 8027 63913 8113 63969
rect 8169 63913 8255 63969
rect 8311 63913 8397 63969
rect 8453 63913 8539 63969
rect 8595 63913 8681 63969
rect 8737 63913 8823 63969
rect 8879 63913 8965 63969
rect 9021 63913 9107 63969
rect 9163 63913 9249 63969
rect 9305 63913 9391 63969
rect 9447 63913 9533 63969
rect 9589 63913 9675 63969
rect 9731 63913 9817 63969
rect 9873 63913 9959 63969
rect 10015 63913 10101 63969
rect 10157 63913 10243 63969
rect 10299 63913 10385 63969
rect 10441 63913 10527 63969
rect 10583 63913 10669 63969
rect 10725 63913 10811 63969
rect 10867 63913 10953 63969
rect 11009 63913 11095 63969
rect 11151 63913 11237 63969
rect 11293 63913 11379 63969
rect 11435 63913 11521 63969
rect 11577 63913 11663 63969
rect 11719 63913 11805 63969
rect 11861 63913 11947 63969
rect 12003 63913 12089 63969
rect 12145 63913 12231 63969
rect 12287 63913 12373 63969
rect 12429 63913 12515 63969
rect 12571 63913 12657 63969
rect 12713 63913 12799 63969
rect 12855 63913 12941 63969
rect 12997 63913 13083 63969
rect 13139 63913 13225 63969
rect 13281 63913 13367 63969
rect 13423 63913 13509 63969
rect 13565 63913 13651 63969
rect 13707 63913 13793 63969
rect 13849 63913 13935 63969
rect 13991 63913 14077 63969
rect 14133 63913 14219 63969
rect 14275 63913 14361 63969
rect 14417 63913 14503 63969
rect 14559 63913 14645 63969
rect 14701 63913 14787 63969
rect 14843 63913 14853 63969
rect 151 63827 14853 63913
rect 151 63771 161 63827
rect 217 63771 303 63827
rect 359 63771 445 63827
rect 501 63771 587 63827
rect 643 63771 729 63827
rect 785 63771 871 63827
rect 927 63771 1013 63827
rect 1069 63771 1155 63827
rect 1211 63771 1297 63827
rect 1353 63771 1439 63827
rect 1495 63771 1581 63827
rect 1637 63771 1723 63827
rect 1779 63771 1865 63827
rect 1921 63771 2007 63827
rect 2063 63771 2149 63827
rect 2205 63771 2291 63827
rect 2347 63771 2433 63827
rect 2489 63771 2575 63827
rect 2631 63771 2717 63827
rect 2773 63771 2859 63827
rect 2915 63771 3001 63827
rect 3057 63771 3143 63827
rect 3199 63771 3285 63827
rect 3341 63771 3427 63827
rect 3483 63771 3569 63827
rect 3625 63771 3711 63827
rect 3767 63771 3853 63827
rect 3909 63771 3995 63827
rect 4051 63771 4137 63827
rect 4193 63771 4279 63827
rect 4335 63771 4421 63827
rect 4477 63771 4563 63827
rect 4619 63771 4705 63827
rect 4761 63771 4847 63827
rect 4903 63771 4989 63827
rect 5045 63771 5131 63827
rect 5187 63771 5273 63827
rect 5329 63771 5415 63827
rect 5471 63771 5557 63827
rect 5613 63771 5699 63827
rect 5755 63771 5841 63827
rect 5897 63771 5983 63827
rect 6039 63771 6125 63827
rect 6181 63771 6267 63827
rect 6323 63771 6409 63827
rect 6465 63771 6551 63827
rect 6607 63771 6693 63827
rect 6749 63771 6835 63827
rect 6891 63771 6977 63827
rect 7033 63771 7119 63827
rect 7175 63771 7261 63827
rect 7317 63771 7403 63827
rect 7459 63771 7545 63827
rect 7601 63771 7687 63827
rect 7743 63771 7829 63827
rect 7885 63771 7971 63827
rect 8027 63771 8113 63827
rect 8169 63771 8255 63827
rect 8311 63771 8397 63827
rect 8453 63771 8539 63827
rect 8595 63771 8681 63827
rect 8737 63771 8823 63827
rect 8879 63771 8965 63827
rect 9021 63771 9107 63827
rect 9163 63771 9249 63827
rect 9305 63771 9391 63827
rect 9447 63771 9533 63827
rect 9589 63771 9675 63827
rect 9731 63771 9817 63827
rect 9873 63771 9959 63827
rect 10015 63771 10101 63827
rect 10157 63771 10243 63827
rect 10299 63771 10385 63827
rect 10441 63771 10527 63827
rect 10583 63771 10669 63827
rect 10725 63771 10811 63827
rect 10867 63771 10953 63827
rect 11009 63771 11095 63827
rect 11151 63771 11237 63827
rect 11293 63771 11379 63827
rect 11435 63771 11521 63827
rect 11577 63771 11663 63827
rect 11719 63771 11805 63827
rect 11861 63771 11947 63827
rect 12003 63771 12089 63827
rect 12145 63771 12231 63827
rect 12287 63771 12373 63827
rect 12429 63771 12515 63827
rect 12571 63771 12657 63827
rect 12713 63771 12799 63827
rect 12855 63771 12941 63827
rect 12997 63771 13083 63827
rect 13139 63771 13225 63827
rect 13281 63771 13367 63827
rect 13423 63771 13509 63827
rect 13565 63771 13651 63827
rect 13707 63771 13793 63827
rect 13849 63771 13935 63827
rect 13991 63771 14077 63827
rect 14133 63771 14219 63827
rect 14275 63771 14361 63827
rect 14417 63771 14503 63827
rect 14559 63771 14645 63827
rect 14701 63771 14787 63827
rect 14843 63771 14853 63827
rect 151 63685 14853 63771
rect 151 63629 161 63685
rect 217 63629 303 63685
rect 359 63629 445 63685
rect 501 63629 587 63685
rect 643 63629 729 63685
rect 785 63629 871 63685
rect 927 63629 1013 63685
rect 1069 63629 1155 63685
rect 1211 63629 1297 63685
rect 1353 63629 1439 63685
rect 1495 63629 1581 63685
rect 1637 63629 1723 63685
rect 1779 63629 1865 63685
rect 1921 63629 2007 63685
rect 2063 63629 2149 63685
rect 2205 63629 2291 63685
rect 2347 63629 2433 63685
rect 2489 63629 2575 63685
rect 2631 63629 2717 63685
rect 2773 63629 2859 63685
rect 2915 63629 3001 63685
rect 3057 63629 3143 63685
rect 3199 63629 3285 63685
rect 3341 63629 3427 63685
rect 3483 63629 3569 63685
rect 3625 63629 3711 63685
rect 3767 63629 3853 63685
rect 3909 63629 3995 63685
rect 4051 63629 4137 63685
rect 4193 63629 4279 63685
rect 4335 63629 4421 63685
rect 4477 63629 4563 63685
rect 4619 63629 4705 63685
rect 4761 63629 4847 63685
rect 4903 63629 4989 63685
rect 5045 63629 5131 63685
rect 5187 63629 5273 63685
rect 5329 63629 5415 63685
rect 5471 63629 5557 63685
rect 5613 63629 5699 63685
rect 5755 63629 5841 63685
rect 5897 63629 5983 63685
rect 6039 63629 6125 63685
rect 6181 63629 6267 63685
rect 6323 63629 6409 63685
rect 6465 63629 6551 63685
rect 6607 63629 6693 63685
rect 6749 63629 6835 63685
rect 6891 63629 6977 63685
rect 7033 63629 7119 63685
rect 7175 63629 7261 63685
rect 7317 63629 7403 63685
rect 7459 63629 7545 63685
rect 7601 63629 7687 63685
rect 7743 63629 7829 63685
rect 7885 63629 7971 63685
rect 8027 63629 8113 63685
rect 8169 63629 8255 63685
rect 8311 63629 8397 63685
rect 8453 63629 8539 63685
rect 8595 63629 8681 63685
rect 8737 63629 8823 63685
rect 8879 63629 8965 63685
rect 9021 63629 9107 63685
rect 9163 63629 9249 63685
rect 9305 63629 9391 63685
rect 9447 63629 9533 63685
rect 9589 63629 9675 63685
rect 9731 63629 9817 63685
rect 9873 63629 9959 63685
rect 10015 63629 10101 63685
rect 10157 63629 10243 63685
rect 10299 63629 10385 63685
rect 10441 63629 10527 63685
rect 10583 63629 10669 63685
rect 10725 63629 10811 63685
rect 10867 63629 10953 63685
rect 11009 63629 11095 63685
rect 11151 63629 11237 63685
rect 11293 63629 11379 63685
rect 11435 63629 11521 63685
rect 11577 63629 11663 63685
rect 11719 63629 11805 63685
rect 11861 63629 11947 63685
rect 12003 63629 12089 63685
rect 12145 63629 12231 63685
rect 12287 63629 12373 63685
rect 12429 63629 12515 63685
rect 12571 63629 12657 63685
rect 12713 63629 12799 63685
rect 12855 63629 12941 63685
rect 12997 63629 13083 63685
rect 13139 63629 13225 63685
rect 13281 63629 13367 63685
rect 13423 63629 13509 63685
rect 13565 63629 13651 63685
rect 13707 63629 13793 63685
rect 13849 63629 13935 63685
rect 13991 63629 14077 63685
rect 14133 63629 14219 63685
rect 14275 63629 14361 63685
rect 14417 63629 14503 63685
rect 14559 63629 14645 63685
rect 14701 63629 14787 63685
rect 14843 63629 14853 63685
rect 151 63619 14853 63629
rect 151 63371 14853 63381
rect 151 63315 161 63371
rect 217 63315 303 63371
rect 359 63315 445 63371
rect 501 63315 587 63371
rect 643 63315 729 63371
rect 785 63315 871 63371
rect 927 63315 1013 63371
rect 1069 63315 1155 63371
rect 1211 63315 1297 63371
rect 1353 63315 1439 63371
rect 1495 63315 1581 63371
rect 1637 63315 1723 63371
rect 1779 63315 1865 63371
rect 1921 63315 2007 63371
rect 2063 63315 2149 63371
rect 2205 63315 2291 63371
rect 2347 63315 2433 63371
rect 2489 63315 2575 63371
rect 2631 63315 2717 63371
rect 2773 63315 2859 63371
rect 2915 63315 3001 63371
rect 3057 63315 3143 63371
rect 3199 63315 3285 63371
rect 3341 63315 3427 63371
rect 3483 63315 3569 63371
rect 3625 63315 3711 63371
rect 3767 63315 3853 63371
rect 3909 63315 3995 63371
rect 4051 63315 4137 63371
rect 4193 63315 4279 63371
rect 4335 63315 4421 63371
rect 4477 63315 4563 63371
rect 4619 63315 4705 63371
rect 4761 63315 4847 63371
rect 4903 63315 4989 63371
rect 5045 63315 5131 63371
rect 5187 63315 5273 63371
rect 5329 63315 5415 63371
rect 5471 63315 5557 63371
rect 5613 63315 5699 63371
rect 5755 63315 5841 63371
rect 5897 63315 5983 63371
rect 6039 63315 6125 63371
rect 6181 63315 6267 63371
rect 6323 63315 6409 63371
rect 6465 63315 6551 63371
rect 6607 63315 6693 63371
rect 6749 63315 6835 63371
rect 6891 63315 6977 63371
rect 7033 63315 7119 63371
rect 7175 63315 7261 63371
rect 7317 63315 7403 63371
rect 7459 63315 7545 63371
rect 7601 63315 7687 63371
rect 7743 63315 7829 63371
rect 7885 63315 7971 63371
rect 8027 63315 8113 63371
rect 8169 63315 8255 63371
rect 8311 63315 8397 63371
rect 8453 63315 8539 63371
rect 8595 63315 8681 63371
rect 8737 63315 8823 63371
rect 8879 63315 8965 63371
rect 9021 63315 9107 63371
rect 9163 63315 9249 63371
rect 9305 63315 9391 63371
rect 9447 63315 9533 63371
rect 9589 63315 9675 63371
rect 9731 63315 9817 63371
rect 9873 63315 9959 63371
rect 10015 63315 10101 63371
rect 10157 63315 10243 63371
rect 10299 63315 10385 63371
rect 10441 63315 10527 63371
rect 10583 63315 10669 63371
rect 10725 63315 10811 63371
rect 10867 63315 10953 63371
rect 11009 63315 11095 63371
rect 11151 63315 11237 63371
rect 11293 63315 11379 63371
rect 11435 63315 11521 63371
rect 11577 63315 11663 63371
rect 11719 63315 11805 63371
rect 11861 63315 11947 63371
rect 12003 63315 12089 63371
rect 12145 63315 12231 63371
rect 12287 63315 12373 63371
rect 12429 63315 12515 63371
rect 12571 63315 12657 63371
rect 12713 63315 12799 63371
rect 12855 63315 12941 63371
rect 12997 63315 13083 63371
rect 13139 63315 13225 63371
rect 13281 63315 13367 63371
rect 13423 63315 13509 63371
rect 13565 63315 13651 63371
rect 13707 63315 13793 63371
rect 13849 63315 13935 63371
rect 13991 63315 14077 63371
rect 14133 63315 14219 63371
rect 14275 63315 14361 63371
rect 14417 63315 14503 63371
rect 14559 63315 14645 63371
rect 14701 63315 14787 63371
rect 14843 63315 14853 63371
rect 151 63229 14853 63315
rect 151 63173 161 63229
rect 217 63173 303 63229
rect 359 63173 445 63229
rect 501 63173 587 63229
rect 643 63173 729 63229
rect 785 63173 871 63229
rect 927 63173 1013 63229
rect 1069 63173 1155 63229
rect 1211 63173 1297 63229
rect 1353 63173 1439 63229
rect 1495 63173 1581 63229
rect 1637 63173 1723 63229
rect 1779 63173 1865 63229
rect 1921 63173 2007 63229
rect 2063 63173 2149 63229
rect 2205 63173 2291 63229
rect 2347 63173 2433 63229
rect 2489 63173 2575 63229
rect 2631 63173 2717 63229
rect 2773 63173 2859 63229
rect 2915 63173 3001 63229
rect 3057 63173 3143 63229
rect 3199 63173 3285 63229
rect 3341 63173 3427 63229
rect 3483 63173 3569 63229
rect 3625 63173 3711 63229
rect 3767 63173 3853 63229
rect 3909 63173 3995 63229
rect 4051 63173 4137 63229
rect 4193 63173 4279 63229
rect 4335 63173 4421 63229
rect 4477 63173 4563 63229
rect 4619 63173 4705 63229
rect 4761 63173 4847 63229
rect 4903 63173 4989 63229
rect 5045 63173 5131 63229
rect 5187 63173 5273 63229
rect 5329 63173 5415 63229
rect 5471 63173 5557 63229
rect 5613 63173 5699 63229
rect 5755 63173 5841 63229
rect 5897 63173 5983 63229
rect 6039 63173 6125 63229
rect 6181 63173 6267 63229
rect 6323 63173 6409 63229
rect 6465 63173 6551 63229
rect 6607 63173 6693 63229
rect 6749 63173 6835 63229
rect 6891 63173 6977 63229
rect 7033 63173 7119 63229
rect 7175 63173 7261 63229
rect 7317 63173 7403 63229
rect 7459 63173 7545 63229
rect 7601 63173 7687 63229
rect 7743 63173 7829 63229
rect 7885 63173 7971 63229
rect 8027 63173 8113 63229
rect 8169 63173 8255 63229
rect 8311 63173 8397 63229
rect 8453 63173 8539 63229
rect 8595 63173 8681 63229
rect 8737 63173 8823 63229
rect 8879 63173 8965 63229
rect 9021 63173 9107 63229
rect 9163 63173 9249 63229
rect 9305 63173 9391 63229
rect 9447 63173 9533 63229
rect 9589 63173 9675 63229
rect 9731 63173 9817 63229
rect 9873 63173 9959 63229
rect 10015 63173 10101 63229
rect 10157 63173 10243 63229
rect 10299 63173 10385 63229
rect 10441 63173 10527 63229
rect 10583 63173 10669 63229
rect 10725 63173 10811 63229
rect 10867 63173 10953 63229
rect 11009 63173 11095 63229
rect 11151 63173 11237 63229
rect 11293 63173 11379 63229
rect 11435 63173 11521 63229
rect 11577 63173 11663 63229
rect 11719 63173 11805 63229
rect 11861 63173 11947 63229
rect 12003 63173 12089 63229
rect 12145 63173 12231 63229
rect 12287 63173 12373 63229
rect 12429 63173 12515 63229
rect 12571 63173 12657 63229
rect 12713 63173 12799 63229
rect 12855 63173 12941 63229
rect 12997 63173 13083 63229
rect 13139 63173 13225 63229
rect 13281 63173 13367 63229
rect 13423 63173 13509 63229
rect 13565 63173 13651 63229
rect 13707 63173 13793 63229
rect 13849 63173 13935 63229
rect 13991 63173 14077 63229
rect 14133 63173 14219 63229
rect 14275 63173 14361 63229
rect 14417 63173 14503 63229
rect 14559 63173 14645 63229
rect 14701 63173 14787 63229
rect 14843 63173 14853 63229
rect 151 63087 14853 63173
rect 151 63031 161 63087
rect 217 63031 303 63087
rect 359 63031 445 63087
rect 501 63031 587 63087
rect 643 63031 729 63087
rect 785 63031 871 63087
rect 927 63031 1013 63087
rect 1069 63031 1155 63087
rect 1211 63031 1297 63087
rect 1353 63031 1439 63087
rect 1495 63031 1581 63087
rect 1637 63031 1723 63087
rect 1779 63031 1865 63087
rect 1921 63031 2007 63087
rect 2063 63031 2149 63087
rect 2205 63031 2291 63087
rect 2347 63031 2433 63087
rect 2489 63031 2575 63087
rect 2631 63031 2717 63087
rect 2773 63031 2859 63087
rect 2915 63031 3001 63087
rect 3057 63031 3143 63087
rect 3199 63031 3285 63087
rect 3341 63031 3427 63087
rect 3483 63031 3569 63087
rect 3625 63031 3711 63087
rect 3767 63031 3853 63087
rect 3909 63031 3995 63087
rect 4051 63031 4137 63087
rect 4193 63031 4279 63087
rect 4335 63031 4421 63087
rect 4477 63031 4563 63087
rect 4619 63031 4705 63087
rect 4761 63031 4847 63087
rect 4903 63031 4989 63087
rect 5045 63031 5131 63087
rect 5187 63031 5273 63087
rect 5329 63031 5415 63087
rect 5471 63031 5557 63087
rect 5613 63031 5699 63087
rect 5755 63031 5841 63087
rect 5897 63031 5983 63087
rect 6039 63031 6125 63087
rect 6181 63031 6267 63087
rect 6323 63031 6409 63087
rect 6465 63031 6551 63087
rect 6607 63031 6693 63087
rect 6749 63031 6835 63087
rect 6891 63031 6977 63087
rect 7033 63031 7119 63087
rect 7175 63031 7261 63087
rect 7317 63031 7403 63087
rect 7459 63031 7545 63087
rect 7601 63031 7687 63087
rect 7743 63031 7829 63087
rect 7885 63031 7971 63087
rect 8027 63031 8113 63087
rect 8169 63031 8255 63087
rect 8311 63031 8397 63087
rect 8453 63031 8539 63087
rect 8595 63031 8681 63087
rect 8737 63031 8823 63087
rect 8879 63031 8965 63087
rect 9021 63031 9107 63087
rect 9163 63031 9249 63087
rect 9305 63031 9391 63087
rect 9447 63031 9533 63087
rect 9589 63031 9675 63087
rect 9731 63031 9817 63087
rect 9873 63031 9959 63087
rect 10015 63031 10101 63087
rect 10157 63031 10243 63087
rect 10299 63031 10385 63087
rect 10441 63031 10527 63087
rect 10583 63031 10669 63087
rect 10725 63031 10811 63087
rect 10867 63031 10953 63087
rect 11009 63031 11095 63087
rect 11151 63031 11237 63087
rect 11293 63031 11379 63087
rect 11435 63031 11521 63087
rect 11577 63031 11663 63087
rect 11719 63031 11805 63087
rect 11861 63031 11947 63087
rect 12003 63031 12089 63087
rect 12145 63031 12231 63087
rect 12287 63031 12373 63087
rect 12429 63031 12515 63087
rect 12571 63031 12657 63087
rect 12713 63031 12799 63087
rect 12855 63031 12941 63087
rect 12997 63031 13083 63087
rect 13139 63031 13225 63087
rect 13281 63031 13367 63087
rect 13423 63031 13509 63087
rect 13565 63031 13651 63087
rect 13707 63031 13793 63087
rect 13849 63031 13935 63087
rect 13991 63031 14077 63087
rect 14133 63031 14219 63087
rect 14275 63031 14361 63087
rect 14417 63031 14503 63087
rect 14559 63031 14645 63087
rect 14701 63031 14787 63087
rect 14843 63031 14853 63087
rect 151 62945 14853 63031
rect 151 62889 161 62945
rect 217 62889 303 62945
rect 359 62889 445 62945
rect 501 62889 587 62945
rect 643 62889 729 62945
rect 785 62889 871 62945
rect 927 62889 1013 62945
rect 1069 62889 1155 62945
rect 1211 62889 1297 62945
rect 1353 62889 1439 62945
rect 1495 62889 1581 62945
rect 1637 62889 1723 62945
rect 1779 62889 1865 62945
rect 1921 62889 2007 62945
rect 2063 62889 2149 62945
rect 2205 62889 2291 62945
rect 2347 62889 2433 62945
rect 2489 62889 2575 62945
rect 2631 62889 2717 62945
rect 2773 62889 2859 62945
rect 2915 62889 3001 62945
rect 3057 62889 3143 62945
rect 3199 62889 3285 62945
rect 3341 62889 3427 62945
rect 3483 62889 3569 62945
rect 3625 62889 3711 62945
rect 3767 62889 3853 62945
rect 3909 62889 3995 62945
rect 4051 62889 4137 62945
rect 4193 62889 4279 62945
rect 4335 62889 4421 62945
rect 4477 62889 4563 62945
rect 4619 62889 4705 62945
rect 4761 62889 4847 62945
rect 4903 62889 4989 62945
rect 5045 62889 5131 62945
rect 5187 62889 5273 62945
rect 5329 62889 5415 62945
rect 5471 62889 5557 62945
rect 5613 62889 5699 62945
rect 5755 62889 5841 62945
rect 5897 62889 5983 62945
rect 6039 62889 6125 62945
rect 6181 62889 6267 62945
rect 6323 62889 6409 62945
rect 6465 62889 6551 62945
rect 6607 62889 6693 62945
rect 6749 62889 6835 62945
rect 6891 62889 6977 62945
rect 7033 62889 7119 62945
rect 7175 62889 7261 62945
rect 7317 62889 7403 62945
rect 7459 62889 7545 62945
rect 7601 62889 7687 62945
rect 7743 62889 7829 62945
rect 7885 62889 7971 62945
rect 8027 62889 8113 62945
rect 8169 62889 8255 62945
rect 8311 62889 8397 62945
rect 8453 62889 8539 62945
rect 8595 62889 8681 62945
rect 8737 62889 8823 62945
rect 8879 62889 8965 62945
rect 9021 62889 9107 62945
rect 9163 62889 9249 62945
rect 9305 62889 9391 62945
rect 9447 62889 9533 62945
rect 9589 62889 9675 62945
rect 9731 62889 9817 62945
rect 9873 62889 9959 62945
rect 10015 62889 10101 62945
rect 10157 62889 10243 62945
rect 10299 62889 10385 62945
rect 10441 62889 10527 62945
rect 10583 62889 10669 62945
rect 10725 62889 10811 62945
rect 10867 62889 10953 62945
rect 11009 62889 11095 62945
rect 11151 62889 11237 62945
rect 11293 62889 11379 62945
rect 11435 62889 11521 62945
rect 11577 62889 11663 62945
rect 11719 62889 11805 62945
rect 11861 62889 11947 62945
rect 12003 62889 12089 62945
rect 12145 62889 12231 62945
rect 12287 62889 12373 62945
rect 12429 62889 12515 62945
rect 12571 62889 12657 62945
rect 12713 62889 12799 62945
rect 12855 62889 12941 62945
rect 12997 62889 13083 62945
rect 13139 62889 13225 62945
rect 13281 62889 13367 62945
rect 13423 62889 13509 62945
rect 13565 62889 13651 62945
rect 13707 62889 13793 62945
rect 13849 62889 13935 62945
rect 13991 62889 14077 62945
rect 14133 62889 14219 62945
rect 14275 62889 14361 62945
rect 14417 62889 14503 62945
rect 14559 62889 14645 62945
rect 14701 62889 14787 62945
rect 14843 62889 14853 62945
rect 151 62803 14853 62889
rect 151 62747 161 62803
rect 217 62747 303 62803
rect 359 62747 445 62803
rect 501 62747 587 62803
rect 643 62747 729 62803
rect 785 62747 871 62803
rect 927 62747 1013 62803
rect 1069 62747 1155 62803
rect 1211 62747 1297 62803
rect 1353 62747 1439 62803
rect 1495 62747 1581 62803
rect 1637 62747 1723 62803
rect 1779 62747 1865 62803
rect 1921 62747 2007 62803
rect 2063 62747 2149 62803
rect 2205 62747 2291 62803
rect 2347 62747 2433 62803
rect 2489 62747 2575 62803
rect 2631 62747 2717 62803
rect 2773 62747 2859 62803
rect 2915 62747 3001 62803
rect 3057 62747 3143 62803
rect 3199 62747 3285 62803
rect 3341 62747 3427 62803
rect 3483 62747 3569 62803
rect 3625 62747 3711 62803
rect 3767 62747 3853 62803
rect 3909 62747 3995 62803
rect 4051 62747 4137 62803
rect 4193 62747 4279 62803
rect 4335 62747 4421 62803
rect 4477 62747 4563 62803
rect 4619 62747 4705 62803
rect 4761 62747 4847 62803
rect 4903 62747 4989 62803
rect 5045 62747 5131 62803
rect 5187 62747 5273 62803
rect 5329 62747 5415 62803
rect 5471 62747 5557 62803
rect 5613 62747 5699 62803
rect 5755 62747 5841 62803
rect 5897 62747 5983 62803
rect 6039 62747 6125 62803
rect 6181 62747 6267 62803
rect 6323 62747 6409 62803
rect 6465 62747 6551 62803
rect 6607 62747 6693 62803
rect 6749 62747 6835 62803
rect 6891 62747 6977 62803
rect 7033 62747 7119 62803
rect 7175 62747 7261 62803
rect 7317 62747 7403 62803
rect 7459 62747 7545 62803
rect 7601 62747 7687 62803
rect 7743 62747 7829 62803
rect 7885 62747 7971 62803
rect 8027 62747 8113 62803
rect 8169 62747 8255 62803
rect 8311 62747 8397 62803
rect 8453 62747 8539 62803
rect 8595 62747 8681 62803
rect 8737 62747 8823 62803
rect 8879 62747 8965 62803
rect 9021 62747 9107 62803
rect 9163 62747 9249 62803
rect 9305 62747 9391 62803
rect 9447 62747 9533 62803
rect 9589 62747 9675 62803
rect 9731 62747 9817 62803
rect 9873 62747 9959 62803
rect 10015 62747 10101 62803
rect 10157 62747 10243 62803
rect 10299 62747 10385 62803
rect 10441 62747 10527 62803
rect 10583 62747 10669 62803
rect 10725 62747 10811 62803
rect 10867 62747 10953 62803
rect 11009 62747 11095 62803
rect 11151 62747 11237 62803
rect 11293 62747 11379 62803
rect 11435 62747 11521 62803
rect 11577 62747 11663 62803
rect 11719 62747 11805 62803
rect 11861 62747 11947 62803
rect 12003 62747 12089 62803
rect 12145 62747 12231 62803
rect 12287 62747 12373 62803
rect 12429 62747 12515 62803
rect 12571 62747 12657 62803
rect 12713 62747 12799 62803
rect 12855 62747 12941 62803
rect 12997 62747 13083 62803
rect 13139 62747 13225 62803
rect 13281 62747 13367 62803
rect 13423 62747 13509 62803
rect 13565 62747 13651 62803
rect 13707 62747 13793 62803
rect 13849 62747 13935 62803
rect 13991 62747 14077 62803
rect 14133 62747 14219 62803
rect 14275 62747 14361 62803
rect 14417 62747 14503 62803
rect 14559 62747 14645 62803
rect 14701 62747 14787 62803
rect 14843 62747 14853 62803
rect 151 62661 14853 62747
rect 151 62605 161 62661
rect 217 62605 303 62661
rect 359 62605 445 62661
rect 501 62605 587 62661
rect 643 62605 729 62661
rect 785 62605 871 62661
rect 927 62605 1013 62661
rect 1069 62605 1155 62661
rect 1211 62605 1297 62661
rect 1353 62605 1439 62661
rect 1495 62605 1581 62661
rect 1637 62605 1723 62661
rect 1779 62605 1865 62661
rect 1921 62605 2007 62661
rect 2063 62605 2149 62661
rect 2205 62605 2291 62661
rect 2347 62605 2433 62661
rect 2489 62605 2575 62661
rect 2631 62605 2717 62661
rect 2773 62605 2859 62661
rect 2915 62605 3001 62661
rect 3057 62605 3143 62661
rect 3199 62605 3285 62661
rect 3341 62605 3427 62661
rect 3483 62605 3569 62661
rect 3625 62605 3711 62661
rect 3767 62605 3853 62661
rect 3909 62605 3995 62661
rect 4051 62605 4137 62661
rect 4193 62605 4279 62661
rect 4335 62605 4421 62661
rect 4477 62605 4563 62661
rect 4619 62605 4705 62661
rect 4761 62605 4847 62661
rect 4903 62605 4989 62661
rect 5045 62605 5131 62661
rect 5187 62605 5273 62661
rect 5329 62605 5415 62661
rect 5471 62605 5557 62661
rect 5613 62605 5699 62661
rect 5755 62605 5841 62661
rect 5897 62605 5983 62661
rect 6039 62605 6125 62661
rect 6181 62605 6267 62661
rect 6323 62605 6409 62661
rect 6465 62605 6551 62661
rect 6607 62605 6693 62661
rect 6749 62605 6835 62661
rect 6891 62605 6977 62661
rect 7033 62605 7119 62661
rect 7175 62605 7261 62661
rect 7317 62605 7403 62661
rect 7459 62605 7545 62661
rect 7601 62605 7687 62661
rect 7743 62605 7829 62661
rect 7885 62605 7971 62661
rect 8027 62605 8113 62661
rect 8169 62605 8255 62661
rect 8311 62605 8397 62661
rect 8453 62605 8539 62661
rect 8595 62605 8681 62661
rect 8737 62605 8823 62661
rect 8879 62605 8965 62661
rect 9021 62605 9107 62661
rect 9163 62605 9249 62661
rect 9305 62605 9391 62661
rect 9447 62605 9533 62661
rect 9589 62605 9675 62661
rect 9731 62605 9817 62661
rect 9873 62605 9959 62661
rect 10015 62605 10101 62661
rect 10157 62605 10243 62661
rect 10299 62605 10385 62661
rect 10441 62605 10527 62661
rect 10583 62605 10669 62661
rect 10725 62605 10811 62661
rect 10867 62605 10953 62661
rect 11009 62605 11095 62661
rect 11151 62605 11237 62661
rect 11293 62605 11379 62661
rect 11435 62605 11521 62661
rect 11577 62605 11663 62661
rect 11719 62605 11805 62661
rect 11861 62605 11947 62661
rect 12003 62605 12089 62661
rect 12145 62605 12231 62661
rect 12287 62605 12373 62661
rect 12429 62605 12515 62661
rect 12571 62605 12657 62661
rect 12713 62605 12799 62661
rect 12855 62605 12941 62661
rect 12997 62605 13083 62661
rect 13139 62605 13225 62661
rect 13281 62605 13367 62661
rect 13423 62605 13509 62661
rect 13565 62605 13651 62661
rect 13707 62605 13793 62661
rect 13849 62605 13935 62661
rect 13991 62605 14077 62661
rect 14133 62605 14219 62661
rect 14275 62605 14361 62661
rect 14417 62605 14503 62661
rect 14559 62605 14645 62661
rect 14701 62605 14787 62661
rect 14843 62605 14853 62661
rect 151 62519 14853 62605
rect 151 62463 161 62519
rect 217 62463 303 62519
rect 359 62463 445 62519
rect 501 62463 587 62519
rect 643 62463 729 62519
rect 785 62463 871 62519
rect 927 62463 1013 62519
rect 1069 62463 1155 62519
rect 1211 62463 1297 62519
rect 1353 62463 1439 62519
rect 1495 62463 1581 62519
rect 1637 62463 1723 62519
rect 1779 62463 1865 62519
rect 1921 62463 2007 62519
rect 2063 62463 2149 62519
rect 2205 62463 2291 62519
rect 2347 62463 2433 62519
rect 2489 62463 2575 62519
rect 2631 62463 2717 62519
rect 2773 62463 2859 62519
rect 2915 62463 3001 62519
rect 3057 62463 3143 62519
rect 3199 62463 3285 62519
rect 3341 62463 3427 62519
rect 3483 62463 3569 62519
rect 3625 62463 3711 62519
rect 3767 62463 3853 62519
rect 3909 62463 3995 62519
rect 4051 62463 4137 62519
rect 4193 62463 4279 62519
rect 4335 62463 4421 62519
rect 4477 62463 4563 62519
rect 4619 62463 4705 62519
rect 4761 62463 4847 62519
rect 4903 62463 4989 62519
rect 5045 62463 5131 62519
rect 5187 62463 5273 62519
rect 5329 62463 5415 62519
rect 5471 62463 5557 62519
rect 5613 62463 5699 62519
rect 5755 62463 5841 62519
rect 5897 62463 5983 62519
rect 6039 62463 6125 62519
rect 6181 62463 6267 62519
rect 6323 62463 6409 62519
rect 6465 62463 6551 62519
rect 6607 62463 6693 62519
rect 6749 62463 6835 62519
rect 6891 62463 6977 62519
rect 7033 62463 7119 62519
rect 7175 62463 7261 62519
rect 7317 62463 7403 62519
rect 7459 62463 7545 62519
rect 7601 62463 7687 62519
rect 7743 62463 7829 62519
rect 7885 62463 7971 62519
rect 8027 62463 8113 62519
rect 8169 62463 8255 62519
rect 8311 62463 8397 62519
rect 8453 62463 8539 62519
rect 8595 62463 8681 62519
rect 8737 62463 8823 62519
rect 8879 62463 8965 62519
rect 9021 62463 9107 62519
rect 9163 62463 9249 62519
rect 9305 62463 9391 62519
rect 9447 62463 9533 62519
rect 9589 62463 9675 62519
rect 9731 62463 9817 62519
rect 9873 62463 9959 62519
rect 10015 62463 10101 62519
rect 10157 62463 10243 62519
rect 10299 62463 10385 62519
rect 10441 62463 10527 62519
rect 10583 62463 10669 62519
rect 10725 62463 10811 62519
rect 10867 62463 10953 62519
rect 11009 62463 11095 62519
rect 11151 62463 11237 62519
rect 11293 62463 11379 62519
rect 11435 62463 11521 62519
rect 11577 62463 11663 62519
rect 11719 62463 11805 62519
rect 11861 62463 11947 62519
rect 12003 62463 12089 62519
rect 12145 62463 12231 62519
rect 12287 62463 12373 62519
rect 12429 62463 12515 62519
rect 12571 62463 12657 62519
rect 12713 62463 12799 62519
rect 12855 62463 12941 62519
rect 12997 62463 13083 62519
rect 13139 62463 13225 62519
rect 13281 62463 13367 62519
rect 13423 62463 13509 62519
rect 13565 62463 13651 62519
rect 13707 62463 13793 62519
rect 13849 62463 13935 62519
rect 13991 62463 14077 62519
rect 14133 62463 14219 62519
rect 14275 62463 14361 62519
rect 14417 62463 14503 62519
rect 14559 62463 14645 62519
rect 14701 62463 14787 62519
rect 14843 62463 14853 62519
rect 151 62377 14853 62463
rect 151 62321 161 62377
rect 217 62321 303 62377
rect 359 62321 445 62377
rect 501 62321 587 62377
rect 643 62321 729 62377
rect 785 62321 871 62377
rect 927 62321 1013 62377
rect 1069 62321 1155 62377
rect 1211 62321 1297 62377
rect 1353 62321 1439 62377
rect 1495 62321 1581 62377
rect 1637 62321 1723 62377
rect 1779 62321 1865 62377
rect 1921 62321 2007 62377
rect 2063 62321 2149 62377
rect 2205 62321 2291 62377
rect 2347 62321 2433 62377
rect 2489 62321 2575 62377
rect 2631 62321 2717 62377
rect 2773 62321 2859 62377
rect 2915 62321 3001 62377
rect 3057 62321 3143 62377
rect 3199 62321 3285 62377
rect 3341 62321 3427 62377
rect 3483 62321 3569 62377
rect 3625 62321 3711 62377
rect 3767 62321 3853 62377
rect 3909 62321 3995 62377
rect 4051 62321 4137 62377
rect 4193 62321 4279 62377
rect 4335 62321 4421 62377
rect 4477 62321 4563 62377
rect 4619 62321 4705 62377
rect 4761 62321 4847 62377
rect 4903 62321 4989 62377
rect 5045 62321 5131 62377
rect 5187 62321 5273 62377
rect 5329 62321 5415 62377
rect 5471 62321 5557 62377
rect 5613 62321 5699 62377
rect 5755 62321 5841 62377
rect 5897 62321 5983 62377
rect 6039 62321 6125 62377
rect 6181 62321 6267 62377
rect 6323 62321 6409 62377
rect 6465 62321 6551 62377
rect 6607 62321 6693 62377
rect 6749 62321 6835 62377
rect 6891 62321 6977 62377
rect 7033 62321 7119 62377
rect 7175 62321 7261 62377
rect 7317 62321 7403 62377
rect 7459 62321 7545 62377
rect 7601 62321 7687 62377
rect 7743 62321 7829 62377
rect 7885 62321 7971 62377
rect 8027 62321 8113 62377
rect 8169 62321 8255 62377
rect 8311 62321 8397 62377
rect 8453 62321 8539 62377
rect 8595 62321 8681 62377
rect 8737 62321 8823 62377
rect 8879 62321 8965 62377
rect 9021 62321 9107 62377
rect 9163 62321 9249 62377
rect 9305 62321 9391 62377
rect 9447 62321 9533 62377
rect 9589 62321 9675 62377
rect 9731 62321 9817 62377
rect 9873 62321 9959 62377
rect 10015 62321 10101 62377
rect 10157 62321 10243 62377
rect 10299 62321 10385 62377
rect 10441 62321 10527 62377
rect 10583 62321 10669 62377
rect 10725 62321 10811 62377
rect 10867 62321 10953 62377
rect 11009 62321 11095 62377
rect 11151 62321 11237 62377
rect 11293 62321 11379 62377
rect 11435 62321 11521 62377
rect 11577 62321 11663 62377
rect 11719 62321 11805 62377
rect 11861 62321 11947 62377
rect 12003 62321 12089 62377
rect 12145 62321 12231 62377
rect 12287 62321 12373 62377
rect 12429 62321 12515 62377
rect 12571 62321 12657 62377
rect 12713 62321 12799 62377
rect 12855 62321 12941 62377
rect 12997 62321 13083 62377
rect 13139 62321 13225 62377
rect 13281 62321 13367 62377
rect 13423 62321 13509 62377
rect 13565 62321 13651 62377
rect 13707 62321 13793 62377
rect 13849 62321 13935 62377
rect 13991 62321 14077 62377
rect 14133 62321 14219 62377
rect 14275 62321 14361 62377
rect 14417 62321 14503 62377
rect 14559 62321 14645 62377
rect 14701 62321 14787 62377
rect 14843 62321 14853 62377
rect 151 62235 14853 62321
rect 151 62179 161 62235
rect 217 62179 303 62235
rect 359 62179 445 62235
rect 501 62179 587 62235
rect 643 62179 729 62235
rect 785 62179 871 62235
rect 927 62179 1013 62235
rect 1069 62179 1155 62235
rect 1211 62179 1297 62235
rect 1353 62179 1439 62235
rect 1495 62179 1581 62235
rect 1637 62179 1723 62235
rect 1779 62179 1865 62235
rect 1921 62179 2007 62235
rect 2063 62179 2149 62235
rect 2205 62179 2291 62235
rect 2347 62179 2433 62235
rect 2489 62179 2575 62235
rect 2631 62179 2717 62235
rect 2773 62179 2859 62235
rect 2915 62179 3001 62235
rect 3057 62179 3143 62235
rect 3199 62179 3285 62235
rect 3341 62179 3427 62235
rect 3483 62179 3569 62235
rect 3625 62179 3711 62235
rect 3767 62179 3853 62235
rect 3909 62179 3995 62235
rect 4051 62179 4137 62235
rect 4193 62179 4279 62235
rect 4335 62179 4421 62235
rect 4477 62179 4563 62235
rect 4619 62179 4705 62235
rect 4761 62179 4847 62235
rect 4903 62179 4989 62235
rect 5045 62179 5131 62235
rect 5187 62179 5273 62235
rect 5329 62179 5415 62235
rect 5471 62179 5557 62235
rect 5613 62179 5699 62235
rect 5755 62179 5841 62235
rect 5897 62179 5983 62235
rect 6039 62179 6125 62235
rect 6181 62179 6267 62235
rect 6323 62179 6409 62235
rect 6465 62179 6551 62235
rect 6607 62179 6693 62235
rect 6749 62179 6835 62235
rect 6891 62179 6977 62235
rect 7033 62179 7119 62235
rect 7175 62179 7261 62235
rect 7317 62179 7403 62235
rect 7459 62179 7545 62235
rect 7601 62179 7687 62235
rect 7743 62179 7829 62235
rect 7885 62179 7971 62235
rect 8027 62179 8113 62235
rect 8169 62179 8255 62235
rect 8311 62179 8397 62235
rect 8453 62179 8539 62235
rect 8595 62179 8681 62235
rect 8737 62179 8823 62235
rect 8879 62179 8965 62235
rect 9021 62179 9107 62235
rect 9163 62179 9249 62235
rect 9305 62179 9391 62235
rect 9447 62179 9533 62235
rect 9589 62179 9675 62235
rect 9731 62179 9817 62235
rect 9873 62179 9959 62235
rect 10015 62179 10101 62235
rect 10157 62179 10243 62235
rect 10299 62179 10385 62235
rect 10441 62179 10527 62235
rect 10583 62179 10669 62235
rect 10725 62179 10811 62235
rect 10867 62179 10953 62235
rect 11009 62179 11095 62235
rect 11151 62179 11237 62235
rect 11293 62179 11379 62235
rect 11435 62179 11521 62235
rect 11577 62179 11663 62235
rect 11719 62179 11805 62235
rect 11861 62179 11947 62235
rect 12003 62179 12089 62235
rect 12145 62179 12231 62235
rect 12287 62179 12373 62235
rect 12429 62179 12515 62235
rect 12571 62179 12657 62235
rect 12713 62179 12799 62235
rect 12855 62179 12941 62235
rect 12997 62179 13083 62235
rect 13139 62179 13225 62235
rect 13281 62179 13367 62235
rect 13423 62179 13509 62235
rect 13565 62179 13651 62235
rect 13707 62179 13793 62235
rect 13849 62179 13935 62235
rect 13991 62179 14077 62235
rect 14133 62179 14219 62235
rect 14275 62179 14361 62235
rect 14417 62179 14503 62235
rect 14559 62179 14645 62235
rect 14701 62179 14787 62235
rect 14843 62179 14853 62235
rect 151 62093 14853 62179
rect 151 62037 161 62093
rect 217 62037 303 62093
rect 359 62037 445 62093
rect 501 62037 587 62093
rect 643 62037 729 62093
rect 785 62037 871 62093
rect 927 62037 1013 62093
rect 1069 62037 1155 62093
rect 1211 62037 1297 62093
rect 1353 62037 1439 62093
rect 1495 62037 1581 62093
rect 1637 62037 1723 62093
rect 1779 62037 1865 62093
rect 1921 62037 2007 62093
rect 2063 62037 2149 62093
rect 2205 62037 2291 62093
rect 2347 62037 2433 62093
rect 2489 62037 2575 62093
rect 2631 62037 2717 62093
rect 2773 62037 2859 62093
rect 2915 62037 3001 62093
rect 3057 62037 3143 62093
rect 3199 62037 3285 62093
rect 3341 62037 3427 62093
rect 3483 62037 3569 62093
rect 3625 62037 3711 62093
rect 3767 62037 3853 62093
rect 3909 62037 3995 62093
rect 4051 62037 4137 62093
rect 4193 62037 4279 62093
rect 4335 62037 4421 62093
rect 4477 62037 4563 62093
rect 4619 62037 4705 62093
rect 4761 62037 4847 62093
rect 4903 62037 4989 62093
rect 5045 62037 5131 62093
rect 5187 62037 5273 62093
rect 5329 62037 5415 62093
rect 5471 62037 5557 62093
rect 5613 62037 5699 62093
rect 5755 62037 5841 62093
rect 5897 62037 5983 62093
rect 6039 62037 6125 62093
rect 6181 62037 6267 62093
rect 6323 62037 6409 62093
rect 6465 62037 6551 62093
rect 6607 62037 6693 62093
rect 6749 62037 6835 62093
rect 6891 62037 6977 62093
rect 7033 62037 7119 62093
rect 7175 62037 7261 62093
rect 7317 62037 7403 62093
rect 7459 62037 7545 62093
rect 7601 62037 7687 62093
rect 7743 62037 7829 62093
rect 7885 62037 7971 62093
rect 8027 62037 8113 62093
rect 8169 62037 8255 62093
rect 8311 62037 8397 62093
rect 8453 62037 8539 62093
rect 8595 62037 8681 62093
rect 8737 62037 8823 62093
rect 8879 62037 8965 62093
rect 9021 62037 9107 62093
rect 9163 62037 9249 62093
rect 9305 62037 9391 62093
rect 9447 62037 9533 62093
rect 9589 62037 9675 62093
rect 9731 62037 9817 62093
rect 9873 62037 9959 62093
rect 10015 62037 10101 62093
rect 10157 62037 10243 62093
rect 10299 62037 10385 62093
rect 10441 62037 10527 62093
rect 10583 62037 10669 62093
rect 10725 62037 10811 62093
rect 10867 62037 10953 62093
rect 11009 62037 11095 62093
rect 11151 62037 11237 62093
rect 11293 62037 11379 62093
rect 11435 62037 11521 62093
rect 11577 62037 11663 62093
rect 11719 62037 11805 62093
rect 11861 62037 11947 62093
rect 12003 62037 12089 62093
rect 12145 62037 12231 62093
rect 12287 62037 12373 62093
rect 12429 62037 12515 62093
rect 12571 62037 12657 62093
rect 12713 62037 12799 62093
rect 12855 62037 12941 62093
rect 12997 62037 13083 62093
rect 13139 62037 13225 62093
rect 13281 62037 13367 62093
rect 13423 62037 13509 62093
rect 13565 62037 13651 62093
rect 13707 62037 13793 62093
rect 13849 62037 13935 62093
rect 13991 62037 14077 62093
rect 14133 62037 14219 62093
rect 14275 62037 14361 62093
rect 14417 62037 14503 62093
rect 14559 62037 14645 62093
rect 14701 62037 14787 62093
rect 14843 62037 14853 62093
rect 151 62027 14853 62037
rect 151 61763 14853 61773
rect 151 61707 161 61763
rect 217 61707 303 61763
rect 359 61707 445 61763
rect 501 61707 587 61763
rect 643 61707 729 61763
rect 785 61707 871 61763
rect 927 61707 1013 61763
rect 1069 61707 1155 61763
rect 1211 61707 1297 61763
rect 1353 61707 1439 61763
rect 1495 61707 1581 61763
rect 1637 61707 1723 61763
rect 1779 61707 1865 61763
rect 1921 61707 2007 61763
rect 2063 61707 2149 61763
rect 2205 61707 2291 61763
rect 2347 61707 2433 61763
rect 2489 61707 2575 61763
rect 2631 61707 2717 61763
rect 2773 61707 2859 61763
rect 2915 61707 3001 61763
rect 3057 61707 3143 61763
rect 3199 61707 3285 61763
rect 3341 61707 3427 61763
rect 3483 61707 3569 61763
rect 3625 61707 3711 61763
rect 3767 61707 3853 61763
rect 3909 61707 3995 61763
rect 4051 61707 4137 61763
rect 4193 61707 4279 61763
rect 4335 61707 4421 61763
rect 4477 61707 4563 61763
rect 4619 61707 4705 61763
rect 4761 61707 4847 61763
rect 4903 61707 4989 61763
rect 5045 61707 5131 61763
rect 5187 61707 5273 61763
rect 5329 61707 5415 61763
rect 5471 61707 5557 61763
rect 5613 61707 5699 61763
rect 5755 61707 5841 61763
rect 5897 61707 5983 61763
rect 6039 61707 6125 61763
rect 6181 61707 6267 61763
rect 6323 61707 6409 61763
rect 6465 61707 6551 61763
rect 6607 61707 6693 61763
rect 6749 61707 6835 61763
rect 6891 61707 6977 61763
rect 7033 61707 7119 61763
rect 7175 61707 7261 61763
rect 7317 61707 7403 61763
rect 7459 61707 7545 61763
rect 7601 61707 7687 61763
rect 7743 61707 7829 61763
rect 7885 61707 7971 61763
rect 8027 61707 8113 61763
rect 8169 61707 8255 61763
rect 8311 61707 8397 61763
rect 8453 61707 8539 61763
rect 8595 61707 8681 61763
rect 8737 61707 8823 61763
rect 8879 61707 8965 61763
rect 9021 61707 9107 61763
rect 9163 61707 9249 61763
rect 9305 61707 9391 61763
rect 9447 61707 9533 61763
rect 9589 61707 9675 61763
rect 9731 61707 9817 61763
rect 9873 61707 9959 61763
rect 10015 61707 10101 61763
rect 10157 61707 10243 61763
rect 10299 61707 10385 61763
rect 10441 61707 10527 61763
rect 10583 61707 10669 61763
rect 10725 61707 10811 61763
rect 10867 61707 10953 61763
rect 11009 61707 11095 61763
rect 11151 61707 11237 61763
rect 11293 61707 11379 61763
rect 11435 61707 11521 61763
rect 11577 61707 11663 61763
rect 11719 61707 11805 61763
rect 11861 61707 11947 61763
rect 12003 61707 12089 61763
rect 12145 61707 12231 61763
rect 12287 61707 12373 61763
rect 12429 61707 12515 61763
rect 12571 61707 12657 61763
rect 12713 61707 12799 61763
rect 12855 61707 12941 61763
rect 12997 61707 13083 61763
rect 13139 61707 13225 61763
rect 13281 61707 13367 61763
rect 13423 61707 13509 61763
rect 13565 61707 13651 61763
rect 13707 61707 13793 61763
rect 13849 61707 13935 61763
rect 13991 61707 14077 61763
rect 14133 61707 14219 61763
rect 14275 61707 14361 61763
rect 14417 61707 14503 61763
rect 14559 61707 14645 61763
rect 14701 61707 14787 61763
rect 14843 61707 14853 61763
rect 151 61621 14853 61707
rect 151 61565 161 61621
rect 217 61565 303 61621
rect 359 61565 445 61621
rect 501 61565 587 61621
rect 643 61565 729 61621
rect 785 61565 871 61621
rect 927 61565 1013 61621
rect 1069 61565 1155 61621
rect 1211 61565 1297 61621
rect 1353 61565 1439 61621
rect 1495 61565 1581 61621
rect 1637 61565 1723 61621
rect 1779 61565 1865 61621
rect 1921 61565 2007 61621
rect 2063 61565 2149 61621
rect 2205 61565 2291 61621
rect 2347 61565 2433 61621
rect 2489 61565 2575 61621
rect 2631 61565 2717 61621
rect 2773 61565 2859 61621
rect 2915 61565 3001 61621
rect 3057 61565 3143 61621
rect 3199 61565 3285 61621
rect 3341 61565 3427 61621
rect 3483 61565 3569 61621
rect 3625 61565 3711 61621
rect 3767 61565 3853 61621
rect 3909 61565 3995 61621
rect 4051 61565 4137 61621
rect 4193 61565 4279 61621
rect 4335 61565 4421 61621
rect 4477 61565 4563 61621
rect 4619 61565 4705 61621
rect 4761 61565 4847 61621
rect 4903 61565 4989 61621
rect 5045 61565 5131 61621
rect 5187 61565 5273 61621
rect 5329 61565 5415 61621
rect 5471 61565 5557 61621
rect 5613 61565 5699 61621
rect 5755 61565 5841 61621
rect 5897 61565 5983 61621
rect 6039 61565 6125 61621
rect 6181 61565 6267 61621
rect 6323 61565 6409 61621
rect 6465 61565 6551 61621
rect 6607 61565 6693 61621
rect 6749 61565 6835 61621
rect 6891 61565 6977 61621
rect 7033 61565 7119 61621
rect 7175 61565 7261 61621
rect 7317 61565 7403 61621
rect 7459 61565 7545 61621
rect 7601 61565 7687 61621
rect 7743 61565 7829 61621
rect 7885 61565 7971 61621
rect 8027 61565 8113 61621
rect 8169 61565 8255 61621
rect 8311 61565 8397 61621
rect 8453 61565 8539 61621
rect 8595 61565 8681 61621
rect 8737 61565 8823 61621
rect 8879 61565 8965 61621
rect 9021 61565 9107 61621
rect 9163 61565 9249 61621
rect 9305 61565 9391 61621
rect 9447 61565 9533 61621
rect 9589 61565 9675 61621
rect 9731 61565 9817 61621
rect 9873 61565 9959 61621
rect 10015 61565 10101 61621
rect 10157 61565 10243 61621
rect 10299 61565 10385 61621
rect 10441 61565 10527 61621
rect 10583 61565 10669 61621
rect 10725 61565 10811 61621
rect 10867 61565 10953 61621
rect 11009 61565 11095 61621
rect 11151 61565 11237 61621
rect 11293 61565 11379 61621
rect 11435 61565 11521 61621
rect 11577 61565 11663 61621
rect 11719 61565 11805 61621
rect 11861 61565 11947 61621
rect 12003 61565 12089 61621
rect 12145 61565 12231 61621
rect 12287 61565 12373 61621
rect 12429 61565 12515 61621
rect 12571 61565 12657 61621
rect 12713 61565 12799 61621
rect 12855 61565 12941 61621
rect 12997 61565 13083 61621
rect 13139 61565 13225 61621
rect 13281 61565 13367 61621
rect 13423 61565 13509 61621
rect 13565 61565 13651 61621
rect 13707 61565 13793 61621
rect 13849 61565 13935 61621
rect 13991 61565 14077 61621
rect 14133 61565 14219 61621
rect 14275 61565 14361 61621
rect 14417 61565 14503 61621
rect 14559 61565 14645 61621
rect 14701 61565 14787 61621
rect 14843 61565 14853 61621
rect 151 61479 14853 61565
rect 151 61423 161 61479
rect 217 61423 303 61479
rect 359 61423 445 61479
rect 501 61423 587 61479
rect 643 61423 729 61479
rect 785 61423 871 61479
rect 927 61423 1013 61479
rect 1069 61423 1155 61479
rect 1211 61423 1297 61479
rect 1353 61423 1439 61479
rect 1495 61423 1581 61479
rect 1637 61423 1723 61479
rect 1779 61423 1865 61479
rect 1921 61423 2007 61479
rect 2063 61423 2149 61479
rect 2205 61423 2291 61479
rect 2347 61423 2433 61479
rect 2489 61423 2575 61479
rect 2631 61423 2717 61479
rect 2773 61423 2859 61479
rect 2915 61423 3001 61479
rect 3057 61423 3143 61479
rect 3199 61423 3285 61479
rect 3341 61423 3427 61479
rect 3483 61423 3569 61479
rect 3625 61423 3711 61479
rect 3767 61423 3853 61479
rect 3909 61423 3995 61479
rect 4051 61423 4137 61479
rect 4193 61423 4279 61479
rect 4335 61423 4421 61479
rect 4477 61423 4563 61479
rect 4619 61423 4705 61479
rect 4761 61423 4847 61479
rect 4903 61423 4989 61479
rect 5045 61423 5131 61479
rect 5187 61423 5273 61479
rect 5329 61423 5415 61479
rect 5471 61423 5557 61479
rect 5613 61423 5699 61479
rect 5755 61423 5841 61479
rect 5897 61423 5983 61479
rect 6039 61423 6125 61479
rect 6181 61423 6267 61479
rect 6323 61423 6409 61479
rect 6465 61423 6551 61479
rect 6607 61423 6693 61479
rect 6749 61423 6835 61479
rect 6891 61423 6977 61479
rect 7033 61423 7119 61479
rect 7175 61423 7261 61479
rect 7317 61423 7403 61479
rect 7459 61423 7545 61479
rect 7601 61423 7687 61479
rect 7743 61423 7829 61479
rect 7885 61423 7971 61479
rect 8027 61423 8113 61479
rect 8169 61423 8255 61479
rect 8311 61423 8397 61479
rect 8453 61423 8539 61479
rect 8595 61423 8681 61479
rect 8737 61423 8823 61479
rect 8879 61423 8965 61479
rect 9021 61423 9107 61479
rect 9163 61423 9249 61479
rect 9305 61423 9391 61479
rect 9447 61423 9533 61479
rect 9589 61423 9675 61479
rect 9731 61423 9817 61479
rect 9873 61423 9959 61479
rect 10015 61423 10101 61479
rect 10157 61423 10243 61479
rect 10299 61423 10385 61479
rect 10441 61423 10527 61479
rect 10583 61423 10669 61479
rect 10725 61423 10811 61479
rect 10867 61423 10953 61479
rect 11009 61423 11095 61479
rect 11151 61423 11237 61479
rect 11293 61423 11379 61479
rect 11435 61423 11521 61479
rect 11577 61423 11663 61479
rect 11719 61423 11805 61479
rect 11861 61423 11947 61479
rect 12003 61423 12089 61479
rect 12145 61423 12231 61479
rect 12287 61423 12373 61479
rect 12429 61423 12515 61479
rect 12571 61423 12657 61479
rect 12713 61423 12799 61479
rect 12855 61423 12941 61479
rect 12997 61423 13083 61479
rect 13139 61423 13225 61479
rect 13281 61423 13367 61479
rect 13423 61423 13509 61479
rect 13565 61423 13651 61479
rect 13707 61423 13793 61479
rect 13849 61423 13935 61479
rect 13991 61423 14077 61479
rect 14133 61423 14219 61479
rect 14275 61423 14361 61479
rect 14417 61423 14503 61479
rect 14559 61423 14645 61479
rect 14701 61423 14787 61479
rect 14843 61423 14853 61479
rect 151 61337 14853 61423
rect 151 61281 161 61337
rect 217 61281 303 61337
rect 359 61281 445 61337
rect 501 61281 587 61337
rect 643 61281 729 61337
rect 785 61281 871 61337
rect 927 61281 1013 61337
rect 1069 61281 1155 61337
rect 1211 61281 1297 61337
rect 1353 61281 1439 61337
rect 1495 61281 1581 61337
rect 1637 61281 1723 61337
rect 1779 61281 1865 61337
rect 1921 61281 2007 61337
rect 2063 61281 2149 61337
rect 2205 61281 2291 61337
rect 2347 61281 2433 61337
rect 2489 61281 2575 61337
rect 2631 61281 2717 61337
rect 2773 61281 2859 61337
rect 2915 61281 3001 61337
rect 3057 61281 3143 61337
rect 3199 61281 3285 61337
rect 3341 61281 3427 61337
rect 3483 61281 3569 61337
rect 3625 61281 3711 61337
rect 3767 61281 3853 61337
rect 3909 61281 3995 61337
rect 4051 61281 4137 61337
rect 4193 61281 4279 61337
rect 4335 61281 4421 61337
rect 4477 61281 4563 61337
rect 4619 61281 4705 61337
rect 4761 61281 4847 61337
rect 4903 61281 4989 61337
rect 5045 61281 5131 61337
rect 5187 61281 5273 61337
rect 5329 61281 5415 61337
rect 5471 61281 5557 61337
rect 5613 61281 5699 61337
rect 5755 61281 5841 61337
rect 5897 61281 5983 61337
rect 6039 61281 6125 61337
rect 6181 61281 6267 61337
rect 6323 61281 6409 61337
rect 6465 61281 6551 61337
rect 6607 61281 6693 61337
rect 6749 61281 6835 61337
rect 6891 61281 6977 61337
rect 7033 61281 7119 61337
rect 7175 61281 7261 61337
rect 7317 61281 7403 61337
rect 7459 61281 7545 61337
rect 7601 61281 7687 61337
rect 7743 61281 7829 61337
rect 7885 61281 7971 61337
rect 8027 61281 8113 61337
rect 8169 61281 8255 61337
rect 8311 61281 8397 61337
rect 8453 61281 8539 61337
rect 8595 61281 8681 61337
rect 8737 61281 8823 61337
rect 8879 61281 8965 61337
rect 9021 61281 9107 61337
rect 9163 61281 9249 61337
rect 9305 61281 9391 61337
rect 9447 61281 9533 61337
rect 9589 61281 9675 61337
rect 9731 61281 9817 61337
rect 9873 61281 9959 61337
rect 10015 61281 10101 61337
rect 10157 61281 10243 61337
rect 10299 61281 10385 61337
rect 10441 61281 10527 61337
rect 10583 61281 10669 61337
rect 10725 61281 10811 61337
rect 10867 61281 10953 61337
rect 11009 61281 11095 61337
rect 11151 61281 11237 61337
rect 11293 61281 11379 61337
rect 11435 61281 11521 61337
rect 11577 61281 11663 61337
rect 11719 61281 11805 61337
rect 11861 61281 11947 61337
rect 12003 61281 12089 61337
rect 12145 61281 12231 61337
rect 12287 61281 12373 61337
rect 12429 61281 12515 61337
rect 12571 61281 12657 61337
rect 12713 61281 12799 61337
rect 12855 61281 12941 61337
rect 12997 61281 13083 61337
rect 13139 61281 13225 61337
rect 13281 61281 13367 61337
rect 13423 61281 13509 61337
rect 13565 61281 13651 61337
rect 13707 61281 13793 61337
rect 13849 61281 13935 61337
rect 13991 61281 14077 61337
rect 14133 61281 14219 61337
rect 14275 61281 14361 61337
rect 14417 61281 14503 61337
rect 14559 61281 14645 61337
rect 14701 61281 14787 61337
rect 14843 61281 14853 61337
rect 151 61195 14853 61281
rect 151 61139 161 61195
rect 217 61139 303 61195
rect 359 61139 445 61195
rect 501 61139 587 61195
rect 643 61139 729 61195
rect 785 61139 871 61195
rect 927 61139 1013 61195
rect 1069 61139 1155 61195
rect 1211 61139 1297 61195
rect 1353 61139 1439 61195
rect 1495 61139 1581 61195
rect 1637 61139 1723 61195
rect 1779 61139 1865 61195
rect 1921 61139 2007 61195
rect 2063 61139 2149 61195
rect 2205 61139 2291 61195
rect 2347 61139 2433 61195
rect 2489 61139 2575 61195
rect 2631 61139 2717 61195
rect 2773 61139 2859 61195
rect 2915 61139 3001 61195
rect 3057 61139 3143 61195
rect 3199 61139 3285 61195
rect 3341 61139 3427 61195
rect 3483 61139 3569 61195
rect 3625 61139 3711 61195
rect 3767 61139 3853 61195
rect 3909 61139 3995 61195
rect 4051 61139 4137 61195
rect 4193 61139 4279 61195
rect 4335 61139 4421 61195
rect 4477 61139 4563 61195
rect 4619 61139 4705 61195
rect 4761 61139 4847 61195
rect 4903 61139 4989 61195
rect 5045 61139 5131 61195
rect 5187 61139 5273 61195
rect 5329 61139 5415 61195
rect 5471 61139 5557 61195
rect 5613 61139 5699 61195
rect 5755 61139 5841 61195
rect 5897 61139 5983 61195
rect 6039 61139 6125 61195
rect 6181 61139 6267 61195
rect 6323 61139 6409 61195
rect 6465 61139 6551 61195
rect 6607 61139 6693 61195
rect 6749 61139 6835 61195
rect 6891 61139 6977 61195
rect 7033 61139 7119 61195
rect 7175 61139 7261 61195
rect 7317 61139 7403 61195
rect 7459 61139 7545 61195
rect 7601 61139 7687 61195
rect 7743 61139 7829 61195
rect 7885 61139 7971 61195
rect 8027 61139 8113 61195
rect 8169 61139 8255 61195
rect 8311 61139 8397 61195
rect 8453 61139 8539 61195
rect 8595 61139 8681 61195
rect 8737 61139 8823 61195
rect 8879 61139 8965 61195
rect 9021 61139 9107 61195
rect 9163 61139 9249 61195
rect 9305 61139 9391 61195
rect 9447 61139 9533 61195
rect 9589 61139 9675 61195
rect 9731 61139 9817 61195
rect 9873 61139 9959 61195
rect 10015 61139 10101 61195
rect 10157 61139 10243 61195
rect 10299 61139 10385 61195
rect 10441 61139 10527 61195
rect 10583 61139 10669 61195
rect 10725 61139 10811 61195
rect 10867 61139 10953 61195
rect 11009 61139 11095 61195
rect 11151 61139 11237 61195
rect 11293 61139 11379 61195
rect 11435 61139 11521 61195
rect 11577 61139 11663 61195
rect 11719 61139 11805 61195
rect 11861 61139 11947 61195
rect 12003 61139 12089 61195
rect 12145 61139 12231 61195
rect 12287 61139 12373 61195
rect 12429 61139 12515 61195
rect 12571 61139 12657 61195
rect 12713 61139 12799 61195
rect 12855 61139 12941 61195
rect 12997 61139 13083 61195
rect 13139 61139 13225 61195
rect 13281 61139 13367 61195
rect 13423 61139 13509 61195
rect 13565 61139 13651 61195
rect 13707 61139 13793 61195
rect 13849 61139 13935 61195
rect 13991 61139 14077 61195
rect 14133 61139 14219 61195
rect 14275 61139 14361 61195
rect 14417 61139 14503 61195
rect 14559 61139 14645 61195
rect 14701 61139 14787 61195
rect 14843 61139 14853 61195
rect 151 61053 14853 61139
rect 151 60997 161 61053
rect 217 60997 303 61053
rect 359 60997 445 61053
rect 501 60997 587 61053
rect 643 60997 729 61053
rect 785 60997 871 61053
rect 927 60997 1013 61053
rect 1069 60997 1155 61053
rect 1211 60997 1297 61053
rect 1353 60997 1439 61053
rect 1495 60997 1581 61053
rect 1637 60997 1723 61053
rect 1779 60997 1865 61053
rect 1921 60997 2007 61053
rect 2063 60997 2149 61053
rect 2205 60997 2291 61053
rect 2347 60997 2433 61053
rect 2489 60997 2575 61053
rect 2631 60997 2717 61053
rect 2773 60997 2859 61053
rect 2915 60997 3001 61053
rect 3057 60997 3143 61053
rect 3199 60997 3285 61053
rect 3341 60997 3427 61053
rect 3483 60997 3569 61053
rect 3625 60997 3711 61053
rect 3767 60997 3853 61053
rect 3909 60997 3995 61053
rect 4051 60997 4137 61053
rect 4193 60997 4279 61053
rect 4335 60997 4421 61053
rect 4477 60997 4563 61053
rect 4619 60997 4705 61053
rect 4761 60997 4847 61053
rect 4903 60997 4989 61053
rect 5045 60997 5131 61053
rect 5187 60997 5273 61053
rect 5329 60997 5415 61053
rect 5471 60997 5557 61053
rect 5613 60997 5699 61053
rect 5755 60997 5841 61053
rect 5897 60997 5983 61053
rect 6039 60997 6125 61053
rect 6181 60997 6267 61053
rect 6323 60997 6409 61053
rect 6465 60997 6551 61053
rect 6607 60997 6693 61053
rect 6749 60997 6835 61053
rect 6891 60997 6977 61053
rect 7033 60997 7119 61053
rect 7175 60997 7261 61053
rect 7317 60997 7403 61053
rect 7459 60997 7545 61053
rect 7601 60997 7687 61053
rect 7743 60997 7829 61053
rect 7885 60997 7971 61053
rect 8027 60997 8113 61053
rect 8169 60997 8255 61053
rect 8311 60997 8397 61053
rect 8453 60997 8539 61053
rect 8595 60997 8681 61053
rect 8737 60997 8823 61053
rect 8879 60997 8965 61053
rect 9021 60997 9107 61053
rect 9163 60997 9249 61053
rect 9305 60997 9391 61053
rect 9447 60997 9533 61053
rect 9589 60997 9675 61053
rect 9731 60997 9817 61053
rect 9873 60997 9959 61053
rect 10015 60997 10101 61053
rect 10157 60997 10243 61053
rect 10299 60997 10385 61053
rect 10441 60997 10527 61053
rect 10583 60997 10669 61053
rect 10725 60997 10811 61053
rect 10867 60997 10953 61053
rect 11009 60997 11095 61053
rect 11151 60997 11237 61053
rect 11293 60997 11379 61053
rect 11435 60997 11521 61053
rect 11577 60997 11663 61053
rect 11719 60997 11805 61053
rect 11861 60997 11947 61053
rect 12003 60997 12089 61053
rect 12145 60997 12231 61053
rect 12287 60997 12373 61053
rect 12429 60997 12515 61053
rect 12571 60997 12657 61053
rect 12713 60997 12799 61053
rect 12855 60997 12941 61053
rect 12997 60997 13083 61053
rect 13139 60997 13225 61053
rect 13281 60997 13367 61053
rect 13423 60997 13509 61053
rect 13565 60997 13651 61053
rect 13707 60997 13793 61053
rect 13849 60997 13935 61053
rect 13991 60997 14077 61053
rect 14133 60997 14219 61053
rect 14275 60997 14361 61053
rect 14417 60997 14503 61053
rect 14559 60997 14645 61053
rect 14701 60997 14787 61053
rect 14843 60997 14853 61053
rect 151 60911 14853 60997
rect 151 60855 161 60911
rect 217 60855 303 60911
rect 359 60855 445 60911
rect 501 60855 587 60911
rect 643 60855 729 60911
rect 785 60855 871 60911
rect 927 60855 1013 60911
rect 1069 60855 1155 60911
rect 1211 60855 1297 60911
rect 1353 60855 1439 60911
rect 1495 60855 1581 60911
rect 1637 60855 1723 60911
rect 1779 60855 1865 60911
rect 1921 60855 2007 60911
rect 2063 60855 2149 60911
rect 2205 60855 2291 60911
rect 2347 60855 2433 60911
rect 2489 60855 2575 60911
rect 2631 60855 2717 60911
rect 2773 60855 2859 60911
rect 2915 60855 3001 60911
rect 3057 60855 3143 60911
rect 3199 60855 3285 60911
rect 3341 60855 3427 60911
rect 3483 60855 3569 60911
rect 3625 60855 3711 60911
rect 3767 60855 3853 60911
rect 3909 60855 3995 60911
rect 4051 60855 4137 60911
rect 4193 60855 4279 60911
rect 4335 60855 4421 60911
rect 4477 60855 4563 60911
rect 4619 60855 4705 60911
rect 4761 60855 4847 60911
rect 4903 60855 4989 60911
rect 5045 60855 5131 60911
rect 5187 60855 5273 60911
rect 5329 60855 5415 60911
rect 5471 60855 5557 60911
rect 5613 60855 5699 60911
rect 5755 60855 5841 60911
rect 5897 60855 5983 60911
rect 6039 60855 6125 60911
rect 6181 60855 6267 60911
rect 6323 60855 6409 60911
rect 6465 60855 6551 60911
rect 6607 60855 6693 60911
rect 6749 60855 6835 60911
rect 6891 60855 6977 60911
rect 7033 60855 7119 60911
rect 7175 60855 7261 60911
rect 7317 60855 7403 60911
rect 7459 60855 7545 60911
rect 7601 60855 7687 60911
rect 7743 60855 7829 60911
rect 7885 60855 7971 60911
rect 8027 60855 8113 60911
rect 8169 60855 8255 60911
rect 8311 60855 8397 60911
rect 8453 60855 8539 60911
rect 8595 60855 8681 60911
rect 8737 60855 8823 60911
rect 8879 60855 8965 60911
rect 9021 60855 9107 60911
rect 9163 60855 9249 60911
rect 9305 60855 9391 60911
rect 9447 60855 9533 60911
rect 9589 60855 9675 60911
rect 9731 60855 9817 60911
rect 9873 60855 9959 60911
rect 10015 60855 10101 60911
rect 10157 60855 10243 60911
rect 10299 60855 10385 60911
rect 10441 60855 10527 60911
rect 10583 60855 10669 60911
rect 10725 60855 10811 60911
rect 10867 60855 10953 60911
rect 11009 60855 11095 60911
rect 11151 60855 11237 60911
rect 11293 60855 11379 60911
rect 11435 60855 11521 60911
rect 11577 60855 11663 60911
rect 11719 60855 11805 60911
rect 11861 60855 11947 60911
rect 12003 60855 12089 60911
rect 12145 60855 12231 60911
rect 12287 60855 12373 60911
rect 12429 60855 12515 60911
rect 12571 60855 12657 60911
rect 12713 60855 12799 60911
rect 12855 60855 12941 60911
rect 12997 60855 13083 60911
rect 13139 60855 13225 60911
rect 13281 60855 13367 60911
rect 13423 60855 13509 60911
rect 13565 60855 13651 60911
rect 13707 60855 13793 60911
rect 13849 60855 13935 60911
rect 13991 60855 14077 60911
rect 14133 60855 14219 60911
rect 14275 60855 14361 60911
rect 14417 60855 14503 60911
rect 14559 60855 14645 60911
rect 14701 60855 14787 60911
rect 14843 60855 14853 60911
rect 151 60769 14853 60855
rect 151 60713 161 60769
rect 217 60713 303 60769
rect 359 60713 445 60769
rect 501 60713 587 60769
rect 643 60713 729 60769
rect 785 60713 871 60769
rect 927 60713 1013 60769
rect 1069 60713 1155 60769
rect 1211 60713 1297 60769
rect 1353 60713 1439 60769
rect 1495 60713 1581 60769
rect 1637 60713 1723 60769
rect 1779 60713 1865 60769
rect 1921 60713 2007 60769
rect 2063 60713 2149 60769
rect 2205 60713 2291 60769
rect 2347 60713 2433 60769
rect 2489 60713 2575 60769
rect 2631 60713 2717 60769
rect 2773 60713 2859 60769
rect 2915 60713 3001 60769
rect 3057 60713 3143 60769
rect 3199 60713 3285 60769
rect 3341 60713 3427 60769
rect 3483 60713 3569 60769
rect 3625 60713 3711 60769
rect 3767 60713 3853 60769
rect 3909 60713 3995 60769
rect 4051 60713 4137 60769
rect 4193 60713 4279 60769
rect 4335 60713 4421 60769
rect 4477 60713 4563 60769
rect 4619 60713 4705 60769
rect 4761 60713 4847 60769
rect 4903 60713 4989 60769
rect 5045 60713 5131 60769
rect 5187 60713 5273 60769
rect 5329 60713 5415 60769
rect 5471 60713 5557 60769
rect 5613 60713 5699 60769
rect 5755 60713 5841 60769
rect 5897 60713 5983 60769
rect 6039 60713 6125 60769
rect 6181 60713 6267 60769
rect 6323 60713 6409 60769
rect 6465 60713 6551 60769
rect 6607 60713 6693 60769
rect 6749 60713 6835 60769
rect 6891 60713 6977 60769
rect 7033 60713 7119 60769
rect 7175 60713 7261 60769
rect 7317 60713 7403 60769
rect 7459 60713 7545 60769
rect 7601 60713 7687 60769
rect 7743 60713 7829 60769
rect 7885 60713 7971 60769
rect 8027 60713 8113 60769
rect 8169 60713 8255 60769
rect 8311 60713 8397 60769
rect 8453 60713 8539 60769
rect 8595 60713 8681 60769
rect 8737 60713 8823 60769
rect 8879 60713 8965 60769
rect 9021 60713 9107 60769
rect 9163 60713 9249 60769
rect 9305 60713 9391 60769
rect 9447 60713 9533 60769
rect 9589 60713 9675 60769
rect 9731 60713 9817 60769
rect 9873 60713 9959 60769
rect 10015 60713 10101 60769
rect 10157 60713 10243 60769
rect 10299 60713 10385 60769
rect 10441 60713 10527 60769
rect 10583 60713 10669 60769
rect 10725 60713 10811 60769
rect 10867 60713 10953 60769
rect 11009 60713 11095 60769
rect 11151 60713 11237 60769
rect 11293 60713 11379 60769
rect 11435 60713 11521 60769
rect 11577 60713 11663 60769
rect 11719 60713 11805 60769
rect 11861 60713 11947 60769
rect 12003 60713 12089 60769
rect 12145 60713 12231 60769
rect 12287 60713 12373 60769
rect 12429 60713 12515 60769
rect 12571 60713 12657 60769
rect 12713 60713 12799 60769
rect 12855 60713 12941 60769
rect 12997 60713 13083 60769
rect 13139 60713 13225 60769
rect 13281 60713 13367 60769
rect 13423 60713 13509 60769
rect 13565 60713 13651 60769
rect 13707 60713 13793 60769
rect 13849 60713 13935 60769
rect 13991 60713 14077 60769
rect 14133 60713 14219 60769
rect 14275 60713 14361 60769
rect 14417 60713 14503 60769
rect 14559 60713 14645 60769
rect 14701 60713 14787 60769
rect 14843 60713 14853 60769
rect 151 60627 14853 60713
rect 151 60571 161 60627
rect 217 60571 303 60627
rect 359 60571 445 60627
rect 501 60571 587 60627
rect 643 60571 729 60627
rect 785 60571 871 60627
rect 927 60571 1013 60627
rect 1069 60571 1155 60627
rect 1211 60571 1297 60627
rect 1353 60571 1439 60627
rect 1495 60571 1581 60627
rect 1637 60571 1723 60627
rect 1779 60571 1865 60627
rect 1921 60571 2007 60627
rect 2063 60571 2149 60627
rect 2205 60571 2291 60627
rect 2347 60571 2433 60627
rect 2489 60571 2575 60627
rect 2631 60571 2717 60627
rect 2773 60571 2859 60627
rect 2915 60571 3001 60627
rect 3057 60571 3143 60627
rect 3199 60571 3285 60627
rect 3341 60571 3427 60627
rect 3483 60571 3569 60627
rect 3625 60571 3711 60627
rect 3767 60571 3853 60627
rect 3909 60571 3995 60627
rect 4051 60571 4137 60627
rect 4193 60571 4279 60627
rect 4335 60571 4421 60627
rect 4477 60571 4563 60627
rect 4619 60571 4705 60627
rect 4761 60571 4847 60627
rect 4903 60571 4989 60627
rect 5045 60571 5131 60627
rect 5187 60571 5273 60627
rect 5329 60571 5415 60627
rect 5471 60571 5557 60627
rect 5613 60571 5699 60627
rect 5755 60571 5841 60627
rect 5897 60571 5983 60627
rect 6039 60571 6125 60627
rect 6181 60571 6267 60627
rect 6323 60571 6409 60627
rect 6465 60571 6551 60627
rect 6607 60571 6693 60627
rect 6749 60571 6835 60627
rect 6891 60571 6977 60627
rect 7033 60571 7119 60627
rect 7175 60571 7261 60627
rect 7317 60571 7403 60627
rect 7459 60571 7545 60627
rect 7601 60571 7687 60627
rect 7743 60571 7829 60627
rect 7885 60571 7971 60627
rect 8027 60571 8113 60627
rect 8169 60571 8255 60627
rect 8311 60571 8397 60627
rect 8453 60571 8539 60627
rect 8595 60571 8681 60627
rect 8737 60571 8823 60627
rect 8879 60571 8965 60627
rect 9021 60571 9107 60627
rect 9163 60571 9249 60627
rect 9305 60571 9391 60627
rect 9447 60571 9533 60627
rect 9589 60571 9675 60627
rect 9731 60571 9817 60627
rect 9873 60571 9959 60627
rect 10015 60571 10101 60627
rect 10157 60571 10243 60627
rect 10299 60571 10385 60627
rect 10441 60571 10527 60627
rect 10583 60571 10669 60627
rect 10725 60571 10811 60627
rect 10867 60571 10953 60627
rect 11009 60571 11095 60627
rect 11151 60571 11237 60627
rect 11293 60571 11379 60627
rect 11435 60571 11521 60627
rect 11577 60571 11663 60627
rect 11719 60571 11805 60627
rect 11861 60571 11947 60627
rect 12003 60571 12089 60627
rect 12145 60571 12231 60627
rect 12287 60571 12373 60627
rect 12429 60571 12515 60627
rect 12571 60571 12657 60627
rect 12713 60571 12799 60627
rect 12855 60571 12941 60627
rect 12997 60571 13083 60627
rect 13139 60571 13225 60627
rect 13281 60571 13367 60627
rect 13423 60571 13509 60627
rect 13565 60571 13651 60627
rect 13707 60571 13793 60627
rect 13849 60571 13935 60627
rect 13991 60571 14077 60627
rect 14133 60571 14219 60627
rect 14275 60571 14361 60627
rect 14417 60571 14503 60627
rect 14559 60571 14645 60627
rect 14701 60571 14787 60627
rect 14843 60571 14853 60627
rect 151 60485 14853 60571
rect 151 60429 161 60485
rect 217 60429 303 60485
rect 359 60429 445 60485
rect 501 60429 587 60485
rect 643 60429 729 60485
rect 785 60429 871 60485
rect 927 60429 1013 60485
rect 1069 60429 1155 60485
rect 1211 60429 1297 60485
rect 1353 60429 1439 60485
rect 1495 60429 1581 60485
rect 1637 60429 1723 60485
rect 1779 60429 1865 60485
rect 1921 60429 2007 60485
rect 2063 60429 2149 60485
rect 2205 60429 2291 60485
rect 2347 60429 2433 60485
rect 2489 60429 2575 60485
rect 2631 60429 2717 60485
rect 2773 60429 2859 60485
rect 2915 60429 3001 60485
rect 3057 60429 3143 60485
rect 3199 60429 3285 60485
rect 3341 60429 3427 60485
rect 3483 60429 3569 60485
rect 3625 60429 3711 60485
rect 3767 60429 3853 60485
rect 3909 60429 3995 60485
rect 4051 60429 4137 60485
rect 4193 60429 4279 60485
rect 4335 60429 4421 60485
rect 4477 60429 4563 60485
rect 4619 60429 4705 60485
rect 4761 60429 4847 60485
rect 4903 60429 4989 60485
rect 5045 60429 5131 60485
rect 5187 60429 5273 60485
rect 5329 60429 5415 60485
rect 5471 60429 5557 60485
rect 5613 60429 5699 60485
rect 5755 60429 5841 60485
rect 5897 60429 5983 60485
rect 6039 60429 6125 60485
rect 6181 60429 6267 60485
rect 6323 60429 6409 60485
rect 6465 60429 6551 60485
rect 6607 60429 6693 60485
rect 6749 60429 6835 60485
rect 6891 60429 6977 60485
rect 7033 60429 7119 60485
rect 7175 60429 7261 60485
rect 7317 60429 7403 60485
rect 7459 60429 7545 60485
rect 7601 60429 7687 60485
rect 7743 60429 7829 60485
rect 7885 60429 7971 60485
rect 8027 60429 8113 60485
rect 8169 60429 8255 60485
rect 8311 60429 8397 60485
rect 8453 60429 8539 60485
rect 8595 60429 8681 60485
rect 8737 60429 8823 60485
rect 8879 60429 8965 60485
rect 9021 60429 9107 60485
rect 9163 60429 9249 60485
rect 9305 60429 9391 60485
rect 9447 60429 9533 60485
rect 9589 60429 9675 60485
rect 9731 60429 9817 60485
rect 9873 60429 9959 60485
rect 10015 60429 10101 60485
rect 10157 60429 10243 60485
rect 10299 60429 10385 60485
rect 10441 60429 10527 60485
rect 10583 60429 10669 60485
rect 10725 60429 10811 60485
rect 10867 60429 10953 60485
rect 11009 60429 11095 60485
rect 11151 60429 11237 60485
rect 11293 60429 11379 60485
rect 11435 60429 11521 60485
rect 11577 60429 11663 60485
rect 11719 60429 11805 60485
rect 11861 60429 11947 60485
rect 12003 60429 12089 60485
rect 12145 60429 12231 60485
rect 12287 60429 12373 60485
rect 12429 60429 12515 60485
rect 12571 60429 12657 60485
rect 12713 60429 12799 60485
rect 12855 60429 12941 60485
rect 12997 60429 13083 60485
rect 13139 60429 13225 60485
rect 13281 60429 13367 60485
rect 13423 60429 13509 60485
rect 13565 60429 13651 60485
rect 13707 60429 13793 60485
rect 13849 60429 13935 60485
rect 13991 60429 14077 60485
rect 14133 60429 14219 60485
rect 14275 60429 14361 60485
rect 14417 60429 14503 60485
rect 14559 60429 14645 60485
rect 14701 60429 14787 60485
rect 14843 60429 14853 60485
rect 151 60419 14853 60429
rect 151 60171 14853 60181
rect 151 60115 161 60171
rect 217 60115 303 60171
rect 359 60115 445 60171
rect 501 60115 587 60171
rect 643 60115 729 60171
rect 785 60115 871 60171
rect 927 60115 1013 60171
rect 1069 60115 1155 60171
rect 1211 60115 1297 60171
rect 1353 60115 1439 60171
rect 1495 60115 1581 60171
rect 1637 60115 1723 60171
rect 1779 60115 1865 60171
rect 1921 60115 2007 60171
rect 2063 60115 2149 60171
rect 2205 60115 2291 60171
rect 2347 60115 2433 60171
rect 2489 60115 2575 60171
rect 2631 60115 2717 60171
rect 2773 60115 2859 60171
rect 2915 60115 3001 60171
rect 3057 60115 3143 60171
rect 3199 60115 3285 60171
rect 3341 60115 3427 60171
rect 3483 60115 3569 60171
rect 3625 60115 3711 60171
rect 3767 60115 3853 60171
rect 3909 60115 3995 60171
rect 4051 60115 4137 60171
rect 4193 60115 4279 60171
rect 4335 60115 4421 60171
rect 4477 60115 4563 60171
rect 4619 60115 4705 60171
rect 4761 60115 4847 60171
rect 4903 60115 4989 60171
rect 5045 60115 5131 60171
rect 5187 60115 5273 60171
rect 5329 60115 5415 60171
rect 5471 60115 5557 60171
rect 5613 60115 5699 60171
rect 5755 60115 5841 60171
rect 5897 60115 5983 60171
rect 6039 60115 6125 60171
rect 6181 60115 6267 60171
rect 6323 60115 6409 60171
rect 6465 60115 6551 60171
rect 6607 60115 6693 60171
rect 6749 60115 6835 60171
rect 6891 60115 6977 60171
rect 7033 60115 7119 60171
rect 7175 60115 7261 60171
rect 7317 60115 7403 60171
rect 7459 60115 7545 60171
rect 7601 60115 7687 60171
rect 7743 60115 7829 60171
rect 7885 60115 7971 60171
rect 8027 60115 8113 60171
rect 8169 60115 8255 60171
rect 8311 60115 8397 60171
rect 8453 60115 8539 60171
rect 8595 60115 8681 60171
rect 8737 60115 8823 60171
rect 8879 60115 8965 60171
rect 9021 60115 9107 60171
rect 9163 60115 9249 60171
rect 9305 60115 9391 60171
rect 9447 60115 9533 60171
rect 9589 60115 9675 60171
rect 9731 60115 9817 60171
rect 9873 60115 9959 60171
rect 10015 60115 10101 60171
rect 10157 60115 10243 60171
rect 10299 60115 10385 60171
rect 10441 60115 10527 60171
rect 10583 60115 10669 60171
rect 10725 60115 10811 60171
rect 10867 60115 10953 60171
rect 11009 60115 11095 60171
rect 11151 60115 11237 60171
rect 11293 60115 11379 60171
rect 11435 60115 11521 60171
rect 11577 60115 11663 60171
rect 11719 60115 11805 60171
rect 11861 60115 11947 60171
rect 12003 60115 12089 60171
rect 12145 60115 12231 60171
rect 12287 60115 12373 60171
rect 12429 60115 12515 60171
rect 12571 60115 12657 60171
rect 12713 60115 12799 60171
rect 12855 60115 12941 60171
rect 12997 60115 13083 60171
rect 13139 60115 13225 60171
rect 13281 60115 13367 60171
rect 13423 60115 13509 60171
rect 13565 60115 13651 60171
rect 13707 60115 13793 60171
rect 13849 60115 13935 60171
rect 13991 60115 14077 60171
rect 14133 60115 14219 60171
rect 14275 60115 14361 60171
rect 14417 60115 14503 60171
rect 14559 60115 14645 60171
rect 14701 60115 14787 60171
rect 14843 60115 14853 60171
rect 151 60029 14853 60115
rect 151 59973 161 60029
rect 217 59973 303 60029
rect 359 59973 445 60029
rect 501 59973 587 60029
rect 643 59973 729 60029
rect 785 59973 871 60029
rect 927 59973 1013 60029
rect 1069 59973 1155 60029
rect 1211 59973 1297 60029
rect 1353 59973 1439 60029
rect 1495 59973 1581 60029
rect 1637 59973 1723 60029
rect 1779 59973 1865 60029
rect 1921 59973 2007 60029
rect 2063 59973 2149 60029
rect 2205 59973 2291 60029
rect 2347 59973 2433 60029
rect 2489 59973 2575 60029
rect 2631 59973 2717 60029
rect 2773 59973 2859 60029
rect 2915 59973 3001 60029
rect 3057 59973 3143 60029
rect 3199 59973 3285 60029
rect 3341 59973 3427 60029
rect 3483 59973 3569 60029
rect 3625 59973 3711 60029
rect 3767 59973 3853 60029
rect 3909 59973 3995 60029
rect 4051 59973 4137 60029
rect 4193 59973 4279 60029
rect 4335 59973 4421 60029
rect 4477 59973 4563 60029
rect 4619 59973 4705 60029
rect 4761 59973 4847 60029
rect 4903 59973 4989 60029
rect 5045 59973 5131 60029
rect 5187 59973 5273 60029
rect 5329 59973 5415 60029
rect 5471 59973 5557 60029
rect 5613 59973 5699 60029
rect 5755 59973 5841 60029
rect 5897 59973 5983 60029
rect 6039 59973 6125 60029
rect 6181 59973 6267 60029
rect 6323 59973 6409 60029
rect 6465 59973 6551 60029
rect 6607 59973 6693 60029
rect 6749 59973 6835 60029
rect 6891 59973 6977 60029
rect 7033 59973 7119 60029
rect 7175 59973 7261 60029
rect 7317 59973 7403 60029
rect 7459 59973 7545 60029
rect 7601 59973 7687 60029
rect 7743 59973 7829 60029
rect 7885 59973 7971 60029
rect 8027 59973 8113 60029
rect 8169 59973 8255 60029
rect 8311 59973 8397 60029
rect 8453 59973 8539 60029
rect 8595 59973 8681 60029
rect 8737 59973 8823 60029
rect 8879 59973 8965 60029
rect 9021 59973 9107 60029
rect 9163 59973 9249 60029
rect 9305 59973 9391 60029
rect 9447 59973 9533 60029
rect 9589 59973 9675 60029
rect 9731 59973 9817 60029
rect 9873 59973 9959 60029
rect 10015 59973 10101 60029
rect 10157 59973 10243 60029
rect 10299 59973 10385 60029
rect 10441 59973 10527 60029
rect 10583 59973 10669 60029
rect 10725 59973 10811 60029
rect 10867 59973 10953 60029
rect 11009 59973 11095 60029
rect 11151 59973 11237 60029
rect 11293 59973 11379 60029
rect 11435 59973 11521 60029
rect 11577 59973 11663 60029
rect 11719 59973 11805 60029
rect 11861 59973 11947 60029
rect 12003 59973 12089 60029
rect 12145 59973 12231 60029
rect 12287 59973 12373 60029
rect 12429 59973 12515 60029
rect 12571 59973 12657 60029
rect 12713 59973 12799 60029
rect 12855 59973 12941 60029
rect 12997 59973 13083 60029
rect 13139 59973 13225 60029
rect 13281 59973 13367 60029
rect 13423 59973 13509 60029
rect 13565 59973 13651 60029
rect 13707 59973 13793 60029
rect 13849 59973 13935 60029
rect 13991 59973 14077 60029
rect 14133 59973 14219 60029
rect 14275 59973 14361 60029
rect 14417 59973 14503 60029
rect 14559 59973 14645 60029
rect 14701 59973 14787 60029
rect 14843 59973 14853 60029
rect 151 59887 14853 59973
rect 151 59831 161 59887
rect 217 59831 303 59887
rect 359 59831 445 59887
rect 501 59831 587 59887
rect 643 59831 729 59887
rect 785 59831 871 59887
rect 927 59831 1013 59887
rect 1069 59831 1155 59887
rect 1211 59831 1297 59887
rect 1353 59831 1439 59887
rect 1495 59831 1581 59887
rect 1637 59831 1723 59887
rect 1779 59831 1865 59887
rect 1921 59831 2007 59887
rect 2063 59831 2149 59887
rect 2205 59831 2291 59887
rect 2347 59831 2433 59887
rect 2489 59831 2575 59887
rect 2631 59831 2717 59887
rect 2773 59831 2859 59887
rect 2915 59831 3001 59887
rect 3057 59831 3143 59887
rect 3199 59831 3285 59887
rect 3341 59831 3427 59887
rect 3483 59831 3569 59887
rect 3625 59831 3711 59887
rect 3767 59831 3853 59887
rect 3909 59831 3995 59887
rect 4051 59831 4137 59887
rect 4193 59831 4279 59887
rect 4335 59831 4421 59887
rect 4477 59831 4563 59887
rect 4619 59831 4705 59887
rect 4761 59831 4847 59887
rect 4903 59831 4989 59887
rect 5045 59831 5131 59887
rect 5187 59831 5273 59887
rect 5329 59831 5415 59887
rect 5471 59831 5557 59887
rect 5613 59831 5699 59887
rect 5755 59831 5841 59887
rect 5897 59831 5983 59887
rect 6039 59831 6125 59887
rect 6181 59831 6267 59887
rect 6323 59831 6409 59887
rect 6465 59831 6551 59887
rect 6607 59831 6693 59887
rect 6749 59831 6835 59887
rect 6891 59831 6977 59887
rect 7033 59831 7119 59887
rect 7175 59831 7261 59887
rect 7317 59831 7403 59887
rect 7459 59831 7545 59887
rect 7601 59831 7687 59887
rect 7743 59831 7829 59887
rect 7885 59831 7971 59887
rect 8027 59831 8113 59887
rect 8169 59831 8255 59887
rect 8311 59831 8397 59887
rect 8453 59831 8539 59887
rect 8595 59831 8681 59887
rect 8737 59831 8823 59887
rect 8879 59831 8965 59887
rect 9021 59831 9107 59887
rect 9163 59831 9249 59887
rect 9305 59831 9391 59887
rect 9447 59831 9533 59887
rect 9589 59831 9675 59887
rect 9731 59831 9817 59887
rect 9873 59831 9959 59887
rect 10015 59831 10101 59887
rect 10157 59831 10243 59887
rect 10299 59831 10385 59887
rect 10441 59831 10527 59887
rect 10583 59831 10669 59887
rect 10725 59831 10811 59887
rect 10867 59831 10953 59887
rect 11009 59831 11095 59887
rect 11151 59831 11237 59887
rect 11293 59831 11379 59887
rect 11435 59831 11521 59887
rect 11577 59831 11663 59887
rect 11719 59831 11805 59887
rect 11861 59831 11947 59887
rect 12003 59831 12089 59887
rect 12145 59831 12231 59887
rect 12287 59831 12373 59887
rect 12429 59831 12515 59887
rect 12571 59831 12657 59887
rect 12713 59831 12799 59887
rect 12855 59831 12941 59887
rect 12997 59831 13083 59887
rect 13139 59831 13225 59887
rect 13281 59831 13367 59887
rect 13423 59831 13509 59887
rect 13565 59831 13651 59887
rect 13707 59831 13793 59887
rect 13849 59831 13935 59887
rect 13991 59831 14077 59887
rect 14133 59831 14219 59887
rect 14275 59831 14361 59887
rect 14417 59831 14503 59887
rect 14559 59831 14645 59887
rect 14701 59831 14787 59887
rect 14843 59831 14853 59887
rect 151 59745 14853 59831
rect 151 59689 161 59745
rect 217 59689 303 59745
rect 359 59689 445 59745
rect 501 59689 587 59745
rect 643 59689 729 59745
rect 785 59689 871 59745
rect 927 59689 1013 59745
rect 1069 59689 1155 59745
rect 1211 59689 1297 59745
rect 1353 59689 1439 59745
rect 1495 59689 1581 59745
rect 1637 59689 1723 59745
rect 1779 59689 1865 59745
rect 1921 59689 2007 59745
rect 2063 59689 2149 59745
rect 2205 59689 2291 59745
rect 2347 59689 2433 59745
rect 2489 59689 2575 59745
rect 2631 59689 2717 59745
rect 2773 59689 2859 59745
rect 2915 59689 3001 59745
rect 3057 59689 3143 59745
rect 3199 59689 3285 59745
rect 3341 59689 3427 59745
rect 3483 59689 3569 59745
rect 3625 59689 3711 59745
rect 3767 59689 3853 59745
rect 3909 59689 3995 59745
rect 4051 59689 4137 59745
rect 4193 59689 4279 59745
rect 4335 59689 4421 59745
rect 4477 59689 4563 59745
rect 4619 59689 4705 59745
rect 4761 59689 4847 59745
rect 4903 59689 4989 59745
rect 5045 59689 5131 59745
rect 5187 59689 5273 59745
rect 5329 59689 5415 59745
rect 5471 59689 5557 59745
rect 5613 59689 5699 59745
rect 5755 59689 5841 59745
rect 5897 59689 5983 59745
rect 6039 59689 6125 59745
rect 6181 59689 6267 59745
rect 6323 59689 6409 59745
rect 6465 59689 6551 59745
rect 6607 59689 6693 59745
rect 6749 59689 6835 59745
rect 6891 59689 6977 59745
rect 7033 59689 7119 59745
rect 7175 59689 7261 59745
rect 7317 59689 7403 59745
rect 7459 59689 7545 59745
rect 7601 59689 7687 59745
rect 7743 59689 7829 59745
rect 7885 59689 7971 59745
rect 8027 59689 8113 59745
rect 8169 59689 8255 59745
rect 8311 59689 8397 59745
rect 8453 59689 8539 59745
rect 8595 59689 8681 59745
rect 8737 59689 8823 59745
rect 8879 59689 8965 59745
rect 9021 59689 9107 59745
rect 9163 59689 9249 59745
rect 9305 59689 9391 59745
rect 9447 59689 9533 59745
rect 9589 59689 9675 59745
rect 9731 59689 9817 59745
rect 9873 59689 9959 59745
rect 10015 59689 10101 59745
rect 10157 59689 10243 59745
rect 10299 59689 10385 59745
rect 10441 59689 10527 59745
rect 10583 59689 10669 59745
rect 10725 59689 10811 59745
rect 10867 59689 10953 59745
rect 11009 59689 11095 59745
rect 11151 59689 11237 59745
rect 11293 59689 11379 59745
rect 11435 59689 11521 59745
rect 11577 59689 11663 59745
rect 11719 59689 11805 59745
rect 11861 59689 11947 59745
rect 12003 59689 12089 59745
rect 12145 59689 12231 59745
rect 12287 59689 12373 59745
rect 12429 59689 12515 59745
rect 12571 59689 12657 59745
rect 12713 59689 12799 59745
rect 12855 59689 12941 59745
rect 12997 59689 13083 59745
rect 13139 59689 13225 59745
rect 13281 59689 13367 59745
rect 13423 59689 13509 59745
rect 13565 59689 13651 59745
rect 13707 59689 13793 59745
rect 13849 59689 13935 59745
rect 13991 59689 14077 59745
rect 14133 59689 14219 59745
rect 14275 59689 14361 59745
rect 14417 59689 14503 59745
rect 14559 59689 14645 59745
rect 14701 59689 14787 59745
rect 14843 59689 14853 59745
rect 151 59603 14853 59689
rect 151 59547 161 59603
rect 217 59547 303 59603
rect 359 59547 445 59603
rect 501 59547 587 59603
rect 643 59547 729 59603
rect 785 59547 871 59603
rect 927 59547 1013 59603
rect 1069 59547 1155 59603
rect 1211 59547 1297 59603
rect 1353 59547 1439 59603
rect 1495 59547 1581 59603
rect 1637 59547 1723 59603
rect 1779 59547 1865 59603
rect 1921 59547 2007 59603
rect 2063 59547 2149 59603
rect 2205 59547 2291 59603
rect 2347 59547 2433 59603
rect 2489 59547 2575 59603
rect 2631 59547 2717 59603
rect 2773 59547 2859 59603
rect 2915 59547 3001 59603
rect 3057 59547 3143 59603
rect 3199 59547 3285 59603
rect 3341 59547 3427 59603
rect 3483 59547 3569 59603
rect 3625 59547 3711 59603
rect 3767 59547 3853 59603
rect 3909 59547 3995 59603
rect 4051 59547 4137 59603
rect 4193 59547 4279 59603
rect 4335 59547 4421 59603
rect 4477 59547 4563 59603
rect 4619 59547 4705 59603
rect 4761 59547 4847 59603
rect 4903 59547 4989 59603
rect 5045 59547 5131 59603
rect 5187 59547 5273 59603
rect 5329 59547 5415 59603
rect 5471 59547 5557 59603
rect 5613 59547 5699 59603
rect 5755 59547 5841 59603
rect 5897 59547 5983 59603
rect 6039 59547 6125 59603
rect 6181 59547 6267 59603
rect 6323 59547 6409 59603
rect 6465 59547 6551 59603
rect 6607 59547 6693 59603
rect 6749 59547 6835 59603
rect 6891 59547 6977 59603
rect 7033 59547 7119 59603
rect 7175 59547 7261 59603
rect 7317 59547 7403 59603
rect 7459 59547 7545 59603
rect 7601 59547 7687 59603
rect 7743 59547 7829 59603
rect 7885 59547 7971 59603
rect 8027 59547 8113 59603
rect 8169 59547 8255 59603
rect 8311 59547 8397 59603
rect 8453 59547 8539 59603
rect 8595 59547 8681 59603
rect 8737 59547 8823 59603
rect 8879 59547 8965 59603
rect 9021 59547 9107 59603
rect 9163 59547 9249 59603
rect 9305 59547 9391 59603
rect 9447 59547 9533 59603
rect 9589 59547 9675 59603
rect 9731 59547 9817 59603
rect 9873 59547 9959 59603
rect 10015 59547 10101 59603
rect 10157 59547 10243 59603
rect 10299 59547 10385 59603
rect 10441 59547 10527 59603
rect 10583 59547 10669 59603
rect 10725 59547 10811 59603
rect 10867 59547 10953 59603
rect 11009 59547 11095 59603
rect 11151 59547 11237 59603
rect 11293 59547 11379 59603
rect 11435 59547 11521 59603
rect 11577 59547 11663 59603
rect 11719 59547 11805 59603
rect 11861 59547 11947 59603
rect 12003 59547 12089 59603
rect 12145 59547 12231 59603
rect 12287 59547 12373 59603
rect 12429 59547 12515 59603
rect 12571 59547 12657 59603
rect 12713 59547 12799 59603
rect 12855 59547 12941 59603
rect 12997 59547 13083 59603
rect 13139 59547 13225 59603
rect 13281 59547 13367 59603
rect 13423 59547 13509 59603
rect 13565 59547 13651 59603
rect 13707 59547 13793 59603
rect 13849 59547 13935 59603
rect 13991 59547 14077 59603
rect 14133 59547 14219 59603
rect 14275 59547 14361 59603
rect 14417 59547 14503 59603
rect 14559 59547 14645 59603
rect 14701 59547 14787 59603
rect 14843 59547 14853 59603
rect 151 59461 14853 59547
rect 151 59405 161 59461
rect 217 59405 303 59461
rect 359 59405 445 59461
rect 501 59405 587 59461
rect 643 59405 729 59461
rect 785 59405 871 59461
rect 927 59405 1013 59461
rect 1069 59405 1155 59461
rect 1211 59405 1297 59461
rect 1353 59405 1439 59461
rect 1495 59405 1581 59461
rect 1637 59405 1723 59461
rect 1779 59405 1865 59461
rect 1921 59405 2007 59461
rect 2063 59405 2149 59461
rect 2205 59405 2291 59461
rect 2347 59405 2433 59461
rect 2489 59405 2575 59461
rect 2631 59405 2717 59461
rect 2773 59405 2859 59461
rect 2915 59405 3001 59461
rect 3057 59405 3143 59461
rect 3199 59405 3285 59461
rect 3341 59405 3427 59461
rect 3483 59405 3569 59461
rect 3625 59405 3711 59461
rect 3767 59405 3853 59461
rect 3909 59405 3995 59461
rect 4051 59405 4137 59461
rect 4193 59405 4279 59461
rect 4335 59405 4421 59461
rect 4477 59405 4563 59461
rect 4619 59405 4705 59461
rect 4761 59405 4847 59461
rect 4903 59405 4989 59461
rect 5045 59405 5131 59461
rect 5187 59405 5273 59461
rect 5329 59405 5415 59461
rect 5471 59405 5557 59461
rect 5613 59405 5699 59461
rect 5755 59405 5841 59461
rect 5897 59405 5983 59461
rect 6039 59405 6125 59461
rect 6181 59405 6267 59461
rect 6323 59405 6409 59461
rect 6465 59405 6551 59461
rect 6607 59405 6693 59461
rect 6749 59405 6835 59461
rect 6891 59405 6977 59461
rect 7033 59405 7119 59461
rect 7175 59405 7261 59461
rect 7317 59405 7403 59461
rect 7459 59405 7545 59461
rect 7601 59405 7687 59461
rect 7743 59405 7829 59461
rect 7885 59405 7971 59461
rect 8027 59405 8113 59461
rect 8169 59405 8255 59461
rect 8311 59405 8397 59461
rect 8453 59405 8539 59461
rect 8595 59405 8681 59461
rect 8737 59405 8823 59461
rect 8879 59405 8965 59461
rect 9021 59405 9107 59461
rect 9163 59405 9249 59461
rect 9305 59405 9391 59461
rect 9447 59405 9533 59461
rect 9589 59405 9675 59461
rect 9731 59405 9817 59461
rect 9873 59405 9959 59461
rect 10015 59405 10101 59461
rect 10157 59405 10243 59461
rect 10299 59405 10385 59461
rect 10441 59405 10527 59461
rect 10583 59405 10669 59461
rect 10725 59405 10811 59461
rect 10867 59405 10953 59461
rect 11009 59405 11095 59461
rect 11151 59405 11237 59461
rect 11293 59405 11379 59461
rect 11435 59405 11521 59461
rect 11577 59405 11663 59461
rect 11719 59405 11805 59461
rect 11861 59405 11947 59461
rect 12003 59405 12089 59461
rect 12145 59405 12231 59461
rect 12287 59405 12373 59461
rect 12429 59405 12515 59461
rect 12571 59405 12657 59461
rect 12713 59405 12799 59461
rect 12855 59405 12941 59461
rect 12997 59405 13083 59461
rect 13139 59405 13225 59461
rect 13281 59405 13367 59461
rect 13423 59405 13509 59461
rect 13565 59405 13651 59461
rect 13707 59405 13793 59461
rect 13849 59405 13935 59461
rect 13991 59405 14077 59461
rect 14133 59405 14219 59461
rect 14275 59405 14361 59461
rect 14417 59405 14503 59461
rect 14559 59405 14645 59461
rect 14701 59405 14787 59461
rect 14843 59405 14853 59461
rect 151 59319 14853 59405
rect 151 59263 161 59319
rect 217 59263 303 59319
rect 359 59263 445 59319
rect 501 59263 587 59319
rect 643 59263 729 59319
rect 785 59263 871 59319
rect 927 59263 1013 59319
rect 1069 59263 1155 59319
rect 1211 59263 1297 59319
rect 1353 59263 1439 59319
rect 1495 59263 1581 59319
rect 1637 59263 1723 59319
rect 1779 59263 1865 59319
rect 1921 59263 2007 59319
rect 2063 59263 2149 59319
rect 2205 59263 2291 59319
rect 2347 59263 2433 59319
rect 2489 59263 2575 59319
rect 2631 59263 2717 59319
rect 2773 59263 2859 59319
rect 2915 59263 3001 59319
rect 3057 59263 3143 59319
rect 3199 59263 3285 59319
rect 3341 59263 3427 59319
rect 3483 59263 3569 59319
rect 3625 59263 3711 59319
rect 3767 59263 3853 59319
rect 3909 59263 3995 59319
rect 4051 59263 4137 59319
rect 4193 59263 4279 59319
rect 4335 59263 4421 59319
rect 4477 59263 4563 59319
rect 4619 59263 4705 59319
rect 4761 59263 4847 59319
rect 4903 59263 4989 59319
rect 5045 59263 5131 59319
rect 5187 59263 5273 59319
rect 5329 59263 5415 59319
rect 5471 59263 5557 59319
rect 5613 59263 5699 59319
rect 5755 59263 5841 59319
rect 5897 59263 5983 59319
rect 6039 59263 6125 59319
rect 6181 59263 6267 59319
rect 6323 59263 6409 59319
rect 6465 59263 6551 59319
rect 6607 59263 6693 59319
rect 6749 59263 6835 59319
rect 6891 59263 6977 59319
rect 7033 59263 7119 59319
rect 7175 59263 7261 59319
rect 7317 59263 7403 59319
rect 7459 59263 7545 59319
rect 7601 59263 7687 59319
rect 7743 59263 7829 59319
rect 7885 59263 7971 59319
rect 8027 59263 8113 59319
rect 8169 59263 8255 59319
rect 8311 59263 8397 59319
rect 8453 59263 8539 59319
rect 8595 59263 8681 59319
rect 8737 59263 8823 59319
rect 8879 59263 8965 59319
rect 9021 59263 9107 59319
rect 9163 59263 9249 59319
rect 9305 59263 9391 59319
rect 9447 59263 9533 59319
rect 9589 59263 9675 59319
rect 9731 59263 9817 59319
rect 9873 59263 9959 59319
rect 10015 59263 10101 59319
rect 10157 59263 10243 59319
rect 10299 59263 10385 59319
rect 10441 59263 10527 59319
rect 10583 59263 10669 59319
rect 10725 59263 10811 59319
rect 10867 59263 10953 59319
rect 11009 59263 11095 59319
rect 11151 59263 11237 59319
rect 11293 59263 11379 59319
rect 11435 59263 11521 59319
rect 11577 59263 11663 59319
rect 11719 59263 11805 59319
rect 11861 59263 11947 59319
rect 12003 59263 12089 59319
rect 12145 59263 12231 59319
rect 12287 59263 12373 59319
rect 12429 59263 12515 59319
rect 12571 59263 12657 59319
rect 12713 59263 12799 59319
rect 12855 59263 12941 59319
rect 12997 59263 13083 59319
rect 13139 59263 13225 59319
rect 13281 59263 13367 59319
rect 13423 59263 13509 59319
rect 13565 59263 13651 59319
rect 13707 59263 13793 59319
rect 13849 59263 13935 59319
rect 13991 59263 14077 59319
rect 14133 59263 14219 59319
rect 14275 59263 14361 59319
rect 14417 59263 14503 59319
rect 14559 59263 14645 59319
rect 14701 59263 14787 59319
rect 14843 59263 14853 59319
rect 151 59177 14853 59263
rect 151 59121 161 59177
rect 217 59121 303 59177
rect 359 59121 445 59177
rect 501 59121 587 59177
rect 643 59121 729 59177
rect 785 59121 871 59177
rect 927 59121 1013 59177
rect 1069 59121 1155 59177
rect 1211 59121 1297 59177
rect 1353 59121 1439 59177
rect 1495 59121 1581 59177
rect 1637 59121 1723 59177
rect 1779 59121 1865 59177
rect 1921 59121 2007 59177
rect 2063 59121 2149 59177
rect 2205 59121 2291 59177
rect 2347 59121 2433 59177
rect 2489 59121 2575 59177
rect 2631 59121 2717 59177
rect 2773 59121 2859 59177
rect 2915 59121 3001 59177
rect 3057 59121 3143 59177
rect 3199 59121 3285 59177
rect 3341 59121 3427 59177
rect 3483 59121 3569 59177
rect 3625 59121 3711 59177
rect 3767 59121 3853 59177
rect 3909 59121 3995 59177
rect 4051 59121 4137 59177
rect 4193 59121 4279 59177
rect 4335 59121 4421 59177
rect 4477 59121 4563 59177
rect 4619 59121 4705 59177
rect 4761 59121 4847 59177
rect 4903 59121 4989 59177
rect 5045 59121 5131 59177
rect 5187 59121 5273 59177
rect 5329 59121 5415 59177
rect 5471 59121 5557 59177
rect 5613 59121 5699 59177
rect 5755 59121 5841 59177
rect 5897 59121 5983 59177
rect 6039 59121 6125 59177
rect 6181 59121 6267 59177
rect 6323 59121 6409 59177
rect 6465 59121 6551 59177
rect 6607 59121 6693 59177
rect 6749 59121 6835 59177
rect 6891 59121 6977 59177
rect 7033 59121 7119 59177
rect 7175 59121 7261 59177
rect 7317 59121 7403 59177
rect 7459 59121 7545 59177
rect 7601 59121 7687 59177
rect 7743 59121 7829 59177
rect 7885 59121 7971 59177
rect 8027 59121 8113 59177
rect 8169 59121 8255 59177
rect 8311 59121 8397 59177
rect 8453 59121 8539 59177
rect 8595 59121 8681 59177
rect 8737 59121 8823 59177
rect 8879 59121 8965 59177
rect 9021 59121 9107 59177
rect 9163 59121 9249 59177
rect 9305 59121 9391 59177
rect 9447 59121 9533 59177
rect 9589 59121 9675 59177
rect 9731 59121 9817 59177
rect 9873 59121 9959 59177
rect 10015 59121 10101 59177
rect 10157 59121 10243 59177
rect 10299 59121 10385 59177
rect 10441 59121 10527 59177
rect 10583 59121 10669 59177
rect 10725 59121 10811 59177
rect 10867 59121 10953 59177
rect 11009 59121 11095 59177
rect 11151 59121 11237 59177
rect 11293 59121 11379 59177
rect 11435 59121 11521 59177
rect 11577 59121 11663 59177
rect 11719 59121 11805 59177
rect 11861 59121 11947 59177
rect 12003 59121 12089 59177
rect 12145 59121 12231 59177
rect 12287 59121 12373 59177
rect 12429 59121 12515 59177
rect 12571 59121 12657 59177
rect 12713 59121 12799 59177
rect 12855 59121 12941 59177
rect 12997 59121 13083 59177
rect 13139 59121 13225 59177
rect 13281 59121 13367 59177
rect 13423 59121 13509 59177
rect 13565 59121 13651 59177
rect 13707 59121 13793 59177
rect 13849 59121 13935 59177
rect 13991 59121 14077 59177
rect 14133 59121 14219 59177
rect 14275 59121 14361 59177
rect 14417 59121 14503 59177
rect 14559 59121 14645 59177
rect 14701 59121 14787 59177
rect 14843 59121 14853 59177
rect 151 59035 14853 59121
rect 151 58979 161 59035
rect 217 58979 303 59035
rect 359 58979 445 59035
rect 501 58979 587 59035
rect 643 58979 729 59035
rect 785 58979 871 59035
rect 927 58979 1013 59035
rect 1069 58979 1155 59035
rect 1211 58979 1297 59035
rect 1353 58979 1439 59035
rect 1495 58979 1581 59035
rect 1637 58979 1723 59035
rect 1779 58979 1865 59035
rect 1921 58979 2007 59035
rect 2063 58979 2149 59035
rect 2205 58979 2291 59035
rect 2347 58979 2433 59035
rect 2489 58979 2575 59035
rect 2631 58979 2717 59035
rect 2773 58979 2859 59035
rect 2915 58979 3001 59035
rect 3057 58979 3143 59035
rect 3199 58979 3285 59035
rect 3341 58979 3427 59035
rect 3483 58979 3569 59035
rect 3625 58979 3711 59035
rect 3767 58979 3853 59035
rect 3909 58979 3995 59035
rect 4051 58979 4137 59035
rect 4193 58979 4279 59035
rect 4335 58979 4421 59035
rect 4477 58979 4563 59035
rect 4619 58979 4705 59035
rect 4761 58979 4847 59035
rect 4903 58979 4989 59035
rect 5045 58979 5131 59035
rect 5187 58979 5273 59035
rect 5329 58979 5415 59035
rect 5471 58979 5557 59035
rect 5613 58979 5699 59035
rect 5755 58979 5841 59035
rect 5897 58979 5983 59035
rect 6039 58979 6125 59035
rect 6181 58979 6267 59035
rect 6323 58979 6409 59035
rect 6465 58979 6551 59035
rect 6607 58979 6693 59035
rect 6749 58979 6835 59035
rect 6891 58979 6977 59035
rect 7033 58979 7119 59035
rect 7175 58979 7261 59035
rect 7317 58979 7403 59035
rect 7459 58979 7545 59035
rect 7601 58979 7687 59035
rect 7743 58979 7829 59035
rect 7885 58979 7971 59035
rect 8027 58979 8113 59035
rect 8169 58979 8255 59035
rect 8311 58979 8397 59035
rect 8453 58979 8539 59035
rect 8595 58979 8681 59035
rect 8737 58979 8823 59035
rect 8879 58979 8965 59035
rect 9021 58979 9107 59035
rect 9163 58979 9249 59035
rect 9305 58979 9391 59035
rect 9447 58979 9533 59035
rect 9589 58979 9675 59035
rect 9731 58979 9817 59035
rect 9873 58979 9959 59035
rect 10015 58979 10101 59035
rect 10157 58979 10243 59035
rect 10299 58979 10385 59035
rect 10441 58979 10527 59035
rect 10583 58979 10669 59035
rect 10725 58979 10811 59035
rect 10867 58979 10953 59035
rect 11009 58979 11095 59035
rect 11151 58979 11237 59035
rect 11293 58979 11379 59035
rect 11435 58979 11521 59035
rect 11577 58979 11663 59035
rect 11719 58979 11805 59035
rect 11861 58979 11947 59035
rect 12003 58979 12089 59035
rect 12145 58979 12231 59035
rect 12287 58979 12373 59035
rect 12429 58979 12515 59035
rect 12571 58979 12657 59035
rect 12713 58979 12799 59035
rect 12855 58979 12941 59035
rect 12997 58979 13083 59035
rect 13139 58979 13225 59035
rect 13281 58979 13367 59035
rect 13423 58979 13509 59035
rect 13565 58979 13651 59035
rect 13707 58979 13793 59035
rect 13849 58979 13935 59035
rect 13991 58979 14077 59035
rect 14133 58979 14219 59035
rect 14275 58979 14361 59035
rect 14417 58979 14503 59035
rect 14559 58979 14645 59035
rect 14701 58979 14787 59035
rect 14843 58979 14853 59035
rect 151 58893 14853 58979
rect 151 58837 161 58893
rect 217 58837 303 58893
rect 359 58837 445 58893
rect 501 58837 587 58893
rect 643 58837 729 58893
rect 785 58837 871 58893
rect 927 58837 1013 58893
rect 1069 58837 1155 58893
rect 1211 58837 1297 58893
rect 1353 58837 1439 58893
rect 1495 58837 1581 58893
rect 1637 58837 1723 58893
rect 1779 58837 1865 58893
rect 1921 58837 2007 58893
rect 2063 58837 2149 58893
rect 2205 58837 2291 58893
rect 2347 58837 2433 58893
rect 2489 58837 2575 58893
rect 2631 58837 2717 58893
rect 2773 58837 2859 58893
rect 2915 58837 3001 58893
rect 3057 58837 3143 58893
rect 3199 58837 3285 58893
rect 3341 58837 3427 58893
rect 3483 58837 3569 58893
rect 3625 58837 3711 58893
rect 3767 58837 3853 58893
rect 3909 58837 3995 58893
rect 4051 58837 4137 58893
rect 4193 58837 4279 58893
rect 4335 58837 4421 58893
rect 4477 58837 4563 58893
rect 4619 58837 4705 58893
rect 4761 58837 4847 58893
rect 4903 58837 4989 58893
rect 5045 58837 5131 58893
rect 5187 58837 5273 58893
rect 5329 58837 5415 58893
rect 5471 58837 5557 58893
rect 5613 58837 5699 58893
rect 5755 58837 5841 58893
rect 5897 58837 5983 58893
rect 6039 58837 6125 58893
rect 6181 58837 6267 58893
rect 6323 58837 6409 58893
rect 6465 58837 6551 58893
rect 6607 58837 6693 58893
rect 6749 58837 6835 58893
rect 6891 58837 6977 58893
rect 7033 58837 7119 58893
rect 7175 58837 7261 58893
rect 7317 58837 7403 58893
rect 7459 58837 7545 58893
rect 7601 58837 7687 58893
rect 7743 58837 7829 58893
rect 7885 58837 7971 58893
rect 8027 58837 8113 58893
rect 8169 58837 8255 58893
rect 8311 58837 8397 58893
rect 8453 58837 8539 58893
rect 8595 58837 8681 58893
rect 8737 58837 8823 58893
rect 8879 58837 8965 58893
rect 9021 58837 9107 58893
rect 9163 58837 9249 58893
rect 9305 58837 9391 58893
rect 9447 58837 9533 58893
rect 9589 58837 9675 58893
rect 9731 58837 9817 58893
rect 9873 58837 9959 58893
rect 10015 58837 10101 58893
rect 10157 58837 10243 58893
rect 10299 58837 10385 58893
rect 10441 58837 10527 58893
rect 10583 58837 10669 58893
rect 10725 58837 10811 58893
rect 10867 58837 10953 58893
rect 11009 58837 11095 58893
rect 11151 58837 11237 58893
rect 11293 58837 11379 58893
rect 11435 58837 11521 58893
rect 11577 58837 11663 58893
rect 11719 58837 11805 58893
rect 11861 58837 11947 58893
rect 12003 58837 12089 58893
rect 12145 58837 12231 58893
rect 12287 58837 12373 58893
rect 12429 58837 12515 58893
rect 12571 58837 12657 58893
rect 12713 58837 12799 58893
rect 12855 58837 12941 58893
rect 12997 58837 13083 58893
rect 13139 58837 13225 58893
rect 13281 58837 13367 58893
rect 13423 58837 13509 58893
rect 13565 58837 13651 58893
rect 13707 58837 13793 58893
rect 13849 58837 13935 58893
rect 13991 58837 14077 58893
rect 14133 58837 14219 58893
rect 14275 58837 14361 58893
rect 14417 58837 14503 58893
rect 14559 58837 14645 58893
rect 14701 58837 14787 58893
rect 14843 58837 14853 58893
rect 151 58827 14853 58837
rect 151 58563 14853 58573
rect 151 58507 161 58563
rect 217 58507 303 58563
rect 359 58507 445 58563
rect 501 58507 587 58563
rect 643 58507 729 58563
rect 785 58507 871 58563
rect 927 58507 1013 58563
rect 1069 58507 1155 58563
rect 1211 58507 1297 58563
rect 1353 58507 1439 58563
rect 1495 58507 1581 58563
rect 1637 58507 1723 58563
rect 1779 58507 1865 58563
rect 1921 58507 2007 58563
rect 2063 58507 2149 58563
rect 2205 58507 2291 58563
rect 2347 58507 2433 58563
rect 2489 58507 2575 58563
rect 2631 58507 2717 58563
rect 2773 58507 2859 58563
rect 2915 58507 3001 58563
rect 3057 58507 3143 58563
rect 3199 58507 3285 58563
rect 3341 58507 3427 58563
rect 3483 58507 3569 58563
rect 3625 58507 3711 58563
rect 3767 58507 3853 58563
rect 3909 58507 3995 58563
rect 4051 58507 4137 58563
rect 4193 58507 4279 58563
rect 4335 58507 4421 58563
rect 4477 58507 4563 58563
rect 4619 58507 4705 58563
rect 4761 58507 4847 58563
rect 4903 58507 4989 58563
rect 5045 58507 5131 58563
rect 5187 58507 5273 58563
rect 5329 58507 5415 58563
rect 5471 58507 5557 58563
rect 5613 58507 5699 58563
rect 5755 58507 5841 58563
rect 5897 58507 5983 58563
rect 6039 58507 6125 58563
rect 6181 58507 6267 58563
rect 6323 58507 6409 58563
rect 6465 58507 6551 58563
rect 6607 58507 6693 58563
rect 6749 58507 6835 58563
rect 6891 58507 6977 58563
rect 7033 58507 7119 58563
rect 7175 58507 7261 58563
rect 7317 58507 7403 58563
rect 7459 58507 7545 58563
rect 7601 58507 7687 58563
rect 7743 58507 7829 58563
rect 7885 58507 7971 58563
rect 8027 58507 8113 58563
rect 8169 58507 8255 58563
rect 8311 58507 8397 58563
rect 8453 58507 8539 58563
rect 8595 58507 8681 58563
rect 8737 58507 8823 58563
rect 8879 58507 8965 58563
rect 9021 58507 9107 58563
rect 9163 58507 9249 58563
rect 9305 58507 9391 58563
rect 9447 58507 9533 58563
rect 9589 58507 9675 58563
rect 9731 58507 9817 58563
rect 9873 58507 9959 58563
rect 10015 58507 10101 58563
rect 10157 58507 10243 58563
rect 10299 58507 10385 58563
rect 10441 58507 10527 58563
rect 10583 58507 10669 58563
rect 10725 58507 10811 58563
rect 10867 58507 10953 58563
rect 11009 58507 11095 58563
rect 11151 58507 11237 58563
rect 11293 58507 11379 58563
rect 11435 58507 11521 58563
rect 11577 58507 11663 58563
rect 11719 58507 11805 58563
rect 11861 58507 11947 58563
rect 12003 58507 12089 58563
rect 12145 58507 12231 58563
rect 12287 58507 12373 58563
rect 12429 58507 12515 58563
rect 12571 58507 12657 58563
rect 12713 58507 12799 58563
rect 12855 58507 12941 58563
rect 12997 58507 13083 58563
rect 13139 58507 13225 58563
rect 13281 58507 13367 58563
rect 13423 58507 13509 58563
rect 13565 58507 13651 58563
rect 13707 58507 13793 58563
rect 13849 58507 13935 58563
rect 13991 58507 14077 58563
rect 14133 58507 14219 58563
rect 14275 58507 14361 58563
rect 14417 58507 14503 58563
rect 14559 58507 14645 58563
rect 14701 58507 14787 58563
rect 14843 58507 14853 58563
rect 151 58421 14853 58507
rect 151 58365 161 58421
rect 217 58365 303 58421
rect 359 58365 445 58421
rect 501 58365 587 58421
rect 643 58365 729 58421
rect 785 58365 871 58421
rect 927 58365 1013 58421
rect 1069 58365 1155 58421
rect 1211 58365 1297 58421
rect 1353 58365 1439 58421
rect 1495 58365 1581 58421
rect 1637 58365 1723 58421
rect 1779 58365 1865 58421
rect 1921 58365 2007 58421
rect 2063 58365 2149 58421
rect 2205 58365 2291 58421
rect 2347 58365 2433 58421
rect 2489 58365 2575 58421
rect 2631 58365 2717 58421
rect 2773 58365 2859 58421
rect 2915 58365 3001 58421
rect 3057 58365 3143 58421
rect 3199 58365 3285 58421
rect 3341 58365 3427 58421
rect 3483 58365 3569 58421
rect 3625 58365 3711 58421
rect 3767 58365 3853 58421
rect 3909 58365 3995 58421
rect 4051 58365 4137 58421
rect 4193 58365 4279 58421
rect 4335 58365 4421 58421
rect 4477 58365 4563 58421
rect 4619 58365 4705 58421
rect 4761 58365 4847 58421
rect 4903 58365 4989 58421
rect 5045 58365 5131 58421
rect 5187 58365 5273 58421
rect 5329 58365 5415 58421
rect 5471 58365 5557 58421
rect 5613 58365 5699 58421
rect 5755 58365 5841 58421
rect 5897 58365 5983 58421
rect 6039 58365 6125 58421
rect 6181 58365 6267 58421
rect 6323 58365 6409 58421
rect 6465 58365 6551 58421
rect 6607 58365 6693 58421
rect 6749 58365 6835 58421
rect 6891 58365 6977 58421
rect 7033 58365 7119 58421
rect 7175 58365 7261 58421
rect 7317 58365 7403 58421
rect 7459 58365 7545 58421
rect 7601 58365 7687 58421
rect 7743 58365 7829 58421
rect 7885 58365 7971 58421
rect 8027 58365 8113 58421
rect 8169 58365 8255 58421
rect 8311 58365 8397 58421
rect 8453 58365 8539 58421
rect 8595 58365 8681 58421
rect 8737 58365 8823 58421
rect 8879 58365 8965 58421
rect 9021 58365 9107 58421
rect 9163 58365 9249 58421
rect 9305 58365 9391 58421
rect 9447 58365 9533 58421
rect 9589 58365 9675 58421
rect 9731 58365 9817 58421
rect 9873 58365 9959 58421
rect 10015 58365 10101 58421
rect 10157 58365 10243 58421
rect 10299 58365 10385 58421
rect 10441 58365 10527 58421
rect 10583 58365 10669 58421
rect 10725 58365 10811 58421
rect 10867 58365 10953 58421
rect 11009 58365 11095 58421
rect 11151 58365 11237 58421
rect 11293 58365 11379 58421
rect 11435 58365 11521 58421
rect 11577 58365 11663 58421
rect 11719 58365 11805 58421
rect 11861 58365 11947 58421
rect 12003 58365 12089 58421
rect 12145 58365 12231 58421
rect 12287 58365 12373 58421
rect 12429 58365 12515 58421
rect 12571 58365 12657 58421
rect 12713 58365 12799 58421
rect 12855 58365 12941 58421
rect 12997 58365 13083 58421
rect 13139 58365 13225 58421
rect 13281 58365 13367 58421
rect 13423 58365 13509 58421
rect 13565 58365 13651 58421
rect 13707 58365 13793 58421
rect 13849 58365 13935 58421
rect 13991 58365 14077 58421
rect 14133 58365 14219 58421
rect 14275 58365 14361 58421
rect 14417 58365 14503 58421
rect 14559 58365 14645 58421
rect 14701 58365 14787 58421
rect 14843 58365 14853 58421
rect 151 58279 14853 58365
rect 151 58223 161 58279
rect 217 58223 303 58279
rect 359 58223 445 58279
rect 501 58223 587 58279
rect 643 58223 729 58279
rect 785 58223 871 58279
rect 927 58223 1013 58279
rect 1069 58223 1155 58279
rect 1211 58223 1297 58279
rect 1353 58223 1439 58279
rect 1495 58223 1581 58279
rect 1637 58223 1723 58279
rect 1779 58223 1865 58279
rect 1921 58223 2007 58279
rect 2063 58223 2149 58279
rect 2205 58223 2291 58279
rect 2347 58223 2433 58279
rect 2489 58223 2575 58279
rect 2631 58223 2717 58279
rect 2773 58223 2859 58279
rect 2915 58223 3001 58279
rect 3057 58223 3143 58279
rect 3199 58223 3285 58279
rect 3341 58223 3427 58279
rect 3483 58223 3569 58279
rect 3625 58223 3711 58279
rect 3767 58223 3853 58279
rect 3909 58223 3995 58279
rect 4051 58223 4137 58279
rect 4193 58223 4279 58279
rect 4335 58223 4421 58279
rect 4477 58223 4563 58279
rect 4619 58223 4705 58279
rect 4761 58223 4847 58279
rect 4903 58223 4989 58279
rect 5045 58223 5131 58279
rect 5187 58223 5273 58279
rect 5329 58223 5415 58279
rect 5471 58223 5557 58279
rect 5613 58223 5699 58279
rect 5755 58223 5841 58279
rect 5897 58223 5983 58279
rect 6039 58223 6125 58279
rect 6181 58223 6267 58279
rect 6323 58223 6409 58279
rect 6465 58223 6551 58279
rect 6607 58223 6693 58279
rect 6749 58223 6835 58279
rect 6891 58223 6977 58279
rect 7033 58223 7119 58279
rect 7175 58223 7261 58279
rect 7317 58223 7403 58279
rect 7459 58223 7545 58279
rect 7601 58223 7687 58279
rect 7743 58223 7829 58279
rect 7885 58223 7971 58279
rect 8027 58223 8113 58279
rect 8169 58223 8255 58279
rect 8311 58223 8397 58279
rect 8453 58223 8539 58279
rect 8595 58223 8681 58279
rect 8737 58223 8823 58279
rect 8879 58223 8965 58279
rect 9021 58223 9107 58279
rect 9163 58223 9249 58279
rect 9305 58223 9391 58279
rect 9447 58223 9533 58279
rect 9589 58223 9675 58279
rect 9731 58223 9817 58279
rect 9873 58223 9959 58279
rect 10015 58223 10101 58279
rect 10157 58223 10243 58279
rect 10299 58223 10385 58279
rect 10441 58223 10527 58279
rect 10583 58223 10669 58279
rect 10725 58223 10811 58279
rect 10867 58223 10953 58279
rect 11009 58223 11095 58279
rect 11151 58223 11237 58279
rect 11293 58223 11379 58279
rect 11435 58223 11521 58279
rect 11577 58223 11663 58279
rect 11719 58223 11805 58279
rect 11861 58223 11947 58279
rect 12003 58223 12089 58279
rect 12145 58223 12231 58279
rect 12287 58223 12373 58279
rect 12429 58223 12515 58279
rect 12571 58223 12657 58279
rect 12713 58223 12799 58279
rect 12855 58223 12941 58279
rect 12997 58223 13083 58279
rect 13139 58223 13225 58279
rect 13281 58223 13367 58279
rect 13423 58223 13509 58279
rect 13565 58223 13651 58279
rect 13707 58223 13793 58279
rect 13849 58223 13935 58279
rect 13991 58223 14077 58279
rect 14133 58223 14219 58279
rect 14275 58223 14361 58279
rect 14417 58223 14503 58279
rect 14559 58223 14645 58279
rect 14701 58223 14787 58279
rect 14843 58223 14853 58279
rect 151 58137 14853 58223
rect 151 58081 161 58137
rect 217 58081 303 58137
rect 359 58081 445 58137
rect 501 58081 587 58137
rect 643 58081 729 58137
rect 785 58081 871 58137
rect 927 58081 1013 58137
rect 1069 58081 1155 58137
rect 1211 58081 1297 58137
rect 1353 58081 1439 58137
rect 1495 58081 1581 58137
rect 1637 58081 1723 58137
rect 1779 58081 1865 58137
rect 1921 58081 2007 58137
rect 2063 58081 2149 58137
rect 2205 58081 2291 58137
rect 2347 58081 2433 58137
rect 2489 58081 2575 58137
rect 2631 58081 2717 58137
rect 2773 58081 2859 58137
rect 2915 58081 3001 58137
rect 3057 58081 3143 58137
rect 3199 58081 3285 58137
rect 3341 58081 3427 58137
rect 3483 58081 3569 58137
rect 3625 58081 3711 58137
rect 3767 58081 3853 58137
rect 3909 58081 3995 58137
rect 4051 58081 4137 58137
rect 4193 58081 4279 58137
rect 4335 58081 4421 58137
rect 4477 58081 4563 58137
rect 4619 58081 4705 58137
rect 4761 58081 4847 58137
rect 4903 58081 4989 58137
rect 5045 58081 5131 58137
rect 5187 58081 5273 58137
rect 5329 58081 5415 58137
rect 5471 58081 5557 58137
rect 5613 58081 5699 58137
rect 5755 58081 5841 58137
rect 5897 58081 5983 58137
rect 6039 58081 6125 58137
rect 6181 58081 6267 58137
rect 6323 58081 6409 58137
rect 6465 58081 6551 58137
rect 6607 58081 6693 58137
rect 6749 58081 6835 58137
rect 6891 58081 6977 58137
rect 7033 58081 7119 58137
rect 7175 58081 7261 58137
rect 7317 58081 7403 58137
rect 7459 58081 7545 58137
rect 7601 58081 7687 58137
rect 7743 58081 7829 58137
rect 7885 58081 7971 58137
rect 8027 58081 8113 58137
rect 8169 58081 8255 58137
rect 8311 58081 8397 58137
rect 8453 58081 8539 58137
rect 8595 58081 8681 58137
rect 8737 58081 8823 58137
rect 8879 58081 8965 58137
rect 9021 58081 9107 58137
rect 9163 58081 9249 58137
rect 9305 58081 9391 58137
rect 9447 58081 9533 58137
rect 9589 58081 9675 58137
rect 9731 58081 9817 58137
rect 9873 58081 9959 58137
rect 10015 58081 10101 58137
rect 10157 58081 10243 58137
rect 10299 58081 10385 58137
rect 10441 58081 10527 58137
rect 10583 58081 10669 58137
rect 10725 58081 10811 58137
rect 10867 58081 10953 58137
rect 11009 58081 11095 58137
rect 11151 58081 11237 58137
rect 11293 58081 11379 58137
rect 11435 58081 11521 58137
rect 11577 58081 11663 58137
rect 11719 58081 11805 58137
rect 11861 58081 11947 58137
rect 12003 58081 12089 58137
rect 12145 58081 12231 58137
rect 12287 58081 12373 58137
rect 12429 58081 12515 58137
rect 12571 58081 12657 58137
rect 12713 58081 12799 58137
rect 12855 58081 12941 58137
rect 12997 58081 13083 58137
rect 13139 58081 13225 58137
rect 13281 58081 13367 58137
rect 13423 58081 13509 58137
rect 13565 58081 13651 58137
rect 13707 58081 13793 58137
rect 13849 58081 13935 58137
rect 13991 58081 14077 58137
rect 14133 58081 14219 58137
rect 14275 58081 14361 58137
rect 14417 58081 14503 58137
rect 14559 58081 14645 58137
rect 14701 58081 14787 58137
rect 14843 58081 14853 58137
rect 151 57995 14853 58081
rect 151 57939 161 57995
rect 217 57939 303 57995
rect 359 57939 445 57995
rect 501 57939 587 57995
rect 643 57939 729 57995
rect 785 57939 871 57995
rect 927 57939 1013 57995
rect 1069 57939 1155 57995
rect 1211 57939 1297 57995
rect 1353 57939 1439 57995
rect 1495 57939 1581 57995
rect 1637 57939 1723 57995
rect 1779 57939 1865 57995
rect 1921 57939 2007 57995
rect 2063 57939 2149 57995
rect 2205 57939 2291 57995
rect 2347 57939 2433 57995
rect 2489 57939 2575 57995
rect 2631 57939 2717 57995
rect 2773 57939 2859 57995
rect 2915 57939 3001 57995
rect 3057 57939 3143 57995
rect 3199 57939 3285 57995
rect 3341 57939 3427 57995
rect 3483 57939 3569 57995
rect 3625 57939 3711 57995
rect 3767 57939 3853 57995
rect 3909 57939 3995 57995
rect 4051 57939 4137 57995
rect 4193 57939 4279 57995
rect 4335 57939 4421 57995
rect 4477 57939 4563 57995
rect 4619 57939 4705 57995
rect 4761 57939 4847 57995
rect 4903 57939 4989 57995
rect 5045 57939 5131 57995
rect 5187 57939 5273 57995
rect 5329 57939 5415 57995
rect 5471 57939 5557 57995
rect 5613 57939 5699 57995
rect 5755 57939 5841 57995
rect 5897 57939 5983 57995
rect 6039 57939 6125 57995
rect 6181 57939 6267 57995
rect 6323 57939 6409 57995
rect 6465 57939 6551 57995
rect 6607 57939 6693 57995
rect 6749 57939 6835 57995
rect 6891 57939 6977 57995
rect 7033 57939 7119 57995
rect 7175 57939 7261 57995
rect 7317 57939 7403 57995
rect 7459 57939 7545 57995
rect 7601 57939 7687 57995
rect 7743 57939 7829 57995
rect 7885 57939 7971 57995
rect 8027 57939 8113 57995
rect 8169 57939 8255 57995
rect 8311 57939 8397 57995
rect 8453 57939 8539 57995
rect 8595 57939 8681 57995
rect 8737 57939 8823 57995
rect 8879 57939 8965 57995
rect 9021 57939 9107 57995
rect 9163 57939 9249 57995
rect 9305 57939 9391 57995
rect 9447 57939 9533 57995
rect 9589 57939 9675 57995
rect 9731 57939 9817 57995
rect 9873 57939 9959 57995
rect 10015 57939 10101 57995
rect 10157 57939 10243 57995
rect 10299 57939 10385 57995
rect 10441 57939 10527 57995
rect 10583 57939 10669 57995
rect 10725 57939 10811 57995
rect 10867 57939 10953 57995
rect 11009 57939 11095 57995
rect 11151 57939 11237 57995
rect 11293 57939 11379 57995
rect 11435 57939 11521 57995
rect 11577 57939 11663 57995
rect 11719 57939 11805 57995
rect 11861 57939 11947 57995
rect 12003 57939 12089 57995
rect 12145 57939 12231 57995
rect 12287 57939 12373 57995
rect 12429 57939 12515 57995
rect 12571 57939 12657 57995
rect 12713 57939 12799 57995
rect 12855 57939 12941 57995
rect 12997 57939 13083 57995
rect 13139 57939 13225 57995
rect 13281 57939 13367 57995
rect 13423 57939 13509 57995
rect 13565 57939 13651 57995
rect 13707 57939 13793 57995
rect 13849 57939 13935 57995
rect 13991 57939 14077 57995
rect 14133 57939 14219 57995
rect 14275 57939 14361 57995
rect 14417 57939 14503 57995
rect 14559 57939 14645 57995
rect 14701 57939 14787 57995
rect 14843 57939 14853 57995
rect 151 57853 14853 57939
rect 151 57797 161 57853
rect 217 57797 303 57853
rect 359 57797 445 57853
rect 501 57797 587 57853
rect 643 57797 729 57853
rect 785 57797 871 57853
rect 927 57797 1013 57853
rect 1069 57797 1155 57853
rect 1211 57797 1297 57853
rect 1353 57797 1439 57853
rect 1495 57797 1581 57853
rect 1637 57797 1723 57853
rect 1779 57797 1865 57853
rect 1921 57797 2007 57853
rect 2063 57797 2149 57853
rect 2205 57797 2291 57853
rect 2347 57797 2433 57853
rect 2489 57797 2575 57853
rect 2631 57797 2717 57853
rect 2773 57797 2859 57853
rect 2915 57797 3001 57853
rect 3057 57797 3143 57853
rect 3199 57797 3285 57853
rect 3341 57797 3427 57853
rect 3483 57797 3569 57853
rect 3625 57797 3711 57853
rect 3767 57797 3853 57853
rect 3909 57797 3995 57853
rect 4051 57797 4137 57853
rect 4193 57797 4279 57853
rect 4335 57797 4421 57853
rect 4477 57797 4563 57853
rect 4619 57797 4705 57853
rect 4761 57797 4847 57853
rect 4903 57797 4989 57853
rect 5045 57797 5131 57853
rect 5187 57797 5273 57853
rect 5329 57797 5415 57853
rect 5471 57797 5557 57853
rect 5613 57797 5699 57853
rect 5755 57797 5841 57853
rect 5897 57797 5983 57853
rect 6039 57797 6125 57853
rect 6181 57797 6267 57853
rect 6323 57797 6409 57853
rect 6465 57797 6551 57853
rect 6607 57797 6693 57853
rect 6749 57797 6835 57853
rect 6891 57797 6977 57853
rect 7033 57797 7119 57853
rect 7175 57797 7261 57853
rect 7317 57797 7403 57853
rect 7459 57797 7545 57853
rect 7601 57797 7687 57853
rect 7743 57797 7829 57853
rect 7885 57797 7971 57853
rect 8027 57797 8113 57853
rect 8169 57797 8255 57853
rect 8311 57797 8397 57853
rect 8453 57797 8539 57853
rect 8595 57797 8681 57853
rect 8737 57797 8823 57853
rect 8879 57797 8965 57853
rect 9021 57797 9107 57853
rect 9163 57797 9249 57853
rect 9305 57797 9391 57853
rect 9447 57797 9533 57853
rect 9589 57797 9675 57853
rect 9731 57797 9817 57853
rect 9873 57797 9959 57853
rect 10015 57797 10101 57853
rect 10157 57797 10243 57853
rect 10299 57797 10385 57853
rect 10441 57797 10527 57853
rect 10583 57797 10669 57853
rect 10725 57797 10811 57853
rect 10867 57797 10953 57853
rect 11009 57797 11095 57853
rect 11151 57797 11237 57853
rect 11293 57797 11379 57853
rect 11435 57797 11521 57853
rect 11577 57797 11663 57853
rect 11719 57797 11805 57853
rect 11861 57797 11947 57853
rect 12003 57797 12089 57853
rect 12145 57797 12231 57853
rect 12287 57797 12373 57853
rect 12429 57797 12515 57853
rect 12571 57797 12657 57853
rect 12713 57797 12799 57853
rect 12855 57797 12941 57853
rect 12997 57797 13083 57853
rect 13139 57797 13225 57853
rect 13281 57797 13367 57853
rect 13423 57797 13509 57853
rect 13565 57797 13651 57853
rect 13707 57797 13793 57853
rect 13849 57797 13935 57853
rect 13991 57797 14077 57853
rect 14133 57797 14219 57853
rect 14275 57797 14361 57853
rect 14417 57797 14503 57853
rect 14559 57797 14645 57853
rect 14701 57797 14787 57853
rect 14843 57797 14853 57853
rect 151 57711 14853 57797
rect 151 57655 161 57711
rect 217 57655 303 57711
rect 359 57655 445 57711
rect 501 57655 587 57711
rect 643 57655 729 57711
rect 785 57655 871 57711
rect 927 57655 1013 57711
rect 1069 57655 1155 57711
rect 1211 57655 1297 57711
rect 1353 57655 1439 57711
rect 1495 57655 1581 57711
rect 1637 57655 1723 57711
rect 1779 57655 1865 57711
rect 1921 57655 2007 57711
rect 2063 57655 2149 57711
rect 2205 57655 2291 57711
rect 2347 57655 2433 57711
rect 2489 57655 2575 57711
rect 2631 57655 2717 57711
rect 2773 57655 2859 57711
rect 2915 57655 3001 57711
rect 3057 57655 3143 57711
rect 3199 57655 3285 57711
rect 3341 57655 3427 57711
rect 3483 57655 3569 57711
rect 3625 57655 3711 57711
rect 3767 57655 3853 57711
rect 3909 57655 3995 57711
rect 4051 57655 4137 57711
rect 4193 57655 4279 57711
rect 4335 57655 4421 57711
rect 4477 57655 4563 57711
rect 4619 57655 4705 57711
rect 4761 57655 4847 57711
rect 4903 57655 4989 57711
rect 5045 57655 5131 57711
rect 5187 57655 5273 57711
rect 5329 57655 5415 57711
rect 5471 57655 5557 57711
rect 5613 57655 5699 57711
rect 5755 57655 5841 57711
rect 5897 57655 5983 57711
rect 6039 57655 6125 57711
rect 6181 57655 6267 57711
rect 6323 57655 6409 57711
rect 6465 57655 6551 57711
rect 6607 57655 6693 57711
rect 6749 57655 6835 57711
rect 6891 57655 6977 57711
rect 7033 57655 7119 57711
rect 7175 57655 7261 57711
rect 7317 57655 7403 57711
rect 7459 57655 7545 57711
rect 7601 57655 7687 57711
rect 7743 57655 7829 57711
rect 7885 57655 7971 57711
rect 8027 57655 8113 57711
rect 8169 57655 8255 57711
rect 8311 57655 8397 57711
rect 8453 57655 8539 57711
rect 8595 57655 8681 57711
rect 8737 57655 8823 57711
rect 8879 57655 8965 57711
rect 9021 57655 9107 57711
rect 9163 57655 9249 57711
rect 9305 57655 9391 57711
rect 9447 57655 9533 57711
rect 9589 57655 9675 57711
rect 9731 57655 9817 57711
rect 9873 57655 9959 57711
rect 10015 57655 10101 57711
rect 10157 57655 10243 57711
rect 10299 57655 10385 57711
rect 10441 57655 10527 57711
rect 10583 57655 10669 57711
rect 10725 57655 10811 57711
rect 10867 57655 10953 57711
rect 11009 57655 11095 57711
rect 11151 57655 11237 57711
rect 11293 57655 11379 57711
rect 11435 57655 11521 57711
rect 11577 57655 11663 57711
rect 11719 57655 11805 57711
rect 11861 57655 11947 57711
rect 12003 57655 12089 57711
rect 12145 57655 12231 57711
rect 12287 57655 12373 57711
rect 12429 57655 12515 57711
rect 12571 57655 12657 57711
rect 12713 57655 12799 57711
rect 12855 57655 12941 57711
rect 12997 57655 13083 57711
rect 13139 57655 13225 57711
rect 13281 57655 13367 57711
rect 13423 57655 13509 57711
rect 13565 57655 13651 57711
rect 13707 57655 13793 57711
rect 13849 57655 13935 57711
rect 13991 57655 14077 57711
rect 14133 57655 14219 57711
rect 14275 57655 14361 57711
rect 14417 57655 14503 57711
rect 14559 57655 14645 57711
rect 14701 57655 14787 57711
rect 14843 57655 14853 57711
rect 151 57569 14853 57655
rect 151 57513 161 57569
rect 217 57513 303 57569
rect 359 57513 445 57569
rect 501 57513 587 57569
rect 643 57513 729 57569
rect 785 57513 871 57569
rect 927 57513 1013 57569
rect 1069 57513 1155 57569
rect 1211 57513 1297 57569
rect 1353 57513 1439 57569
rect 1495 57513 1581 57569
rect 1637 57513 1723 57569
rect 1779 57513 1865 57569
rect 1921 57513 2007 57569
rect 2063 57513 2149 57569
rect 2205 57513 2291 57569
rect 2347 57513 2433 57569
rect 2489 57513 2575 57569
rect 2631 57513 2717 57569
rect 2773 57513 2859 57569
rect 2915 57513 3001 57569
rect 3057 57513 3143 57569
rect 3199 57513 3285 57569
rect 3341 57513 3427 57569
rect 3483 57513 3569 57569
rect 3625 57513 3711 57569
rect 3767 57513 3853 57569
rect 3909 57513 3995 57569
rect 4051 57513 4137 57569
rect 4193 57513 4279 57569
rect 4335 57513 4421 57569
rect 4477 57513 4563 57569
rect 4619 57513 4705 57569
rect 4761 57513 4847 57569
rect 4903 57513 4989 57569
rect 5045 57513 5131 57569
rect 5187 57513 5273 57569
rect 5329 57513 5415 57569
rect 5471 57513 5557 57569
rect 5613 57513 5699 57569
rect 5755 57513 5841 57569
rect 5897 57513 5983 57569
rect 6039 57513 6125 57569
rect 6181 57513 6267 57569
rect 6323 57513 6409 57569
rect 6465 57513 6551 57569
rect 6607 57513 6693 57569
rect 6749 57513 6835 57569
rect 6891 57513 6977 57569
rect 7033 57513 7119 57569
rect 7175 57513 7261 57569
rect 7317 57513 7403 57569
rect 7459 57513 7545 57569
rect 7601 57513 7687 57569
rect 7743 57513 7829 57569
rect 7885 57513 7971 57569
rect 8027 57513 8113 57569
rect 8169 57513 8255 57569
rect 8311 57513 8397 57569
rect 8453 57513 8539 57569
rect 8595 57513 8681 57569
rect 8737 57513 8823 57569
rect 8879 57513 8965 57569
rect 9021 57513 9107 57569
rect 9163 57513 9249 57569
rect 9305 57513 9391 57569
rect 9447 57513 9533 57569
rect 9589 57513 9675 57569
rect 9731 57513 9817 57569
rect 9873 57513 9959 57569
rect 10015 57513 10101 57569
rect 10157 57513 10243 57569
rect 10299 57513 10385 57569
rect 10441 57513 10527 57569
rect 10583 57513 10669 57569
rect 10725 57513 10811 57569
rect 10867 57513 10953 57569
rect 11009 57513 11095 57569
rect 11151 57513 11237 57569
rect 11293 57513 11379 57569
rect 11435 57513 11521 57569
rect 11577 57513 11663 57569
rect 11719 57513 11805 57569
rect 11861 57513 11947 57569
rect 12003 57513 12089 57569
rect 12145 57513 12231 57569
rect 12287 57513 12373 57569
rect 12429 57513 12515 57569
rect 12571 57513 12657 57569
rect 12713 57513 12799 57569
rect 12855 57513 12941 57569
rect 12997 57513 13083 57569
rect 13139 57513 13225 57569
rect 13281 57513 13367 57569
rect 13423 57513 13509 57569
rect 13565 57513 13651 57569
rect 13707 57513 13793 57569
rect 13849 57513 13935 57569
rect 13991 57513 14077 57569
rect 14133 57513 14219 57569
rect 14275 57513 14361 57569
rect 14417 57513 14503 57569
rect 14559 57513 14645 57569
rect 14701 57513 14787 57569
rect 14843 57513 14853 57569
rect 151 57427 14853 57513
rect 151 57371 161 57427
rect 217 57371 303 57427
rect 359 57371 445 57427
rect 501 57371 587 57427
rect 643 57371 729 57427
rect 785 57371 871 57427
rect 927 57371 1013 57427
rect 1069 57371 1155 57427
rect 1211 57371 1297 57427
rect 1353 57371 1439 57427
rect 1495 57371 1581 57427
rect 1637 57371 1723 57427
rect 1779 57371 1865 57427
rect 1921 57371 2007 57427
rect 2063 57371 2149 57427
rect 2205 57371 2291 57427
rect 2347 57371 2433 57427
rect 2489 57371 2575 57427
rect 2631 57371 2717 57427
rect 2773 57371 2859 57427
rect 2915 57371 3001 57427
rect 3057 57371 3143 57427
rect 3199 57371 3285 57427
rect 3341 57371 3427 57427
rect 3483 57371 3569 57427
rect 3625 57371 3711 57427
rect 3767 57371 3853 57427
rect 3909 57371 3995 57427
rect 4051 57371 4137 57427
rect 4193 57371 4279 57427
rect 4335 57371 4421 57427
rect 4477 57371 4563 57427
rect 4619 57371 4705 57427
rect 4761 57371 4847 57427
rect 4903 57371 4989 57427
rect 5045 57371 5131 57427
rect 5187 57371 5273 57427
rect 5329 57371 5415 57427
rect 5471 57371 5557 57427
rect 5613 57371 5699 57427
rect 5755 57371 5841 57427
rect 5897 57371 5983 57427
rect 6039 57371 6125 57427
rect 6181 57371 6267 57427
rect 6323 57371 6409 57427
rect 6465 57371 6551 57427
rect 6607 57371 6693 57427
rect 6749 57371 6835 57427
rect 6891 57371 6977 57427
rect 7033 57371 7119 57427
rect 7175 57371 7261 57427
rect 7317 57371 7403 57427
rect 7459 57371 7545 57427
rect 7601 57371 7687 57427
rect 7743 57371 7829 57427
rect 7885 57371 7971 57427
rect 8027 57371 8113 57427
rect 8169 57371 8255 57427
rect 8311 57371 8397 57427
rect 8453 57371 8539 57427
rect 8595 57371 8681 57427
rect 8737 57371 8823 57427
rect 8879 57371 8965 57427
rect 9021 57371 9107 57427
rect 9163 57371 9249 57427
rect 9305 57371 9391 57427
rect 9447 57371 9533 57427
rect 9589 57371 9675 57427
rect 9731 57371 9817 57427
rect 9873 57371 9959 57427
rect 10015 57371 10101 57427
rect 10157 57371 10243 57427
rect 10299 57371 10385 57427
rect 10441 57371 10527 57427
rect 10583 57371 10669 57427
rect 10725 57371 10811 57427
rect 10867 57371 10953 57427
rect 11009 57371 11095 57427
rect 11151 57371 11237 57427
rect 11293 57371 11379 57427
rect 11435 57371 11521 57427
rect 11577 57371 11663 57427
rect 11719 57371 11805 57427
rect 11861 57371 11947 57427
rect 12003 57371 12089 57427
rect 12145 57371 12231 57427
rect 12287 57371 12373 57427
rect 12429 57371 12515 57427
rect 12571 57371 12657 57427
rect 12713 57371 12799 57427
rect 12855 57371 12941 57427
rect 12997 57371 13083 57427
rect 13139 57371 13225 57427
rect 13281 57371 13367 57427
rect 13423 57371 13509 57427
rect 13565 57371 13651 57427
rect 13707 57371 13793 57427
rect 13849 57371 13935 57427
rect 13991 57371 14077 57427
rect 14133 57371 14219 57427
rect 14275 57371 14361 57427
rect 14417 57371 14503 57427
rect 14559 57371 14645 57427
rect 14701 57371 14787 57427
rect 14843 57371 14853 57427
rect 151 57285 14853 57371
rect 151 57229 161 57285
rect 217 57229 303 57285
rect 359 57229 445 57285
rect 501 57229 587 57285
rect 643 57229 729 57285
rect 785 57229 871 57285
rect 927 57229 1013 57285
rect 1069 57229 1155 57285
rect 1211 57229 1297 57285
rect 1353 57229 1439 57285
rect 1495 57229 1581 57285
rect 1637 57229 1723 57285
rect 1779 57229 1865 57285
rect 1921 57229 2007 57285
rect 2063 57229 2149 57285
rect 2205 57229 2291 57285
rect 2347 57229 2433 57285
rect 2489 57229 2575 57285
rect 2631 57229 2717 57285
rect 2773 57229 2859 57285
rect 2915 57229 3001 57285
rect 3057 57229 3143 57285
rect 3199 57229 3285 57285
rect 3341 57229 3427 57285
rect 3483 57229 3569 57285
rect 3625 57229 3711 57285
rect 3767 57229 3853 57285
rect 3909 57229 3995 57285
rect 4051 57229 4137 57285
rect 4193 57229 4279 57285
rect 4335 57229 4421 57285
rect 4477 57229 4563 57285
rect 4619 57229 4705 57285
rect 4761 57229 4847 57285
rect 4903 57229 4989 57285
rect 5045 57229 5131 57285
rect 5187 57229 5273 57285
rect 5329 57229 5415 57285
rect 5471 57229 5557 57285
rect 5613 57229 5699 57285
rect 5755 57229 5841 57285
rect 5897 57229 5983 57285
rect 6039 57229 6125 57285
rect 6181 57229 6267 57285
rect 6323 57229 6409 57285
rect 6465 57229 6551 57285
rect 6607 57229 6693 57285
rect 6749 57229 6835 57285
rect 6891 57229 6977 57285
rect 7033 57229 7119 57285
rect 7175 57229 7261 57285
rect 7317 57229 7403 57285
rect 7459 57229 7545 57285
rect 7601 57229 7687 57285
rect 7743 57229 7829 57285
rect 7885 57229 7971 57285
rect 8027 57229 8113 57285
rect 8169 57229 8255 57285
rect 8311 57229 8397 57285
rect 8453 57229 8539 57285
rect 8595 57229 8681 57285
rect 8737 57229 8823 57285
rect 8879 57229 8965 57285
rect 9021 57229 9107 57285
rect 9163 57229 9249 57285
rect 9305 57229 9391 57285
rect 9447 57229 9533 57285
rect 9589 57229 9675 57285
rect 9731 57229 9817 57285
rect 9873 57229 9959 57285
rect 10015 57229 10101 57285
rect 10157 57229 10243 57285
rect 10299 57229 10385 57285
rect 10441 57229 10527 57285
rect 10583 57229 10669 57285
rect 10725 57229 10811 57285
rect 10867 57229 10953 57285
rect 11009 57229 11095 57285
rect 11151 57229 11237 57285
rect 11293 57229 11379 57285
rect 11435 57229 11521 57285
rect 11577 57229 11663 57285
rect 11719 57229 11805 57285
rect 11861 57229 11947 57285
rect 12003 57229 12089 57285
rect 12145 57229 12231 57285
rect 12287 57229 12373 57285
rect 12429 57229 12515 57285
rect 12571 57229 12657 57285
rect 12713 57229 12799 57285
rect 12855 57229 12941 57285
rect 12997 57229 13083 57285
rect 13139 57229 13225 57285
rect 13281 57229 13367 57285
rect 13423 57229 13509 57285
rect 13565 57229 13651 57285
rect 13707 57229 13793 57285
rect 13849 57229 13935 57285
rect 13991 57229 14077 57285
rect 14133 57229 14219 57285
rect 14275 57229 14361 57285
rect 14417 57229 14503 57285
rect 14559 57229 14645 57285
rect 14701 57229 14787 57285
rect 14843 57229 14853 57285
rect 151 57219 14853 57229
rect 151 56971 14853 56981
rect 151 56915 161 56971
rect 217 56915 303 56971
rect 359 56915 445 56971
rect 501 56915 587 56971
rect 643 56915 729 56971
rect 785 56915 871 56971
rect 927 56915 1013 56971
rect 1069 56915 1155 56971
rect 1211 56915 1297 56971
rect 1353 56915 1439 56971
rect 1495 56915 1581 56971
rect 1637 56915 1723 56971
rect 1779 56915 1865 56971
rect 1921 56915 2007 56971
rect 2063 56915 2149 56971
rect 2205 56915 2291 56971
rect 2347 56915 2433 56971
rect 2489 56915 2575 56971
rect 2631 56915 2717 56971
rect 2773 56915 2859 56971
rect 2915 56915 3001 56971
rect 3057 56915 3143 56971
rect 3199 56915 3285 56971
rect 3341 56915 3427 56971
rect 3483 56915 3569 56971
rect 3625 56915 3711 56971
rect 3767 56915 3853 56971
rect 3909 56915 3995 56971
rect 4051 56915 4137 56971
rect 4193 56915 4279 56971
rect 4335 56915 4421 56971
rect 4477 56915 4563 56971
rect 4619 56915 4705 56971
rect 4761 56915 4847 56971
rect 4903 56915 4989 56971
rect 5045 56915 5131 56971
rect 5187 56915 5273 56971
rect 5329 56915 5415 56971
rect 5471 56915 5557 56971
rect 5613 56915 5699 56971
rect 5755 56915 5841 56971
rect 5897 56915 5983 56971
rect 6039 56915 6125 56971
rect 6181 56915 6267 56971
rect 6323 56915 6409 56971
rect 6465 56915 6551 56971
rect 6607 56915 6693 56971
rect 6749 56915 6835 56971
rect 6891 56915 6977 56971
rect 7033 56915 7119 56971
rect 7175 56915 7261 56971
rect 7317 56915 7403 56971
rect 7459 56915 7545 56971
rect 7601 56915 7687 56971
rect 7743 56915 7829 56971
rect 7885 56915 7971 56971
rect 8027 56915 8113 56971
rect 8169 56915 8255 56971
rect 8311 56915 8397 56971
rect 8453 56915 8539 56971
rect 8595 56915 8681 56971
rect 8737 56915 8823 56971
rect 8879 56915 8965 56971
rect 9021 56915 9107 56971
rect 9163 56915 9249 56971
rect 9305 56915 9391 56971
rect 9447 56915 9533 56971
rect 9589 56915 9675 56971
rect 9731 56915 9817 56971
rect 9873 56915 9959 56971
rect 10015 56915 10101 56971
rect 10157 56915 10243 56971
rect 10299 56915 10385 56971
rect 10441 56915 10527 56971
rect 10583 56915 10669 56971
rect 10725 56915 10811 56971
rect 10867 56915 10953 56971
rect 11009 56915 11095 56971
rect 11151 56915 11237 56971
rect 11293 56915 11379 56971
rect 11435 56915 11521 56971
rect 11577 56915 11663 56971
rect 11719 56915 11805 56971
rect 11861 56915 11947 56971
rect 12003 56915 12089 56971
rect 12145 56915 12231 56971
rect 12287 56915 12373 56971
rect 12429 56915 12515 56971
rect 12571 56915 12657 56971
rect 12713 56915 12799 56971
rect 12855 56915 12941 56971
rect 12997 56915 13083 56971
rect 13139 56915 13225 56971
rect 13281 56915 13367 56971
rect 13423 56915 13509 56971
rect 13565 56915 13651 56971
rect 13707 56915 13793 56971
rect 13849 56915 13935 56971
rect 13991 56915 14077 56971
rect 14133 56915 14219 56971
rect 14275 56915 14361 56971
rect 14417 56915 14503 56971
rect 14559 56915 14645 56971
rect 14701 56915 14787 56971
rect 14843 56915 14853 56971
rect 151 56829 14853 56915
rect 151 56773 161 56829
rect 217 56773 303 56829
rect 359 56773 445 56829
rect 501 56773 587 56829
rect 643 56773 729 56829
rect 785 56773 871 56829
rect 927 56773 1013 56829
rect 1069 56773 1155 56829
rect 1211 56773 1297 56829
rect 1353 56773 1439 56829
rect 1495 56773 1581 56829
rect 1637 56773 1723 56829
rect 1779 56773 1865 56829
rect 1921 56773 2007 56829
rect 2063 56773 2149 56829
rect 2205 56773 2291 56829
rect 2347 56773 2433 56829
rect 2489 56773 2575 56829
rect 2631 56773 2717 56829
rect 2773 56773 2859 56829
rect 2915 56773 3001 56829
rect 3057 56773 3143 56829
rect 3199 56773 3285 56829
rect 3341 56773 3427 56829
rect 3483 56773 3569 56829
rect 3625 56773 3711 56829
rect 3767 56773 3853 56829
rect 3909 56773 3995 56829
rect 4051 56773 4137 56829
rect 4193 56773 4279 56829
rect 4335 56773 4421 56829
rect 4477 56773 4563 56829
rect 4619 56773 4705 56829
rect 4761 56773 4847 56829
rect 4903 56773 4989 56829
rect 5045 56773 5131 56829
rect 5187 56773 5273 56829
rect 5329 56773 5415 56829
rect 5471 56773 5557 56829
rect 5613 56773 5699 56829
rect 5755 56773 5841 56829
rect 5897 56773 5983 56829
rect 6039 56773 6125 56829
rect 6181 56773 6267 56829
rect 6323 56773 6409 56829
rect 6465 56773 6551 56829
rect 6607 56773 6693 56829
rect 6749 56773 6835 56829
rect 6891 56773 6977 56829
rect 7033 56773 7119 56829
rect 7175 56773 7261 56829
rect 7317 56773 7403 56829
rect 7459 56773 7545 56829
rect 7601 56773 7687 56829
rect 7743 56773 7829 56829
rect 7885 56773 7971 56829
rect 8027 56773 8113 56829
rect 8169 56773 8255 56829
rect 8311 56773 8397 56829
rect 8453 56773 8539 56829
rect 8595 56773 8681 56829
rect 8737 56773 8823 56829
rect 8879 56773 8965 56829
rect 9021 56773 9107 56829
rect 9163 56773 9249 56829
rect 9305 56773 9391 56829
rect 9447 56773 9533 56829
rect 9589 56773 9675 56829
rect 9731 56773 9817 56829
rect 9873 56773 9959 56829
rect 10015 56773 10101 56829
rect 10157 56773 10243 56829
rect 10299 56773 10385 56829
rect 10441 56773 10527 56829
rect 10583 56773 10669 56829
rect 10725 56773 10811 56829
rect 10867 56773 10953 56829
rect 11009 56773 11095 56829
rect 11151 56773 11237 56829
rect 11293 56773 11379 56829
rect 11435 56773 11521 56829
rect 11577 56773 11663 56829
rect 11719 56773 11805 56829
rect 11861 56773 11947 56829
rect 12003 56773 12089 56829
rect 12145 56773 12231 56829
rect 12287 56773 12373 56829
rect 12429 56773 12515 56829
rect 12571 56773 12657 56829
rect 12713 56773 12799 56829
rect 12855 56773 12941 56829
rect 12997 56773 13083 56829
rect 13139 56773 13225 56829
rect 13281 56773 13367 56829
rect 13423 56773 13509 56829
rect 13565 56773 13651 56829
rect 13707 56773 13793 56829
rect 13849 56773 13935 56829
rect 13991 56773 14077 56829
rect 14133 56773 14219 56829
rect 14275 56773 14361 56829
rect 14417 56773 14503 56829
rect 14559 56773 14645 56829
rect 14701 56773 14787 56829
rect 14843 56773 14853 56829
rect 151 56687 14853 56773
rect 151 56631 161 56687
rect 217 56631 303 56687
rect 359 56631 445 56687
rect 501 56631 587 56687
rect 643 56631 729 56687
rect 785 56631 871 56687
rect 927 56631 1013 56687
rect 1069 56631 1155 56687
rect 1211 56631 1297 56687
rect 1353 56631 1439 56687
rect 1495 56631 1581 56687
rect 1637 56631 1723 56687
rect 1779 56631 1865 56687
rect 1921 56631 2007 56687
rect 2063 56631 2149 56687
rect 2205 56631 2291 56687
rect 2347 56631 2433 56687
rect 2489 56631 2575 56687
rect 2631 56631 2717 56687
rect 2773 56631 2859 56687
rect 2915 56631 3001 56687
rect 3057 56631 3143 56687
rect 3199 56631 3285 56687
rect 3341 56631 3427 56687
rect 3483 56631 3569 56687
rect 3625 56631 3711 56687
rect 3767 56631 3853 56687
rect 3909 56631 3995 56687
rect 4051 56631 4137 56687
rect 4193 56631 4279 56687
rect 4335 56631 4421 56687
rect 4477 56631 4563 56687
rect 4619 56631 4705 56687
rect 4761 56631 4847 56687
rect 4903 56631 4989 56687
rect 5045 56631 5131 56687
rect 5187 56631 5273 56687
rect 5329 56631 5415 56687
rect 5471 56631 5557 56687
rect 5613 56631 5699 56687
rect 5755 56631 5841 56687
rect 5897 56631 5983 56687
rect 6039 56631 6125 56687
rect 6181 56631 6267 56687
rect 6323 56631 6409 56687
rect 6465 56631 6551 56687
rect 6607 56631 6693 56687
rect 6749 56631 6835 56687
rect 6891 56631 6977 56687
rect 7033 56631 7119 56687
rect 7175 56631 7261 56687
rect 7317 56631 7403 56687
rect 7459 56631 7545 56687
rect 7601 56631 7687 56687
rect 7743 56631 7829 56687
rect 7885 56631 7971 56687
rect 8027 56631 8113 56687
rect 8169 56631 8255 56687
rect 8311 56631 8397 56687
rect 8453 56631 8539 56687
rect 8595 56631 8681 56687
rect 8737 56631 8823 56687
rect 8879 56631 8965 56687
rect 9021 56631 9107 56687
rect 9163 56631 9249 56687
rect 9305 56631 9391 56687
rect 9447 56631 9533 56687
rect 9589 56631 9675 56687
rect 9731 56631 9817 56687
rect 9873 56631 9959 56687
rect 10015 56631 10101 56687
rect 10157 56631 10243 56687
rect 10299 56631 10385 56687
rect 10441 56631 10527 56687
rect 10583 56631 10669 56687
rect 10725 56631 10811 56687
rect 10867 56631 10953 56687
rect 11009 56631 11095 56687
rect 11151 56631 11237 56687
rect 11293 56631 11379 56687
rect 11435 56631 11521 56687
rect 11577 56631 11663 56687
rect 11719 56631 11805 56687
rect 11861 56631 11947 56687
rect 12003 56631 12089 56687
rect 12145 56631 12231 56687
rect 12287 56631 12373 56687
rect 12429 56631 12515 56687
rect 12571 56631 12657 56687
rect 12713 56631 12799 56687
rect 12855 56631 12941 56687
rect 12997 56631 13083 56687
rect 13139 56631 13225 56687
rect 13281 56631 13367 56687
rect 13423 56631 13509 56687
rect 13565 56631 13651 56687
rect 13707 56631 13793 56687
rect 13849 56631 13935 56687
rect 13991 56631 14077 56687
rect 14133 56631 14219 56687
rect 14275 56631 14361 56687
rect 14417 56631 14503 56687
rect 14559 56631 14645 56687
rect 14701 56631 14787 56687
rect 14843 56631 14853 56687
rect 151 56545 14853 56631
rect 151 56489 161 56545
rect 217 56489 303 56545
rect 359 56489 445 56545
rect 501 56489 587 56545
rect 643 56489 729 56545
rect 785 56489 871 56545
rect 927 56489 1013 56545
rect 1069 56489 1155 56545
rect 1211 56489 1297 56545
rect 1353 56489 1439 56545
rect 1495 56489 1581 56545
rect 1637 56489 1723 56545
rect 1779 56489 1865 56545
rect 1921 56489 2007 56545
rect 2063 56489 2149 56545
rect 2205 56489 2291 56545
rect 2347 56489 2433 56545
rect 2489 56489 2575 56545
rect 2631 56489 2717 56545
rect 2773 56489 2859 56545
rect 2915 56489 3001 56545
rect 3057 56489 3143 56545
rect 3199 56489 3285 56545
rect 3341 56489 3427 56545
rect 3483 56489 3569 56545
rect 3625 56489 3711 56545
rect 3767 56489 3853 56545
rect 3909 56489 3995 56545
rect 4051 56489 4137 56545
rect 4193 56489 4279 56545
rect 4335 56489 4421 56545
rect 4477 56489 4563 56545
rect 4619 56489 4705 56545
rect 4761 56489 4847 56545
rect 4903 56489 4989 56545
rect 5045 56489 5131 56545
rect 5187 56489 5273 56545
rect 5329 56489 5415 56545
rect 5471 56489 5557 56545
rect 5613 56489 5699 56545
rect 5755 56489 5841 56545
rect 5897 56489 5983 56545
rect 6039 56489 6125 56545
rect 6181 56489 6267 56545
rect 6323 56489 6409 56545
rect 6465 56489 6551 56545
rect 6607 56489 6693 56545
rect 6749 56489 6835 56545
rect 6891 56489 6977 56545
rect 7033 56489 7119 56545
rect 7175 56489 7261 56545
rect 7317 56489 7403 56545
rect 7459 56489 7545 56545
rect 7601 56489 7687 56545
rect 7743 56489 7829 56545
rect 7885 56489 7971 56545
rect 8027 56489 8113 56545
rect 8169 56489 8255 56545
rect 8311 56489 8397 56545
rect 8453 56489 8539 56545
rect 8595 56489 8681 56545
rect 8737 56489 8823 56545
rect 8879 56489 8965 56545
rect 9021 56489 9107 56545
rect 9163 56489 9249 56545
rect 9305 56489 9391 56545
rect 9447 56489 9533 56545
rect 9589 56489 9675 56545
rect 9731 56489 9817 56545
rect 9873 56489 9959 56545
rect 10015 56489 10101 56545
rect 10157 56489 10243 56545
rect 10299 56489 10385 56545
rect 10441 56489 10527 56545
rect 10583 56489 10669 56545
rect 10725 56489 10811 56545
rect 10867 56489 10953 56545
rect 11009 56489 11095 56545
rect 11151 56489 11237 56545
rect 11293 56489 11379 56545
rect 11435 56489 11521 56545
rect 11577 56489 11663 56545
rect 11719 56489 11805 56545
rect 11861 56489 11947 56545
rect 12003 56489 12089 56545
rect 12145 56489 12231 56545
rect 12287 56489 12373 56545
rect 12429 56489 12515 56545
rect 12571 56489 12657 56545
rect 12713 56489 12799 56545
rect 12855 56489 12941 56545
rect 12997 56489 13083 56545
rect 13139 56489 13225 56545
rect 13281 56489 13367 56545
rect 13423 56489 13509 56545
rect 13565 56489 13651 56545
rect 13707 56489 13793 56545
rect 13849 56489 13935 56545
rect 13991 56489 14077 56545
rect 14133 56489 14219 56545
rect 14275 56489 14361 56545
rect 14417 56489 14503 56545
rect 14559 56489 14645 56545
rect 14701 56489 14787 56545
rect 14843 56489 14853 56545
rect 151 56403 14853 56489
rect 151 56347 161 56403
rect 217 56347 303 56403
rect 359 56347 445 56403
rect 501 56347 587 56403
rect 643 56347 729 56403
rect 785 56347 871 56403
rect 927 56347 1013 56403
rect 1069 56347 1155 56403
rect 1211 56347 1297 56403
rect 1353 56347 1439 56403
rect 1495 56347 1581 56403
rect 1637 56347 1723 56403
rect 1779 56347 1865 56403
rect 1921 56347 2007 56403
rect 2063 56347 2149 56403
rect 2205 56347 2291 56403
rect 2347 56347 2433 56403
rect 2489 56347 2575 56403
rect 2631 56347 2717 56403
rect 2773 56347 2859 56403
rect 2915 56347 3001 56403
rect 3057 56347 3143 56403
rect 3199 56347 3285 56403
rect 3341 56347 3427 56403
rect 3483 56347 3569 56403
rect 3625 56347 3711 56403
rect 3767 56347 3853 56403
rect 3909 56347 3995 56403
rect 4051 56347 4137 56403
rect 4193 56347 4279 56403
rect 4335 56347 4421 56403
rect 4477 56347 4563 56403
rect 4619 56347 4705 56403
rect 4761 56347 4847 56403
rect 4903 56347 4989 56403
rect 5045 56347 5131 56403
rect 5187 56347 5273 56403
rect 5329 56347 5415 56403
rect 5471 56347 5557 56403
rect 5613 56347 5699 56403
rect 5755 56347 5841 56403
rect 5897 56347 5983 56403
rect 6039 56347 6125 56403
rect 6181 56347 6267 56403
rect 6323 56347 6409 56403
rect 6465 56347 6551 56403
rect 6607 56347 6693 56403
rect 6749 56347 6835 56403
rect 6891 56347 6977 56403
rect 7033 56347 7119 56403
rect 7175 56347 7261 56403
rect 7317 56347 7403 56403
rect 7459 56347 7545 56403
rect 7601 56347 7687 56403
rect 7743 56347 7829 56403
rect 7885 56347 7971 56403
rect 8027 56347 8113 56403
rect 8169 56347 8255 56403
rect 8311 56347 8397 56403
rect 8453 56347 8539 56403
rect 8595 56347 8681 56403
rect 8737 56347 8823 56403
rect 8879 56347 8965 56403
rect 9021 56347 9107 56403
rect 9163 56347 9249 56403
rect 9305 56347 9391 56403
rect 9447 56347 9533 56403
rect 9589 56347 9675 56403
rect 9731 56347 9817 56403
rect 9873 56347 9959 56403
rect 10015 56347 10101 56403
rect 10157 56347 10243 56403
rect 10299 56347 10385 56403
rect 10441 56347 10527 56403
rect 10583 56347 10669 56403
rect 10725 56347 10811 56403
rect 10867 56347 10953 56403
rect 11009 56347 11095 56403
rect 11151 56347 11237 56403
rect 11293 56347 11379 56403
rect 11435 56347 11521 56403
rect 11577 56347 11663 56403
rect 11719 56347 11805 56403
rect 11861 56347 11947 56403
rect 12003 56347 12089 56403
rect 12145 56347 12231 56403
rect 12287 56347 12373 56403
rect 12429 56347 12515 56403
rect 12571 56347 12657 56403
rect 12713 56347 12799 56403
rect 12855 56347 12941 56403
rect 12997 56347 13083 56403
rect 13139 56347 13225 56403
rect 13281 56347 13367 56403
rect 13423 56347 13509 56403
rect 13565 56347 13651 56403
rect 13707 56347 13793 56403
rect 13849 56347 13935 56403
rect 13991 56347 14077 56403
rect 14133 56347 14219 56403
rect 14275 56347 14361 56403
rect 14417 56347 14503 56403
rect 14559 56347 14645 56403
rect 14701 56347 14787 56403
rect 14843 56347 14853 56403
rect 151 56261 14853 56347
rect 151 56205 161 56261
rect 217 56205 303 56261
rect 359 56205 445 56261
rect 501 56205 587 56261
rect 643 56205 729 56261
rect 785 56205 871 56261
rect 927 56205 1013 56261
rect 1069 56205 1155 56261
rect 1211 56205 1297 56261
rect 1353 56205 1439 56261
rect 1495 56205 1581 56261
rect 1637 56205 1723 56261
rect 1779 56205 1865 56261
rect 1921 56205 2007 56261
rect 2063 56205 2149 56261
rect 2205 56205 2291 56261
rect 2347 56205 2433 56261
rect 2489 56205 2575 56261
rect 2631 56205 2717 56261
rect 2773 56205 2859 56261
rect 2915 56205 3001 56261
rect 3057 56205 3143 56261
rect 3199 56205 3285 56261
rect 3341 56205 3427 56261
rect 3483 56205 3569 56261
rect 3625 56205 3711 56261
rect 3767 56205 3853 56261
rect 3909 56205 3995 56261
rect 4051 56205 4137 56261
rect 4193 56205 4279 56261
rect 4335 56205 4421 56261
rect 4477 56205 4563 56261
rect 4619 56205 4705 56261
rect 4761 56205 4847 56261
rect 4903 56205 4989 56261
rect 5045 56205 5131 56261
rect 5187 56205 5273 56261
rect 5329 56205 5415 56261
rect 5471 56205 5557 56261
rect 5613 56205 5699 56261
rect 5755 56205 5841 56261
rect 5897 56205 5983 56261
rect 6039 56205 6125 56261
rect 6181 56205 6267 56261
rect 6323 56205 6409 56261
rect 6465 56205 6551 56261
rect 6607 56205 6693 56261
rect 6749 56205 6835 56261
rect 6891 56205 6977 56261
rect 7033 56205 7119 56261
rect 7175 56205 7261 56261
rect 7317 56205 7403 56261
rect 7459 56205 7545 56261
rect 7601 56205 7687 56261
rect 7743 56205 7829 56261
rect 7885 56205 7971 56261
rect 8027 56205 8113 56261
rect 8169 56205 8255 56261
rect 8311 56205 8397 56261
rect 8453 56205 8539 56261
rect 8595 56205 8681 56261
rect 8737 56205 8823 56261
rect 8879 56205 8965 56261
rect 9021 56205 9107 56261
rect 9163 56205 9249 56261
rect 9305 56205 9391 56261
rect 9447 56205 9533 56261
rect 9589 56205 9675 56261
rect 9731 56205 9817 56261
rect 9873 56205 9959 56261
rect 10015 56205 10101 56261
rect 10157 56205 10243 56261
rect 10299 56205 10385 56261
rect 10441 56205 10527 56261
rect 10583 56205 10669 56261
rect 10725 56205 10811 56261
rect 10867 56205 10953 56261
rect 11009 56205 11095 56261
rect 11151 56205 11237 56261
rect 11293 56205 11379 56261
rect 11435 56205 11521 56261
rect 11577 56205 11663 56261
rect 11719 56205 11805 56261
rect 11861 56205 11947 56261
rect 12003 56205 12089 56261
rect 12145 56205 12231 56261
rect 12287 56205 12373 56261
rect 12429 56205 12515 56261
rect 12571 56205 12657 56261
rect 12713 56205 12799 56261
rect 12855 56205 12941 56261
rect 12997 56205 13083 56261
rect 13139 56205 13225 56261
rect 13281 56205 13367 56261
rect 13423 56205 13509 56261
rect 13565 56205 13651 56261
rect 13707 56205 13793 56261
rect 13849 56205 13935 56261
rect 13991 56205 14077 56261
rect 14133 56205 14219 56261
rect 14275 56205 14361 56261
rect 14417 56205 14503 56261
rect 14559 56205 14645 56261
rect 14701 56205 14787 56261
rect 14843 56205 14853 56261
rect 151 56119 14853 56205
rect 151 56063 161 56119
rect 217 56063 303 56119
rect 359 56063 445 56119
rect 501 56063 587 56119
rect 643 56063 729 56119
rect 785 56063 871 56119
rect 927 56063 1013 56119
rect 1069 56063 1155 56119
rect 1211 56063 1297 56119
rect 1353 56063 1439 56119
rect 1495 56063 1581 56119
rect 1637 56063 1723 56119
rect 1779 56063 1865 56119
rect 1921 56063 2007 56119
rect 2063 56063 2149 56119
rect 2205 56063 2291 56119
rect 2347 56063 2433 56119
rect 2489 56063 2575 56119
rect 2631 56063 2717 56119
rect 2773 56063 2859 56119
rect 2915 56063 3001 56119
rect 3057 56063 3143 56119
rect 3199 56063 3285 56119
rect 3341 56063 3427 56119
rect 3483 56063 3569 56119
rect 3625 56063 3711 56119
rect 3767 56063 3853 56119
rect 3909 56063 3995 56119
rect 4051 56063 4137 56119
rect 4193 56063 4279 56119
rect 4335 56063 4421 56119
rect 4477 56063 4563 56119
rect 4619 56063 4705 56119
rect 4761 56063 4847 56119
rect 4903 56063 4989 56119
rect 5045 56063 5131 56119
rect 5187 56063 5273 56119
rect 5329 56063 5415 56119
rect 5471 56063 5557 56119
rect 5613 56063 5699 56119
rect 5755 56063 5841 56119
rect 5897 56063 5983 56119
rect 6039 56063 6125 56119
rect 6181 56063 6267 56119
rect 6323 56063 6409 56119
rect 6465 56063 6551 56119
rect 6607 56063 6693 56119
rect 6749 56063 6835 56119
rect 6891 56063 6977 56119
rect 7033 56063 7119 56119
rect 7175 56063 7261 56119
rect 7317 56063 7403 56119
rect 7459 56063 7545 56119
rect 7601 56063 7687 56119
rect 7743 56063 7829 56119
rect 7885 56063 7971 56119
rect 8027 56063 8113 56119
rect 8169 56063 8255 56119
rect 8311 56063 8397 56119
rect 8453 56063 8539 56119
rect 8595 56063 8681 56119
rect 8737 56063 8823 56119
rect 8879 56063 8965 56119
rect 9021 56063 9107 56119
rect 9163 56063 9249 56119
rect 9305 56063 9391 56119
rect 9447 56063 9533 56119
rect 9589 56063 9675 56119
rect 9731 56063 9817 56119
rect 9873 56063 9959 56119
rect 10015 56063 10101 56119
rect 10157 56063 10243 56119
rect 10299 56063 10385 56119
rect 10441 56063 10527 56119
rect 10583 56063 10669 56119
rect 10725 56063 10811 56119
rect 10867 56063 10953 56119
rect 11009 56063 11095 56119
rect 11151 56063 11237 56119
rect 11293 56063 11379 56119
rect 11435 56063 11521 56119
rect 11577 56063 11663 56119
rect 11719 56063 11805 56119
rect 11861 56063 11947 56119
rect 12003 56063 12089 56119
rect 12145 56063 12231 56119
rect 12287 56063 12373 56119
rect 12429 56063 12515 56119
rect 12571 56063 12657 56119
rect 12713 56063 12799 56119
rect 12855 56063 12941 56119
rect 12997 56063 13083 56119
rect 13139 56063 13225 56119
rect 13281 56063 13367 56119
rect 13423 56063 13509 56119
rect 13565 56063 13651 56119
rect 13707 56063 13793 56119
rect 13849 56063 13935 56119
rect 13991 56063 14077 56119
rect 14133 56063 14219 56119
rect 14275 56063 14361 56119
rect 14417 56063 14503 56119
rect 14559 56063 14645 56119
rect 14701 56063 14787 56119
rect 14843 56063 14853 56119
rect 151 55977 14853 56063
rect 151 55921 161 55977
rect 217 55921 303 55977
rect 359 55921 445 55977
rect 501 55921 587 55977
rect 643 55921 729 55977
rect 785 55921 871 55977
rect 927 55921 1013 55977
rect 1069 55921 1155 55977
rect 1211 55921 1297 55977
rect 1353 55921 1439 55977
rect 1495 55921 1581 55977
rect 1637 55921 1723 55977
rect 1779 55921 1865 55977
rect 1921 55921 2007 55977
rect 2063 55921 2149 55977
rect 2205 55921 2291 55977
rect 2347 55921 2433 55977
rect 2489 55921 2575 55977
rect 2631 55921 2717 55977
rect 2773 55921 2859 55977
rect 2915 55921 3001 55977
rect 3057 55921 3143 55977
rect 3199 55921 3285 55977
rect 3341 55921 3427 55977
rect 3483 55921 3569 55977
rect 3625 55921 3711 55977
rect 3767 55921 3853 55977
rect 3909 55921 3995 55977
rect 4051 55921 4137 55977
rect 4193 55921 4279 55977
rect 4335 55921 4421 55977
rect 4477 55921 4563 55977
rect 4619 55921 4705 55977
rect 4761 55921 4847 55977
rect 4903 55921 4989 55977
rect 5045 55921 5131 55977
rect 5187 55921 5273 55977
rect 5329 55921 5415 55977
rect 5471 55921 5557 55977
rect 5613 55921 5699 55977
rect 5755 55921 5841 55977
rect 5897 55921 5983 55977
rect 6039 55921 6125 55977
rect 6181 55921 6267 55977
rect 6323 55921 6409 55977
rect 6465 55921 6551 55977
rect 6607 55921 6693 55977
rect 6749 55921 6835 55977
rect 6891 55921 6977 55977
rect 7033 55921 7119 55977
rect 7175 55921 7261 55977
rect 7317 55921 7403 55977
rect 7459 55921 7545 55977
rect 7601 55921 7687 55977
rect 7743 55921 7829 55977
rect 7885 55921 7971 55977
rect 8027 55921 8113 55977
rect 8169 55921 8255 55977
rect 8311 55921 8397 55977
rect 8453 55921 8539 55977
rect 8595 55921 8681 55977
rect 8737 55921 8823 55977
rect 8879 55921 8965 55977
rect 9021 55921 9107 55977
rect 9163 55921 9249 55977
rect 9305 55921 9391 55977
rect 9447 55921 9533 55977
rect 9589 55921 9675 55977
rect 9731 55921 9817 55977
rect 9873 55921 9959 55977
rect 10015 55921 10101 55977
rect 10157 55921 10243 55977
rect 10299 55921 10385 55977
rect 10441 55921 10527 55977
rect 10583 55921 10669 55977
rect 10725 55921 10811 55977
rect 10867 55921 10953 55977
rect 11009 55921 11095 55977
rect 11151 55921 11237 55977
rect 11293 55921 11379 55977
rect 11435 55921 11521 55977
rect 11577 55921 11663 55977
rect 11719 55921 11805 55977
rect 11861 55921 11947 55977
rect 12003 55921 12089 55977
rect 12145 55921 12231 55977
rect 12287 55921 12373 55977
rect 12429 55921 12515 55977
rect 12571 55921 12657 55977
rect 12713 55921 12799 55977
rect 12855 55921 12941 55977
rect 12997 55921 13083 55977
rect 13139 55921 13225 55977
rect 13281 55921 13367 55977
rect 13423 55921 13509 55977
rect 13565 55921 13651 55977
rect 13707 55921 13793 55977
rect 13849 55921 13935 55977
rect 13991 55921 14077 55977
rect 14133 55921 14219 55977
rect 14275 55921 14361 55977
rect 14417 55921 14503 55977
rect 14559 55921 14645 55977
rect 14701 55921 14787 55977
rect 14843 55921 14853 55977
rect 151 55835 14853 55921
rect 151 55779 161 55835
rect 217 55779 303 55835
rect 359 55779 445 55835
rect 501 55779 587 55835
rect 643 55779 729 55835
rect 785 55779 871 55835
rect 927 55779 1013 55835
rect 1069 55779 1155 55835
rect 1211 55779 1297 55835
rect 1353 55779 1439 55835
rect 1495 55779 1581 55835
rect 1637 55779 1723 55835
rect 1779 55779 1865 55835
rect 1921 55779 2007 55835
rect 2063 55779 2149 55835
rect 2205 55779 2291 55835
rect 2347 55779 2433 55835
rect 2489 55779 2575 55835
rect 2631 55779 2717 55835
rect 2773 55779 2859 55835
rect 2915 55779 3001 55835
rect 3057 55779 3143 55835
rect 3199 55779 3285 55835
rect 3341 55779 3427 55835
rect 3483 55779 3569 55835
rect 3625 55779 3711 55835
rect 3767 55779 3853 55835
rect 3909 55779 3995 55835
rect 4051 55779 4137 55835
rect 4193 55779 4279 55835
rect 4335 55779 4421 55835
rect 4477 55779 4563 55835
rect 4619 55779 4705 55835
rect 4761 55779 4847 55835
rect 4903 55779 4989 55835
rect 5045 55779 5131 55835
rect 5187 55779 5273 55835
rect 5329 55779 5415 55835
rect 5471 55779 5557 55835
rect 5613 55779 5699 55835
rect 5755 55779 5841 55835
rect 5897 55779 5983 55835
rect 6039 55779 6125 55835
rect 6181 55779 6267 55835
rect 6323 55779 6409 55835
rect 6465 55779 6551 55835
rect 6607 55779 6693 55835
rect 6749 55779 6835 55835
rect 6891 55779 6977 55835
rect 7033 55779 7119 55835
rect 7175 55779 7261 55835
rect 7317 55779 7403 55835
rect 7459 55779 7545 55835
rect 7601 55779 7687 55835
rect 7743 55779 7829 55835
rect 7885 55779 7971 55835
rect 8027 55779 8113 55835
rect 8169 55779 8255 55835
rect 8311 55779 8397 55835
rect 8453 55779 8539 55835
rect 8595 55779 8681 55835
rect 8737 55779 8823 55835
rect 8879 55779 8965 55835
rect 9021 55779 9107 55835
rect 9163 55779 9249 55835
rect 9305 55779 9391 55835
rect 9447 55779 9533 55835
rect 9589 55779 9675 55835
rect 9731 55779 9817 55835
rect 9873 55779 9959 55835
rect 10015 55779 10101 55835
rect 10157 55779 10243 55835
rect 10299 55779 10385 55835
rect 10441 55779 10527 55835
rect 10583 55779 10669 55835
rect 10725 55779 10811 55835
rect 10867 55779 10953 55835
rect 11009 55779 11095 55835
rect 11151 55779 11237 55835
rect 11293 55779 11379 55835
rect 11435 55779 11521 55835
rect 11577 55779 11663 55835
rect 11719 55779 11805 55835
rect 11861 55779 11947 55835
rect 12003 55779 12089 55835
rect 12145 55779 12231 55835
rect 12287 55779 12373 55835
rect 12429 55779 12515 55835
rect 12571 55779 12657 55835
rect 12713 55779 12799 55835
rect 12855 55779 12941 55835
rect 12997 55779 13083 55835
rect 13139 55779 13225 55835
rect 13281 55779 13367 55835
rect 13423 55779 13509 55835
rect 13565 55779 13651 55835
rect 13707 55779 13793 55835
rect 13849 55779 13935 55835
rect 13991 55779 14077 55835
rect 14133 55779 14219 55835
rect 14275 55779 14361 55835
rect 14417 55779 14503 55835
rect 14559 55779 14645 55835
rect 14701 55779 14787 55835
rect 14843 55779 14853 55835
rect 151 55693 14853 55779
rect 151 55637 161 55693
rect 217 55637 303 55693
rect 359 55637 445 55693
rect 501 55637 587 55693
rect 643 55637 729 55693
rect 785 55637 871 55693
rect 927 55637 1013 55693
rect 1069 55637 1155 55693
rect 1211 55637 1297 55693
rect 1353 55637 1439 55693
rect 1495 55637 1581 55693
rect 1637 55637 1723 55693
rect 1779 55637 1865 55693
rect 1921 55637 2007 55693
rect 2063 55637 2149 55693
rect 2205 55637 2291 55693
rect 2347 55637 2433 55693
rect 2489 55637 2575 55693
rect 2631 55637 2717 55693
rect 2773 55637 2859 55693
rect 2915 55637 3001 55693
rect 3057 55637 3143 55693
rect 3199 55637 3285 55693
rect 3341 55637 3427 55693
rect 3483 55637 3569 55693
rect 3625 55637 3711 55693
rect 3767 55637 3853 55693
rect 3909 55637 3995 55693
rect 4051 55637 4137 55693
rect 4193 55637 4279 55693
rect 4335 55637 4421 55693
rect 4477 55637 4563 55693
rect 4619 55637 4705 55693
rect 4761 55637 4847 55693
rect 4903 55637 4989 55693
rect 5045 55637 5131 55693
rect 5187 55637 5273 55693
rect 5329 55637 5415 55693
rect 5471 55637 5557 55693
rect 5613 55637 5699 55693
rect 5755 55637 5841 55693
rect 5897 55637 5983 55693
rect 6039 55637 6125 55693
rect 6181 55637 6267 55693
rect 6323 55637 6409 55693
rect 6465 55637 6551 55693
rect 6607 55637 6693 55693
rect 6749 55637 6835 55693
rect 6891 55637 6977 55693
rect 7033 55637 7119 55693
rect 7175 55637 7261 55693
rect 7317 55637 7403 55693
rect 7459 55637 7545 55693
rect 7601 55637 7687 55693
rect 7743 55637 7829 55693
rect 7885 55637 7971 55693
rect 8027 55637 8113 55693
rect 8169 55637 8255 55693
rect 8311 55637 8397 55693
rect 8453 55637 8539 55693
rect 8595 55637 8681 55693
rect 8737 55637 8823 55693
rect 8879 55637 8965 55693
rect 9021 55637 9107 55693
rect 9163 55637 9249 55693
rect 9305 55637 9391 55693
rect 9447 55637 9533 55693
rect 9589 55637 9675 55693
rect 9731 55637 9817 55693
rect 9873 55637 9959 55693
rect 10015 55637 10101 55693
rect 10157 55637 10243 55693
rect 10299 55637 10385 55693
rect 10441 55637 10527 55693
rect 10583 55637 10669 55693
rect 10725 55637 10811 55693
rect 10867 55637 10953 55693
rect 11009 55637 11095 55693
rect 11151 55637 11237 55693
rect 11293 55637 11379 55693
rect 11435 55637 11521 55693
rect 11577 55637 11663 55693
rect 11719 55637 11805 55693
rect 11861 55637 11947 55693
rect 12003 55637 12089 55693
rect 12145 55637 12231 55693
rect 12287 55637 12373 55693
rect 12429 55637 12515 55693
rect 12571 55637 12657 55693
rect 12713 55637 12799 55693
rect 12855 55637 12941 55693
rect 12997 55637 13083 55693
rect 13139 55637 13225 55693
rect 13281 55637 13367 55693
rect 13423 55637 13509 55693
rect 13565 55637 13651 55693
rect 13707 55637 13793 55693
rect 13849 55637 13935 55693
rect 13991 55637 14077 55693
rect 14133 55637 14219 55693
rect 14275 55637 14361 55693
rect 14417 55637 14503 55693
rect 14559 55637 14645 55693
rect 14701 55637 14787 55693
rect 14843 55637 14853 55693
rect 151 55627 14853 55637
rect 151 55363 14853 55373
rect 151 55307 161 55363
rect 217 55307 303 55363
rect 359 55307 445 55363
rect 501 55307 587 55363
rect 643 55307 729 55363
rect 785 55307 871 55363
rect 927 55307 1013 55363
rect 1069 55307 1155 55363
rect 1211 55307 1297 55363
rect 1353 55307 1439 55363
rect 1495 55307 1581 55363
rect 1637 55307 1723 55363
rect 1779 55307 1865 55363
rect 1921 55307 2007 55363
rect 2063 55307 2149 55363
rect 2205 55307 2291 55363
rect 2347 55307 2433 55363
rect 2489 55307 2575 55363
rect 2631 55307 2717 55363
rect 2773 55307 2859 55363
rect 2915 55307 3001 55363
rect 3057 55307 3143 55363
rect 3199 55307 3285 55363
rect 3341 55307 3427 55363
rect 3483 55307 3569 55363
rect 3625 55307 3711 55363
rect 3767 55307 3853 55363
rect 3909 55307 3995 55363
rect 4051 55307 4137 55363
rect 4193 55307 4279 55363
rect 4335 55307 4421 55363
rect 4477 55307 4563 55363
rect 4619 55307 4705 55363
rect 4761 55307 4847 55363
rect 4903 55307 4989 55363
rect 5045 55307 5131 55363
rect 5187 55307 5273 55363
rect 5329 55307 5415 55363
rect 5471 55307 5557 55363
rect 5613 55307 5699 55363
rect 5755 55307 5841 55363
rect 5897 55307 5983 55363
rect 6039 55307 6125 55363
rect 6181 55307 6267 55363
rect 6323 55307 6409 55363
rect 6465 55307 6551 55363
rect 6607 55307 6693 55363
rect 6749 55307 6835 55363
rect 6891 55307 6977 55363
rect 7033 55307 7119 55363
rect 7175 55307 7261 55363
rect 7317 55307 7403 55363
rect 7459 55307 7545 55363
rect 7601 55307 7687 55363
rect 7743 55307 7829 55363
rect 7885 55307 7971 55363
rect 8027 55307 8113 55363
rect 8169 55307 8255 55363
rect 8311 55307 8397 55363
rect 8453 55307 8539 55363
rect 8595 55307 8681 55363
rect 8737 55307 8823 55363
rect 8879 55307 8965 55363
rect 9021 55307 9107 55363
rect 9163 55307 9249 55363
rect 9305 55307 9391 55363
rect 9447 55307 9533 55363
rect 9589 55307 9675 55363
rect 9731 55307 9817 55363
rect 9873 55307 9959 55363
rect 10015 55307 10101 55363
rect 10157 55307 10243 55363
rect 10299 55307 10385 55363
rect 10441 55307 10527 55363
rect 10583 55307 10669 55363
rect 10725 55307 10811 55363
rect 10867 55307 10953 55363
rect 11009 55307 11095 55363
rect 11151 55307 11237 55363
rect 11293 55307 11379 55363
rect 11435 55307 11521 55363
rect 11577 55307 11663 55363
rect 11719 55307 11805 55363
rect 11861 55307 11947 55363
rect 12003 55307 12089 55363
rect 12145 55307 12231 55363
rect 12287 55307 12373 55363
rect 12429 55307 12515 55363
rect 12571 55307 12657 55363
rect 12713 55307 12799 55363
rect 12855 55307 12941 55363
rect 12997 55307 13083 55363
rect 13139 55307 13225 55363
rect 13281 55307 13367 55363
rect 13423 55307 13509 55363
rect 13565 55307 13651 55363
rect 13707 55307 13793 55363
rect 13849 55307 13935 55363
rect 13991 55307 14077 55363
rect 14133 55307 14219 55363
rect 14275 55307 14361 55363
rect 14417 55307 14503 55363
rect 14559 55307 14645 55363
rect 14701 55307 14787 55363
rect 14843 55307 14853 55363
rect 151 55221 14853 55307
rect 151 55165 161 55221
rect 217 55165 303 55221
rect 359 55165 445 55221
rect 501 55165 587 55221
rect 643 55165 729 55221
rect 785 55165 871 55221
rect 927 55165 1013 55221
rect 1069 55165 1155 55221
rect 1211 55165 1297 55221
rect 1353 55165 1439 55221
rect 1495 55165 1581 55221
rect 1637 55165 1723 55221
rect 1779 55165 1865 55221
rect 1921 55165 2007 55221
rect 2063 55165 2149 55221
rect 2205 55165 2291 55221
rect 2347 55165 2433 55221
rect 2489 55165 2575 55221
rect 2631 55165 2717 55221
rect 2773 55165 2859 55221
rect 2915 55165 3001 55221
rect 3057 55165 3143 55221
rect 3199 55165 3285 55221
rect 3341 55165 3427 55221
rect 3483 55165 3569 55221
rect 3625 55165 3711 55221
rect 3767 55165 3853 55221
rect 3909 55165 3995 55221
rect 4051 55165 4137 55221
rect 4193 55165 4279 55221
rect 4335 55165 4421 55221
rect 4477 55165 4563 55221
rect 4619 55165 4705 55221
rect 4761 55165 4847 55221
rect 4903 55165 4989 55221
rect 5045 55165 5131 55221
rect 5187 55165 5273 55221
rect 5329 55165 5415 55221
rect 5471 55165 5557 55221
rect 5613 55165 5699 55221
rect 5755 55165 5841 55221
rect 5897 55165 5983 55221
rect 6039 55165 6125 55221
rect 6181 55165 6267 55221
rect 6323 55165 6409 55221
rect 6465 55165 6551 55221
rect 6607 55165 6693 55221
rect 6749 55165 6835 55221
rect 6891 55165 6977 55221
rect 7033 55165 7119 55221
rect 7175 55165 7261 55221
rect 7317 55165 7403 55221
rect 7459 55165 7545 55221
rect 7601 55165 7687 55221
rect 7743 55165 7829 55221
rect 7885 55165 7971 55221
rect 8027 55165 8113 55221
rect 8169 55165 8255 55221
rect 8311 55165 8397 55221
rect 8453 55165 8539 55221
rect 8595 55165 8681 55221
rect 8737 55165 8823 55221
rect 8879 55165 8965 55221
rect 9021 55165 9107 55221
rect 9163 55165 9249 55221
rect 9305 55165 9391 55221
rect 9447 55165 9533 55221
rect 9589 55165 9675 55221
rect 9731 55165 9817 55221
rect 9873 55165 9959 55221
rect 10015 55165 10101 55221
rect 10157 55165 10243 55221
rect 10299 55165 10385 55221
rect 10441 55165 10527 55221
rect 10583 55165 10669 55221
rect 10725 55165 10811 55221
rect 10867 55165 10953 55221
rect 11009 55165 11095 55221
rect 11151 55165 11237 55221
rect 11293 55165 11379 55221
rect 11435 55165 11521 55221
rect 11577 55165 11663 55221
rect 11719 55165 11805 55221
rect 11861 55165 11947 55221
rect 12003 55165 12089 55221
rect 12145 55165 12231 55221
rect 12287 55165 12373 55221
rect 12429 55165 12515 55221
rect 12571 55165 12657 55221
rect 12713 55165 12799 55221
rect 12855 55165 12941 55221
rect 12997 55165 13083 55221
rect 13139 55165 13225 55221
rect 13281 55165 13367 55221
rect 13423 55165 13509 55221
rect 13565 55165 13651 55221
rect 13707 55165 13793 55221
rect 13849 55165 13935 55221
rect 13991 55165 14077 55221
rect 14133 55165 14219 55221
rect 14275 55165 14361 55221
rect 14417 55165 14503 55221
rect 14559 55165 14645 55221
rect 14701 55165 14787 55221
rect 14843 55165 14853 55221
rect 151 55079 14853 55165
rect 151 55023 161 55079
rect 217 55023 303 55079
rect 359 55023 445 55079
rect 501 55023 587 55079
rect 643 55023 729 55079
rect 785 55023 871 55079
rect 927 55023 1013 55079
rect 1069 55023 1155 55079
rect 1211 55023 1297 55079
rect 1353 55023 1439 55079
rect 1495 55023 1581 55079
rect 1637 55023 1723 55079
rect 1779 55023 1865 55079
rect 1921 55023 2007 55079
rect 2063 55023 2149 55079
rect 2205 55023 2291 55079
rect 2347 55023 2433 55079
rect 2489 55023 2575 55079
rect 2631 55023 2717 55079
rect 2773 55023 2859 55079
rect 2915 55023 3001 55079
rect 3057 55023 3143 55079
rect 3199 55023 3285 55079
rect 3341 55023 3427 55079
rect 3483 55023 3569 55079
rect 3625 55023 3711 55079
rect 3767 55023 3853 55079
rect 3909 55023 3995 55079
rect 4051 55023 4137 55079
rect 4193 55023 4279 55079
rect 4335 55023 4421 55079
rect 4477 55023 4563 55079
rect 4619 55023 4705 55079
rect 4761 55023 4847 55079
rect 4903 55023 4989 55079
rect 5045 55023 5131 55079
rect 5187 55023 5273 55079
rect 5329 55023 5415 55079
rect 5471 55023 5557 55079
rect 5613 55023 5699 55079
rect 5755 55023 5841 55079
rect 5897 55023 5983 55079
rect 6039 55023 6125 55079
rect 6181 55023 6267 55079
rect 6323 55023 6409 55079
rect 6465 55023 6551 55079
rect 6607 55023 6693 55079
rect 6749 55023 6835 55079
rect 6891 55023 6977 55079
rect 7033 55023 7119 55079
rect 7175 55023 7261 55079
rect 7317 55023 7403 55079
rect 7459 55023 7545 55079
rect 7601 55023 7687 55079
rect 7743 55023 7829 55079
rect 7885 55023 7971 55079
rect 8027 55023 8113 55079
rect 8169 55023 8255 55079
rect 8311 55023 8397 55079
rect 8453 55023 8539 55079
rect 8595 55023 8681 55079
rect 8737 55023 8823 55079
rect 8879 55023 8965 55079
rect 9021 55023 9107 55079
rect 9163 55023 9249 55079
rect 9305 55023 9391 55079
rect 9447 55023 9533 55079
rect 9589 55023 9675 55079
rect 9731 55023 9817 55079
rect 9873 55023 9959 55079
rect 10015 55023 10101 55079
rect 10157 55023 10243 55079
rect 10299 55023 10385 55079
rect 10441 55023 10527 55079
rect 10583 55023 10669 55079
rect 10725 55023 10811 55079
rect 10867 55023 10953 55079
rect 11009 55023 11095 55079
rect 11151 55023 11237 55079
rect 11293 55023 11379 55079
rect 11435 55023 11521 55079
rect 11577 55023 11663 55079
rect 11719 55023 11805 55079
rect 11861 55023 11947 55079
rect 12003 55023 12089 55079
rect 12145 55023 12231 55079
rect 12287 55023 12373 55079
rect 12429 55023 12515 55079
rect 12571 55023 12657 55079
rect 12713 55023 12799 55079
rect 12855 55023 12941 55079
rect 12997 55023 13083 55079
rect 13139 55023 13225 55079
rect 13281 55023 13367 55079
rect 13423 55023 13509 55079
rect 13565 55023 13651 55079
rect 13707 55023 13793 55079
rect 13849 55023 13935 55079
rect 13991 55023 14077 55079
rect 14133 55023 14219 55079
rect 14275 55023 14361 55079
rect 14417 55023 14503 55079
rect 14559 55023 14645 55079
rect 14701 55023 14787 55079
rect 14843 55023 14853 55079
rect 151 54937 14853 55023
rect 151 54881 161 54937
rect 217 54881 303 54937
rect 359 54881 445 54937
rect 501 54881 587 54937
rect 643 54881 729 54937
rect 785 54881 871 54937
rect 927 54881 1013 54937
rect 1069 54881 1155 54937
rect 1211 54881 1297 54937
rect 1353 54881 1439 54937
rect 1495 54881 1581 54937
rect 1637 54881 1723 54937
rect 1779 54881 1865 54937
rect 1921 54881 2007 54937
rect 2063 54881 2149 54937
rect 2205 54881 2291 54937
rect 2347 54881 2433 54937
rect 2489 54881 2575 54937
rect 2631 54881 2717 54937
rect 2773 54881 2859 54937
rect 2915 54881 3001 54937
rect 3057 54881 3143 54937
rect 3199 54881 3285 54937
rect 3341 54881 3427 54937
rect 3483 54881 3569 54937
rect 3625 54881 3711 54937
rect 3767 54881 3853 54937
rect 3909 54881 3995 54937
rect 4051 54881 4137 54937
rect 4193 54881 4279 54937
rect 4335 54881 4421 54937
rect 4477 54881 4563 54937
rect 4619 54881 4705 54937
rect 4761 54881 4847 54937
rect 4903 54881 4989 54937
rect 5045 54881 5131 54937
rect 5187 54881 5273 54937
rect 5329 54881 5415 54937
rect 5471 54881 5557 54937
rect 5613 54881 5699 54937
rect 5755 54881 5841 54937
rect 5897 54881 5983 54937
rect 6039 54881 6125 54937
rect 6181 54881 6267 54937
rect 6323 54881 6409 54937
rect 6465 54881 6551 54937
rect 6607 54881 6693 54937
rect 6749 54881 6835 54937
rect 6891 54881 6977 54937
rect 7033 54881 7119 54937
rect 7175 54881 7261 54937
rect 7317 54881 7403 54937
rect 7459 54881 7545 54937
rect 7601 54881 7687 54937
rect 7743 54881 7829 54937
rect 7885 54881 7971 54937
rect 8027 54881 8113 54937
rect 8169 54881 8255 54937
rect 8311 54881 8397 54937
rect 8453 54881 8539 54937
rect 8595 54881 8681 54937
rect 8737 54881 8823 54937
rect 8879 54881 8965 54937
rect 9021 54881 9107 54937
rect 9163 54881 9249 54937
rect 9305 54881 9391 54937
rect 9447 54881 9533 54937
rect 9589 54881 9675 54937
rect 9731 54881 9817 54937
rect 9873 54881 9959 54937
rect 10015 54881 10101 54937
rect 10157 54881 10243 54937
rect 10299 54881 10385 54937
rect 10441 54881 10527 54937
rect 10583 54881 10669 54937
rect 10725 54881 10811 54937
rect 10867 54881 10953 54937
rect 11009 54881 11095 54937
rect 11151 54881 11237 54937
rect 11293 54881 11379 54937
rect 11435 54881 11521 54937
rect 11577 54881 11663 54937
rect 11719 54881 11805 54937
rect 11861 54881 11947 54937
rect 12003 54881 12089 54937
rect 12145 54881 12231 54937
rect 12287 54881 12373 54937
rect 12429 54881 12515 54937
rect 12571 54881 12657 54937
rect 12713 54881 12799 54937
rect 12855 54881 12941 54937
rect 12997 54881 13083 54937
rect 13139 54881 13225 54937
rect 13281 54881 13367 54937
rect 13423 54881 13509 54937
rect 13565 54881 13651 54937
rect 13707 54881 13793 54937
rect 13849 54881 13935 54937
rect 13991 54881 14077 54937
rect 14133 54881 14219 54937
rect 14275 54881 14361 54937
rect 14417 54881 14503 54937
rect 14559 54881 14645 54937
rect 14701 54881 14787 54937
rect 14843 54881 14853 54937
rect 151 54795 14853 54881
rect 151 54739 161 54795
rect 217 54739 303 54795
rect 359 54739 445 54795
rect 501 54739 587 54795
rect 643 54739 729 54795
rect 785 54739 871 54795
rect 927 54739 1013 54795
rect 1069 54739 1155 54795
rect 1211 54739 1297 54795
rect 1353 54739 1439 54795
rect 1495 54739 1581 54795
rect 1637 54739 1723 54795
rect 1779 54739 1865 54795
rect 1921 54739 2007 54795
rect 2063 54739 2149 54795
rect 2205 54739 2291 54795
rect 2347 54739 2433 54795
rect 2489 54739 2575 54795
rect 2631 54739 2717 54795
rect 2773 54739 2859 54795
rect 2915 54739 3001 54795
rect 3057 54739 3143 54795
rect 3199 54739 3285 54795
rect 3341 54739 3427 54795
rect 3483 54739 3569 54795
rect 3625 54739 3711 54795
rect 3767 54739 3853 54795
rect 3909 54739 3995 54795
rect 4051 54739 4137 54795
rect 4193 54739 4279 54795
rect 4335 54739 4421 54795
rect 4477 54739 4563 54795
rect 4619 54739 4705 54795
rect 4761 54739 4847 54795
rect 4903 54739 4989 54795
rect 5045 54739 5131 54795
rect 5187 54739 5273 54795
rect 5329 54739 5415 54795
rect 5471 54739 5557 54795
rect 5613 54739 5699 54795
rect 5755 54739 5841 54795
rect 5897 54739 5983 54795
rect 6039 54739 6125 54795
rect 6181 54739 6267 54795
rect 6323 54739 6409 54795
rect 6465 54739 6551 54795
rect 6607 54739 6693 54795
rect 6749 54739 6835 54795
rect 6891 54739 6977 54795
rect 7033 54739 7119 54795
rect 7175 54739 7261 54795
rect 7317 54739 7403 54795
rect 7459 54739 7545 54795
rect 7601 54739 7687 54795
rect 7743 54739 7829 54795
rect 7885 54739 7971 54795
rect 8027 54739 8113 54795
rect 8169 54739 8255 54795
rect 8311 54739 8397 54795
rect 8453 54739 8539 54795
rect 8595 54739 8681 54795
rect 8737 54739 8823 54795
rect 8879 54739 8965 54795
rect 9021 54739 9107 54795
rect 9163 54739 9249 54795
rect 9305 54739 9391 54795
rect 9447 54739 9533 54795
rect 9589 54739 9675 54795
rect 9731 54739 9817 54795
rect 9873 54739 9959 54795
rect 10015 54739 10101 54795
rect 10157 54739 10243 54795
rect 10299 54739 10385 54795
rect 10441 54739 10527 54795
rect 10583 54739 10669 54795
rect 10725 54739 10811 54795
rect 10867 54739 10953 54795
rect 11009 54739 11095 54795
rect 11151 54739 11237 54795
rect 11293 54739 11379 54795
rect 11435 54739 11521 54795
rect 11577 54739 11663 54795
rect 11719 54739 11805 54795
rect 11861 54739 11947 54795
rect 12003 54739 12089 54795
rect 12145 54739 12231 54795
rect 12287 54739 12373 54795
rect 12429 54739 12515 54795
rect 12571 54739 12657 54795
rect 12713 54739 12799 54795
rect 12855 54739 12941 54795
rect 12997 54739 13083 54795
rect 13139 54739 13225 54795
rect 13281 54739 13367 54795
rect 13423 54739 13509 54795
rect 13565 54739 13651 54795
rect 13707 54739 13793 54795
rect 13849 54739 13935 54795
rect 13991 54739 14077 54795
rect 14133 54739 14219 54795
rect 14275 54739 14361 54795
rect 14417 54739 14503 54795
rect 14559 54739 14645 54795
rect 14701 54739 14787 54795
rect 14843 54739 14853 54795
rect 151 54653 14853 54739
rect 151 54597 161 54653
rect 217 54597 303 54653
rect 359 54597 445 54653
rect 501 54597 587 54653
rect 643 54597 729 54653
rect 785 54597 871 54653
rect 927 54597 1013 54653
rect 1069 54597 1155 54653
rect 1211 54597 1297 54653
rect 1353 54597 1439 54653
rect 1495 54597 1581 54653
rect 1637 54597 1723 54653
rect 1779 54597 1865 54653
rect 1921 54597 2007 54653
rect 2063 54597 2149 54653
rect 2205 54597 2291 54653
rect 2347 54597 2433 54653
rect 2489 54597 2575 54653
rect 2631 54597 2717 54653
rect 2773 54597 2859 54653
rect 2915 54597 3001 54653
rect 3057 54597 3143 54653
rect 3199 54597 3285 54653
rect 3341 54597 3427 54653
rect 3483 54597 3569 54653
rect 3625 54597 3711 54653
rect 3767 54597 3853 54653
rect 3909 54597 3995 54653
rect 4051 54597 4137 54653
rect 4193 54597 4279 54653
rect 4335 54597 4421 54653
rect 4477 54597 4563 54653
rect 4619 54597 4705 54653
rect 4761 54597 4847 54653
rect 4903 54597 4989 54653
rect 5045 54597 5131 54653
rect 5187 54597 5273 54653
rect 5329 54597 5415 54653
rect 5471 54597 5557 54653
rect 5613 54597 5699 54653
rect 5755 54597 5841 54653
rect 5897 54597 5983 54653
rect 6039 54597 6125 54653
rect 6181 54597 6267 54653
rect 6323 54597 6409 54653
rect 6465 54597 6551 54653
rect 6607 54597 6693 54653
rect 6749 54597 6835 54653
rect 6891 54597 6977 54653
rect 7033 54597 7119 54653
rect 7175 54597 7261 54653
rect 7317 54597 7403 54653
rect 7459 54597 7545 54653
rect 7601 54597 7687 54653
rect 7743 54597 7829 54653
rect 7885 54597 7971 54653
rect 8027 54597 8113 54653
rect 8169 54597 8255 54653
rect 8311 54597 8397 54653
rect 8453 54597 8539 54653
rect 8595 54597 8681 54653
rect 8737 54597 8823 54653
rect 8879 54597 8965 54653
rect 9021 54597 9107 54653
rect 9163 54597 9249 54653
rect 9305 54597 9391 54653
rect 9447 54597 9533 54653
rect 9589 54597 9675 54653
rect 9731 54597 9817 54653
rect 9873 54597 9959 54653
rect 10015 54597 10101 54653
rect 10157 54597 10243 54653
rect 10299 54597 10385 54653
rect 10441 54597 10527 54653
rect 10583 54597 10669 54653
rect 10725 54597 10811 54653
rect 10867 54597 10953 54653
rect 11009 54597 11095 54653
rect 11151 54597 11237 54653
rect 11293 54597 11379 54653
rect 11435 54597 11521 54653
rect 11577 54597 11663 54653
rect 11719 54597 11805 54653
rect 11861 54597 11947 54653
rect 12003 54597 12089 54653
rect 12145 54597 12231 54653
rect 12287 54597 12373 54653
rect 12429 54597 12515 54653
rect 12571 54597 12657 54653
rect 12713 54597 12799 54653
rect 12855 54597 12941 54653
rect 12997 54597 13083 54653
rect 13139 54597 13225 54653
rect 13281 54597 13367 54653
rect 13423 54597 13509 54653
rect 13565 54597 13651 54653
rect 13707 54597 13793 54653
rect 13849 54597 13935 54653
rect 13991 54597 14077 54653
rect 14133 54597 14219 54653
rect 14275 54597 14361 54653
rect 14417 54597 14503 54653
rect 14559 54597 14645 54653
rect 14701 54597 14787 54653
rect 14843 54597 14853 54653
rect 151 54511 14853 54597
rect 151 54455 161 54511
rect 217 54455 303 54511
rect 359 54455 445 54511
rect 501 54455 587 54511
rect 643 54455 729 54511
rect 785 54455 871 54511
rect 927 54455 1013 54511
rect 1069 54455 1155 54511
rect 1211 54455 1297 54511
rect 1353 54455 1439 54511
rect 1495 54455 1581 54511
rect 1637 54455 1723 54511
rect 1779 54455 1865 54511
rect 1921 54455 2007 54511
rect 2063 54455 2149 54511
rect 2205 54455 2291 54511
rect 2347 54455 2433 54511
rect 2489 54455 2575 54511
rect 2631 54455 2717 54511
rect 2773 54455 2859 54511
rect 2915 54455 3001 54511
rect 3057 54455 3143 54511
rect 3199 54455 3285 54511
rect 3341 54455 3427 54511
rect 3483 54455 3569 54511
rect 3625 54455 3711 54511
rect 3767 54455 3853 54511
rect 3909 54455 3995 54511
rect 4051 54455 4137 54511
rect 4193 54455 4279 54511
rect 4335 54455 4421 54511
rect 4477 54455 4563 54511
rect 4619 54455 4705 54511
rect 4761 54455 4847 54511
rect 4903 54455 4989 54511
rect 5045 54455 5131 54511
rect 5187 54455 5273 54511
rect 5329 54455 5415 54511
rect 5471 54455 5557 54511
rect 5613 54455 5699 54511
rect 5755 54455 5841 54511
rect 5897 54455 5983 54511
rect 6039 54455 6125 54511
rect 6181 54455 6267 54511
rect 6323 54455 6409 54511
rect 6465 54455 6551 54511
rect 6607 54455 6693 54511
rect 6749 54455 6835 54511
rect 6891 54455 6977 54511
rect 7033 54455 7119 54511
rect 7175 54455 7261 54511
rect 7317 54455 7403 54511
rect 7459 54455 7545 54511
rect 7601 54455 7687 54511
rect 7743 54455 7829 54511
rect 7885 54455 7971 54511
rect 8027 54455 8113 54511
rect 8169 54455 8255 54511
rect 8311 54455 8397 54511
rect 8453 54455 8539 54511
rect 8595 54455 8681 54511
rect 8737 54455 8823 54511
rect 8879 54455 8965 54511
rect 9021 54455 9107 54511
rect 9163 54455 9249 54511
rect 9305 54455 9391 54511
rect 9447 54455 9533 54511
rect 9589 54455 9675 54511
rect 9731 54455 9817 54511
rect 9873 54455 9959 54511
rect 10015 54455 10101 54511
rect 10157 54455 10243 54511
rect 10299 54455 10385 54511
rect 10441 54455 10527 54511
rect 10583 54455 10669 54511
rect 10725 54455 10811 54511
rect 10867 54455 10953 54511
rect 11009 54455 11095 54511
rect 11151 54455 11237 54511
rect 11293 54455 11379 54511
rect 11435 54455 11521 54511
rect 11577 54455 11663 54511
rect 11719 54455 11805 54511
rect 11861 54455 11947 54511
rect 12003 54455 12089 54511
rect 12145 54455 12231 54511
rect 12287 54455 12373 54511
rect 12429 54455 12515 54511
rect 12571 54455 12657 54511
rect 12713 54455 12799 54511
rect 12855 54455 12941 54511
rect 12997 54455 13083 54511
rect 13139 54455 13225 54511
rect 13281 54455 13367 54511
rect 13423 54455 13509 54511
rect 13565 54455 13651 54511
rect 13707 54455 13793 54511
rect 13849 54455 13935 54511
rect 13991 54455 14077 54511
rect 14133 54455 14219 54511
rect 14275 54455 14361 54511
rect 14417 54455 14503 54511
rect 14559 54455 14645 54511
rect 14701 54455 14787 54511
rect 14843 54455 14853 54511
rect 151 54369 14853 54455
rect 151 54313 161 54369
rect 217 54313 303 54369
rect 359 54313 445 54369
rect 501 54313 587 54369
rect 643 54313 729 54369
rect 785 54313 871 54369
rect 927 54313 1013 54369
rect 1069 54313 1155 54369
rect 1211 54313 1297 54369
rect 1353 54313 1439 54369
rect 1495 54313 1581 54369
rect 1637 54313 1723 54369
rect 1779 54313 1865 54369
rect 1921 54313 2007 54369
rect 2063 54313 2149 54369
rect 2205 54313 2291 54369
rect 2347 54313 2433 54369
rect 2489 54313 2575 54369
rect 2631 54313 2717 54369
rect 2773 54313 2859 54369
rect 2915 54313 3001 54369
rect 3057 54313 3143 54369
rect 3199 54313 3285 54369
rect 3341 54313 3427 54369
rect 3483 54313 3569 54369
rect 3625 54313 3711 54369
rect 3767 54313 3853 54369
rect 3909 54313 3995 54369
rect 4051 54313 4137 54369
rect 4193 54313 4279 54369
rect 4335 54313 4421 54369
rect 4477 54313 4563 54369
rect 4619 54313 4705 54369
rect 4761 54313 4847 54369
rect 4903 54313 4989 54369
rect 5045 54313 5131 54369
rect 5187 54313 5273 54369
rect 5329 54313 5415 54369
rect 5471 54313 5557 54369
rect 5613 54313 5699 54369
rect 5755 54313 5841 54369
rect 5897 54313 5983 54369
rect 6039 54313 6125 54369
rect 6181 54313 6267 54369
rect 6323 54313 6409 54369
rect 6465 54313 6551 54369
rect 6607 54313 6693 54369
rect 6749 54313 6835 54369
rect 6891 54313 6977 54369
rect 7033 54313 7119 54369
rect 7175 54313 7261 54369
rect 7317 54313 7403 54369
rect 7459 54313 7545 54369
rect 7601 54313 7687 54369
rect 7743 54313 7829 54369
rect 7885 54313 7971 54369
rect 8027 54313 8113 54369
rect 8169 54313 8255 54369
rect 8311 54313 8397 54369
rect 8453 54313 8539 54369
rect 8595 54313 8681 54369
rect 8737 54313 8823 54369
rect 8879 54313 8965 54369
rect 9021 54313 9107 54369
rect 9163 54313 9249 54369
rect 9305 54313 9391 54369
rect 9447 54313 9533 54369
rect 9589 54313 9675 54369
rect 9731 54313 9817 54369
rect 9873 54313 9959 54369
rect 10015 54313 10101 54369
rect 10157 54313 10243 54369
rect 10299 54313 10385 54369
rect 10441 54313 10527 54369
rect 10583 54313 10669 54369
rect 10725 54313 10811 54369
rect 10867 54313 10953 54369
rect 11009 54313 11095 54369
rect 11151 54313 11237 54369
rect 11293 54313 11379 54369
rect 11435 54313 11521 54369
rect 11577 54313 11663 54369
rect 11719 54313 11805 54369
rect 11861 54313 11947 54369
rect 12003 54313 12089 54369
rect 12145 54313 12231 54369
rect 12287 54313 12373 54369
rect 12429 54313 12515 54369
rect 12571 54313 12657 54369
rect 12713 54313 12799 54369
rect 12855 54313 12941 54369
rect 12997 54313 13083 54369
rect 13139 54313 13225 54369
rect 13281 54313 13367 54369
rect 13423 54313 13509 54369
rect 13565 54313 13651 54369
rect 13707 54313 13793 54369
rect 13849 54313 13935 54369
rect 13991 54313 14077 54369
rect 14133 54313 14219 54369
rect 14275 54313 14361 54369
rect 14417 54313 14503 54369
rect 14559 54313 14645 54369
rect 14701 54313 14787 54369
rect 14843 54313 14853 54369
rect 151 54227 14853 54313
rect 151 54171 161 54227
rect 217 54171 303 54227
rect 359 54171 445 54227
rect 501 54171 587 54227
rect 643 54171 729 54227
rect 785 54171 871 54227
rect 927 54171 1013 54227
rect 1069 54171 1155 54227
rect 1211 54171 1297 54227
rect 1353 54171 1439 54227
rect 1495 54171 1581 54227
rect 1637 54171 1723 54227
rect 1779 54171 1865 54227
rect 1921 54171 2007 54227
rect 2063 54171 2149 54227
rect 2205 54171 2291 54227
rect 2347 54171 2433 54227
rect 2489 54171 2575 54227
rect 2631 54171 2717 54227
rect 2773 54171 2859 54227
rect 2915 54171 3001 54227
rect 3057 54171 3143 54227
rect 3199 54171 3285 54227
rect 3341 54171 3427 54227
rect 3483 54171 3569 54227
rect 3625 54171 3711 54227
rect 3767 54171 3853 54227
rect 3909 54171 3995 54227
rect 4051 54171 4137 54227
rect 4193 54171 4279 54227
rect 4335 54171 4421 54227
rect 4477 54171 4563 54227
rect 4619 54171 4705 54227
rect 4761 54171 4847 54227
rect 4903 54171 4989 54227
rect 5045 54171 5131 54227
rect 5187 54171 5273 54227
rect 5329 54171 5415 54227
rect 5471 54171 5557 54227
rect 5613 54171 5699 54227
rect 5755 54171 5841 54227
rect 5897 54171 5983 54227
rect 6039 54171 6125 54227
rect 6181 54171 6267 54227
rect 6323 54171 6409 54227
rect 6465 54171 6551 54227
rect 6607 54171 6693 54227
rect 6749 54171 6835 54227
rect 6891 54171 6977 54227
rect 7033 54171 7119 54227
rect 7175 54171 7261 54227
rect 7317 54171 7403 54227
rect 7459 54171 7545 54227
rect 7601 54171 7687 54227
rect 7743 54171 7829 54227
rect 7885 54171 7971 54227
rect 8027 54171 8113 54227
rect 8169 54171 8255 54227
rect 8311 54171 8397 54227
rect 8453 54171 8539 54227
rect 8595 54171 8681 54227
rect 8737 54171 8823 54227
rect 8879 54171 8965 54227
rect 9021 54171 9107 54227
rect 9163 54171 9249 54227
rect 9305 54171 9391 54227
rect 9447 54171 9533 54227
rect 9589 54171 9675 54227
rect 9731 54171 9817 54227
rect 9873 54171 9959 54227
rect 10015 54171 10101 54227
rect 10157 54171 10243 54227
rect 10299 54171 10385 54227
rect 10441 54171 10527 54227
rect 10583 54171 10669 54227
rect 10725 54171 10811 54227
rect 10867 54171 10953 54227
rect 11009 54171 11095 54227
rect 11151 54171 11237 54227
rect 11293 54171 11379 54227
rect 11435 54171 11521 54227
rect 11577 54171 11663 54227
rect 11719 54171 11805 54227
rect 11861 54171 11947 54227
rect 12003 54171 12089 54227
rect 12145 54171 12231 54227
rect 12287 54171 12373 54227
rect 12429 54171 12515 54227
rect 12571 54171 12657 54227
rect 12713 54171 12799 54227
rect 12855 54171 12941 54227
rect 12997 54171 13083 54227
rect 13139 54171 13225 54227
rect 13281 54171 13367 54227
rect 13423 54171 13509 54227
rect 13565 54171 13651 54227
rect 13707 54171 13793 54227
rect 13849 54171 13935 54227
rect 13991 54171 14077 54227
rect 14133 54171 14219 54227
rect 14275 54171 14361 54227
rect 14417 54171 14503 54227
rect 14559 54171 14645 54227
rect 14701 54171 14787 54227
rect 14843 54171 14853 54227
rect 151 54085 14853 54171
rect 151 54029 161 54085
rect 217 54029 303 54085
rect 359 54029 445 54085
rect 501 54029 587 54085
rect 643 54029 729 54085
rect 785 54029 871 54085
rect 927 54029 1013 54085
rect 1069 54029 1155 54085
rect 1211 54029 1297 54085
rect 1353 54029 1439 54085
rect 1495 54029 1581 54085
rect 1637 54029 1723 54085
rect 1779 54029 1865 54085
rect 1921 54029 2007 54085
rect 2063 54029 2149 54085
rect 2205 54029 2291 54085
rect 2347 54029 2433 54085
rect 2489 54029 2575 54085
rect 2631 54029 2717 54085
rect 2773 54029 2859 54085
rect 2915 54029 3001 54085
rect 3057 54029 3143 54085
rect 3199 54029 3285 54085
rect 3341 54029 3427 54085
rect 3483 54029 3569 54085
rect 3625 54029 3711 54085
rect 3767 54029 3853 54085
rect 3909 54029 3995 54085
rect 4051 54029 4137 54085
rect 4193 54029 4279 54085
rect 4335 54029 4421 54085
rect 4477 54029 4563 54085
rect 4619 54029 4705 54085
rect 4761 54029 4847 54085
rect 4903 54029 4989 54085
rect 5045 54029 5131 54085
rect 5187 54029 5273 54085
rect 5329 54029 5415 54085
rect 5471 54029 5557 54085
rect 5613 54029 5699 54085
rect 5755 54029 5841 54085
rect 5897 54029 5983 54085
rect 6039 54029 6125 54085
rect 6181 54029 6267 54085
rect 6323 54029 6409 54085
rect 6465 54029 6551 54085
rect 6607 54029 6693 54085
rect 6749 54029 6835 54085
rect 6891 54029 6977 54085
rect 7033 54029 7119 54085
rect 7175 54029 7261 54085
rect 7317 54029 7403 54085
rect 7459 54029 7545 54085
rect 7601 54029 7687 54085
rect 7743 54029 7829 54085
rect 7885 54029 7971 54085
rect 8027 54029 8113 54085
rect 8169 54029 8255 54085
rect 8311 54029 8397 54085
rect 8453 54029 8539 54085
rect 8595 54029 8681 54085
rect 8737 54029 8823 54085
rect 8879 54029 8965 54085
rect 9021 54029 9107 54085
rect 9163 54029 9249 54085
rect 9305 54029 9391 54085
rect 9447 54029 9533 54085
rect 9589 54029 9675 54085
rect 9731 54029 9817 54085
rect 9873 54029 9959 54085
rect 10015 54029 10101 54085
rect 10157 54029 10243 54085
rect 10299 54029 10385 54085
rect 10441 54029 10527 54085
rect 10583 54029 10669 54085
rect 10725 54029 10811 54085
rect 10867 54029 10953 54085
rect 11009 54029 11095 54085
rect 11151 54029 11237 54085
rect 11293 54029 11379 54085
rect 11435 54029 11521 54085
rect 11577 54029 11663 54085
rect 11719 54029 11805 54085
rect 11861 54029 11947 54085
rect 12003 54029 12089 54085
rect 12145 54029 12231 54085
rect 12287 54029 12373 54085
rect 12429 54029 12515 54085
rect 12571 54029 12657 54085
rect 12713 54029 12799 54085
rect 12855 54029 12941 54085
rect 12997 54029 13083 54085
rect 13139 54029 13225 54085
rect 13281 54029 13367 54085
rect 13423 54029 13509 54085
rect 13565 54029 13651 54085
rect 13707 54029 13793 54085
rect 13849 54029 13935 54085
rect 13991 54029 14077 54085
rect 14133 54029 14219 54085
rect 14275 54029 14361 54085
rect 14417 54029 14503 54085
rect 14559 54029 14645 54085
rect 14701 54029 14787 54085
rect 14843 54029 14853 54085
rect 151 54019 14853 54029
rect 151 53771 14853 53781
rect 151 53715 161 53771
rect 217 53715 303 53771
rect 359 53715 445 53771
rect 501 53715 587 53771
rect 643 53715 729 53771
rect 785 53715 871 53771
rect 927 53715 1013 53771
rect 1069 53715 1155 53771
rect 1211 53715 1297 53771
rect 1353 53715 1439 53771
rect 1495 53715 1581 53771
rect 1637 53715 1723 53771
rect 1779 53715 1865 53771
rect 1921 53715 2007 53771
rect 2063 53715 2149 53771
rect 2205 53715 2291 53771
rect 2347 53715 2433 53771
rect 2489 53715 2575 53771
rect 2631 53715 2717 53771
rect 2773 53715 2859 53771
rect 2915 53715 3001 53771
rect 3057 53715 3143 53771
rect 3199 53715 3285 53771
rect 3341 53715 3427 53771
rect 3483 53715 3569 53771
rect 3625 53715 3711 53771
rect 3767 53715 3853 53771
rect 3909 53715 3995 53771
rect 4051 53715 4137 53771
rect 4193 53715 4279 53771
rect 4335 53715 4421 53771
rect 4477 53715 4563 53771
rect 4619 53715 4705 53771
rect 4761 53715 4847 53771
rect 4903 53715 4989 53771
rect 5045 53715 5131 53771
rect 5187 53715 5273 53771
rect 5329 53715 5415 53771
rect 5471 53715 5557 53771
rect 5613 53715 5699 53771
rect 5755 53715 5841 53771
rect 5897 53715 5983 53771
rect 6039 53715 6125 53771
rect 6181 53715 6267 53771
rect 6323 53715 6409 53771
rect 6465 53715 6551 53771
rect 6607 53715 6693 53771
rect 6749 53715 6835 53771
rect 6891 53715 6977 53771
rect 7033 53715 7119 53771
rect 7175 53715 7261 53771
rect 7317 53715 7403 53771
rect 7459 53715 7545 53771
rect 7601 53715 7687 53771
rect 7743 53715 7829 53771
rect 7885 53715 7971 53771
rect 8027 53715 8113 53771
rect 8169 53715 8255 53771
rect 8311 53715 8397 53771
rect 8453 53715 8539 53771
rect 8595 53715 8681 53771
rect 8737 53715 8823 53771
rect 8879 53715 8965 53771
rect 9021 53715 9107 53771
rect 9163 53715 9249 53771
rect 9305 53715 9391 53771
rect 9447 53715 9533 53771
rect 9589 53715 9675 53771
rect 9731 53715 9817 53771
rect 9873 53715 9959 53771
rect 10015 53715 10101 53771
rect 10157 53715 10243 53771
rect 10299 53715 10385 53771
rect 10441 53715 10527 53771
rect 10583 53715 10669 53771
rect 10725 53715 10811 53771
rect 10867 53715 10953 53771
rect 11009 53715 11095 53771
rect 11151 53715 11237 53771
rect 11293 53715 11379 53771
rect 11435 53715 11521 53771
rect 11577 53715 11663 53771
rect 11719 53715 11805 53771
rect 11861 53715 11947 53771
rect 12003 53715 12089 53771
rect 12145 53715 12231 53771
rect 12287 53715 12373 53771
rect 12429 53715 12515 53771
rect 12571 53715 12657 53771
rect 12713 53715 12799 53771
rect 12855 53715 12941 53771
rect 12997 53715 13083 53771
rect 13139 53715 13225 53771
rect 13281 53715 13367 53771
rect 13423 53715 13509 53771
rect 13565 53715 13651 53771
rect 13707 53715 13793 53771
rect 13849 53715 13935 53771
rect 13991 53715 14077 53771
rect 14133 53715 14219 53771
rect 14275 53715 14361 53771
rect 14417 53715 14503 53771
rect 14559 53715 14645 53771
rect 14701 53715 14787 53771
rect 14843 53715 14853 53771
rect 151 53629 14853 53715
rect 151 53573 161 53629
rect 217 53573 303 53629
rect 359 53573 445 53629
rect 501 53573 587 53629
rect 643 53573 729 53629
rect 785 53573 871 53629
rect 927 53573 1013 53629
rect 1069 53573 1155 53629
rect 1211 53573 1297 53629
rect 1353 53573 1439 53629
rect 1495 53573 1581 53629
rect 1637 53573 1723 53629
rect 1779 53573 1865 53629
rect 1921 53573 2007 53629
rect 2063 53573 2149 53629
rect 2205 53573 2291 53629
rect 2347 53573 2433 53629
rect 2489 53573 2575 53629
rect 2631 53573 2717 53629
rect 2773 53573 2859 53629
rect 2915 53573 3001 53629
rect 3057 53573 3143 53629
rect 3199 53573 3285 53629
rect 3341 53573 3427 53629
rect 3483 53573 3569 53629
rect 3625 53573 3711 53629
rect 3767 53573 3853 53629
rect 3909 53573 3995 53629
rect 4051 53573 4137 53629
rect 4193 53573 4279 53629
rect 4335 53573 4421 53629
rect 4477 53573 4563 53629
rect 4619 53573 4705 53629
rect 4761 53573 4847 53629
rect 4903 53573 4989 53629
rect 5045 53573 5131 53629
rect 5187 53573 5273 53629
rect 5329 53573 5415 53629
rect 5471 53573 5557 53629
rect 5613 53573 5699 53629
rect 5755 53573 5841 53629
rect 5897 53573 5983 53629
rect 6039 53573 6125 53629
rect 6181 53573 6267 53629
rect 6323 53573 6409 53629
rect 6465 53573 6551 53629
rect 6607 53573 6693 53629
rect 6749 53573 6835 53629
rect 6891 53573 6977 53629
rect 7033 53573 7119 53629
rect 7175 53573 7261 53629
rect 7317 53573 7403 53629
rect 7459 53573 7545 53629
rect 7601 53573 7687 53629
rect 7743 53573 7829 53629
rect 7885 53573 7971 53629
rect 8027 53573 8113 53629
rect 8169 53573 8255 53629
rect 8311 53573 8397 53629
rect 8453 53573 8539 53629
rect 8595 53573 8681 53629
rect 8737 53573 8823 53629
rect 8879 53573 8965 53629
rect 9021 53573 9107 53629
rect 9163 53573 9249 53629
rect 9305 53573 9391 53629
rect 9447 53573 9533 53629
rect 9589 53573 9675 53629
rect 9731 53573 9817 53629
rect 9873 53573 9959 53629
rect 10015 53573 10101 53629
rect 10157 53573 10243 53629
rect 10299 53573 10385 53629
rect 10441 53573 10527 53629
rect 10583 53573 10669 53629
rect 10725 53573 10811 53629
rect 10867 53573 10953 53629
rect 11009 53573 11095 53629
rect 11151 53573 11237 53629
rect 11293 53573 11379 53629
rect 11435 53573 11521 53629
rect 11577 53573 11663 53629
rect 11719 53573 11805 53629
rect 11861 53573 11947 53629
rect 12003 53573 12089 53629
rect 12145 53573 12231 53629
rect 12287 53573 12373 53629
rect 12429 53573 12515 53629
rect 12571 53573 12657 53629
rect 12713 53573 12799 53629
rect 12855 53573 12941 53629
rect 12997 53573 13083 53629
rect 13139 53573 13225 53629
rect 13281 53573 13367 53629
rect 13423 53573 13509 53629
rect 13565 53573 13651 53629
rect 13707 53573 13793 53629
rect 13849 53573 13935 53629
rect 13991 53573 14077 53629
rect 14133 53573 14219 53629
rect 14275 53573 14361 53629
rect 14417 53573 14503 53629
rect 14559 53573 14645 53629
rect 14701 53573 14787 53629
rect 14843 53573 14853 53629
rect 151 53487 14853 53573
rect 151 53431 161 53487
rect 217 53431 303 53487
rect 359 53431 445 53487
rect 501 53431 587 53487
rect 643 53431 729 53487
rect 785 53431 871 53487
rect 927 53431 1013 53487
rect 1069 53431 1155 53487
rect 1211 53431 1297 53487
rect 1353 53431 1439 53487
rect 1495 53431 1581 53487
rect 1637 53431 1723 53487
rect 1779 53431 1865 53487
rect 1921 53431 2007 53487
rect 2063 53431 2149 53487
rect 2205 53431 2291 53487
rect 2347 53431 2433 53487
rect 2489 53431 2575 53487
rect 2631 53431 2717 53487
rect 2773 53431 2859 53487
rect 2915 53431 3001 53487
rect 3057 53431 3143 53487
rect 3199 53431 3285 53487
rect 3341 53431 3427 53487
rect 3483 53431 3569 53487
rect 3625 53431 3711 53487
rect 3767 53431 3853 53487
rect 3909 53431 3995 53487
rect 4051 53431 4137 53487
rect 4193 53431 4279 53487
rect 4335 53431 4421 53487
rect 4477 53431 4563 53487
rect 4619 53431 4705 53487
rect 4761 53431 4847 53487
rect 4903 53431 4989 53487
rect 5045 53431 5131 53487
rect 5187 53431 5273 53487
rect 5329 53431 5415 53487
rect 5471 53431 5557 53487
rect 5613 53431 5699 53487
rect 5755 53431 5841 53487
rect 5897 53431 5983 53487
rect 6039 53431 6125 53487
rect 6181 53431 6267 53487
rect 6323 53431 6409 53487
rect 6465 53431 6551 53487
rect 6607 53431 6693 53487
rect 6749 53431 6835 53487
rect 6891 53431 6977 53487
rect 7033 53431 7119 53487
rect 7175 53431 7261 53487
rect 7317 53431 7403 53487
rect 7459 53431 7545 53487
rect 7601 53431 7687 53487
rect 7743 53431 7829 53487
rect 7885 53431 7971 53487
rect 8027 53431 8113 53487
rect 8169 53431 8255 53487
rect 8311 53431 8397 53487
rect 8453 53431 8539 53487
rect 8595 53431 8681 53487
rect 8737 53431 8823 53487
rect 8879 53431 8965 53487
rect 9021 53431 9107 53487
rect 9163 53431 9249 53487
rect 9305 53431 9391 53487
rect 9447 53431 9533 53487
rect 9589 53431 9675 53487
rect 9731 53431 9817 53487
rect 9873 53431 9959 53487
rect 10015 53431 10101 53487
rect 10157 53431 10243 53487
rect 10299 53431 10385 53487
rect 10441 53431 10527 53487
rect 10583 53431 10669 53487
rect 10725 53431 10811 53487
rect 10867 53431 10953 53487
rect 11009 53431 11095 53487
rect 11151 53431 11237 53487
rect 11293 53431 11379 53487
rect 11435 53431 11521 53487
rect 11577 53431 11663 53487
rect 11719 53431 11805 53487
rect 11861 53431 11947 53487
rect 12003 53431 12089 53487
rect 12145 53431 12231 53487
rect 12287 53431 12373 53487
rect 12429 53431 12515 53487
rect 12571 53431 12657 53487
rect 12713 53431 12799 53487
rect 12855 53431 12941 53487
rect 12997 53431 13083 53487
rect 13139 53431 13225 53487
rect 13281 53431 13367 53487
rect 13423 53431 13509 53487
rect 13565 53431 13651 53487
rect 13707 53431 13793 53487
rect 13849 53431 13935 53487
rect 13991 53431 14077 53487
rect 14133 53431 14219 53487
rect 14275 53431 14361 53487
rect 14417 53431 14503 53487
rect 14559 53431 14645 53487
rect 14701 53431 14787 53487
rect 14843 53431 14853 53487
rect 151 53345 14853 53431
rect 151 53289 161 53345
rect 217 53289 303 53345
rect 359 53289 445 53345
rect 501 53289 587 53345
rect 643 53289 729 53345
rect 785 53289 871 53345
rect 927 53289 1013 53345
rect 1069 53289 1155 53345
rect 1211 53289 1297 53345
rect 1353 53289 1439 53345
rect 1495 53289 1581 53345
rect 1637 53289 1723 53345
rect 1779 53289 1865 53345
rect 1921 53289 2007 53345
rect 2063 53289 2149 53345
rect 2205 53289 2291 53345
rect 2347 53289 2433 53345
rect 2489 53289 2575 53345
rect 2631 53289 2717 53345
rect 2773 53289 2859 53345
rect 2915 53289 3001 53345
rect 3057 53289 3143 53345
rect 3199 53289 3285 53345
rect 3341 53289 3427 53345
rect 3483 53289 3569 53345
rect 3625 53289 3711 53345
rect 3767 53289 3853 53345
rect 3909 53289 3995 53345
rect 4051 53289 4137 53345
rect 4193 53289 4279 53345
rect 4335 53289 4421 53345
rect 4477 53289 4563 53345
rect 4619 53289 4705 53345
rect 4761 53289 4847 53345
rect 4903 53289 4989 53345
rect 5045 53289 5131 53345
rect 5187 53289 5273 53345
rect 5329 53289 5415 53345
rect 5471 53289 5557 53345
rect 5613 53289 5699 53345
rect 5755 53289 5841 53345
rect 5897 53289 5983 53345
rect 6039 53289 6125 53345
rect 6181 53289 6267 53345
rect 6323 53289 6409 53345
rect 6465 53289 6551 53345
rect 6607 53289 6693 53345
rect 6749 53289 6835 53345
rect 6891 53289 6977 53345
rect 7033 53289 7119 53345
rect 7175 53289 7261 53345
rect 7317 53289 7403 53345
rect 7459 53289 7545 53345
rect 7601 53289 7687 53345
rect 7743 53289 7829 53345
rect 7885 53289 7971 53345
rect 8027 53289 8113 53345
rect 8169 53289 8255 53345
rect 8311 53289 8397 53345
rect 8453 53289 8539 53345
rect 8595 53289 8681 53345
rect 8737 53289 8823 53345
rect 8879 53289 8965 53345
rect 9021 53289 9107 53345
rect 9163 53289 9249 53345
rect 9305 53289 9391 53345
rect 9447 53289 9533 53345
rect 9589 53289 9675 53345
rect 9731 53289 9817 53345
rect 9873 53289 9959 53345
rect 10015 53289 10101 53345
rect 10157 53289 10243 53345
rect 10299 53289 10385 53345
rect 10441 53289 10527 53345
rect 10583 53289 10669 53345
rect 10725 53289 10811 53345
rect 10867 53289 10953 53345
rect 11009 53289 11095 53345
rect 11151 53289 11237 53345
rect 11293 53289 11379 53345
rect 11435 53289 11521 53345
rect 11577 53289 11663 53345
rect 11719 53289 11805 53345
rect 11861 53289 11947 53345
rect 12003 53289 12089 53345
rect 12145 53289 12231 53345
rect 12287 53289 12373 53345
rect 12429 53289 12515 53345
rect 12571 53289 12657 53345
rect 12713 53289 12799 53345
rect 12855 53289 12941 53345
rect 12997 53289 13083 53345
rect 13139 53289 13225 53345
rect 13281 53289 13367 53345
rect 13423 53289 13509 53345
rect 13565 53289 13651 53345
rect 13707 53289 13793 53345
rect 13849 53289 13935 53345
rect 13991 53289 14077 53345
rect 14133 53289 14219 53345
rect 14275 53289 14361 53345
rect 14417 53289 14503 53345
rect 14559 53289 14645 53345
rect 14701 53289 14787 53345
rect 14843 53289 14853 53345
rect 151 53203 14853 53289
rect 151 53147 161 53203
rect 217 53147 303 53203
rect 359 53147 445 53203
rect 501 53147 587 53203
rect 643 53147 729 53203
rect 785 53147 871 53203
rect 927 53147 1013 53203
rect 1069 53147 1155 53203
rect 1211 53147 1297 53203
rect 1353 53147 1439 53203
rect 1495 53147 1581 53203
rect 1637 53147 1723 53203
rect 1779 53147 1865 53203
rect 1921 53147 2007 53203
rect 2063 53147 2149 53203
rect 2205 53147 2291 53203
rect 2347 53147 2433 53203
rect 2489 53147 2575 53203
rect 2631 53147 2717 53203
rect 2773 53147 2859 53203
rect 2915 53147 3001 53203
rect 3057 53147 3143 53203
rect 3199 53147 3285 53203
rect 3341 53147 3427 53203
rect 3483 53147 3569 53203
rect 3625 53147 3711 53203
rect 3767 53147 3853 53203
rect 3909 53147 3995 53203
rect 4051 53147 4137 53203
rect 4193 53147 4279 53203
rect 4335 53147 4421 53203
rect 4477 53147 4563 53203
rect 4619 53147 4705 53203
rect 4761 53147 4847 53203
rect 4903 53147 4989 53203
rect 5045 53147 5131 53203
rect 5187 53147 5273 53203
rect 5329 53147 5415 53203
rect 5471 53147 5557 53203
rect 5613 53147 5699 53203
rect 5755 53147 5841 53203
rect 5897 53147 5983 53203
rect 6039 53147 6125 53203
rect 6181 53147 6267 53203
rect 6323 53147 6409 53203
rect 6465 53147 6551 53203
rect 6607 53147 6693 53203
rect 6749 53147 6835 53203
rect 6891 53147 6977 53203
rect 7033 53147 7119 53203
rect 7175 53147 7261 53203
rect 7317 53147 7403 53203
rect 7459 53147 7545 53203
rect 7601 53147 7687 53203
rect 7743 53147 7829 53203
rect 7885 53147 7971 53203
rect 8027 53147 8113 53203
rect 8169 53147 8255 53203
rect 8311 53147 8397 53203
rect 8453 53147 8539 53203
rect 8595 53147 8681 53203
rect 8737 53147 8823 53203
rect 8879 53147 8965 53203
rect 9021 53147 9107 53203
rect 9163 53147 9249 53203
rect 9305 53147 9391 53203
rect 9447 53147 9533 53203
rect 9589 53147 9675 53203
rect 9731 53147 9817 53203
rect 9873 53147 9959 53203
rect 10015 53147 10101 53203
rect 10157 53147 10243 53203
rect 10299 53147 10385 53203
rect 10441 53147 10527 53203
rect 10583 53147 10669 53203
rect 10725 53147 10811 53203
rect 10867 53147 10953 53203
rect 11009 53147 11095 53203
rect 11151 53147 11237 53203
rect 11293 53147 11379 53203
rect 11435 53147 11521 53203
rect 11577 53147 11663 53203
rect 11719 53147 11805 53203
rect 11861 53147 11947 53203
rect 12003 53147 12089 53203
rect 12145 53147 12231 53203
rect 12287 53147 12373 53203
rect 12429 53147 12515 53203
rect 12571 53147 12657 53203
rect 12713 53147 12799 53203
rect 12855 53147 12941 53203
rect 12997 53147 13083 53203
rect 13139 53147 13225 53203
rect 13281 53147 13367 53203
rect 13423 53147 13509 53203
rect 13565 53147 13651 53203
rect 13707 53147 13793 53203
rect 13849 53147 13935 53203
rect 13991 53147 14077 53203
rect 14133 53147 14219 53203
rect 14275 53147 14361 53203
rect 14417 53147 14503 53203
rect 14559 53147 14645 53203
rect 14701 53147 14787 53203
rect 14843 53147 14853 53203
rect 151 53061 14853 53147
rect 151 53005 161 53061
rect 217 53005 303 53061
rect 359 53005 445 53061
rect 501 53005 587 53061
rect 643 53005 729 53061
rect 785 53005 871 53061
rect 927 53005 1013 53061
rect 1069 53005 1155 53061
rect 1211 53005 1297 53061
rect 1353 53005 1439 53061
rect 1495 53005 1581 53061
rect 1637 53005 1723 53061
rect 1779 53005 1865 53061
rect 1921 53005 2007 53061
rect 2063 53005 2149 53061
rect 2205 53005 2291 53061
rect 2347 53005 2433 53061
rect 2489 53005 2575 53061
rect 2631 53005 2717 53061
rect 2773 53005 2859 53061
rect 2915 53005 3001 53061
rect 3057 53005 3143 53061
rect 3199 53005 3285 53061
rect 3341 53005 3427 53061
rect 3483 53005 3569 53061
rect 3625 53005 3711 53061
rect 3767 53005 3853 53061
rect 3909 53005 3995 53061
rect 4051 53005 4137 53061
rect 4193 53005 4279 53061
rect 4335 53005 4421 53061
rect 4477 53005 4563 53061
rect 4619 53005 4705 53061
rect 4761 53005 4847 53061
rect 4903 53005 4989 53061
rect 5045 53005 5131 53061
rect 5187 53005 5273 53061
rect 5329 53005 5415 53061
rect 5471 53005 5557 53061
rect 5613 53005 5699 53061
rect 5755 53005 5841 53061
rect 5897 53005 5983 53061
rect 6039 53005 6125 53061
rect 6181 53005 6267 53061
rect 6323 53005 6409 53061
rect 6465 53005 6551 53061
rect 6607 53005 6693 53061
rect 6749 53005 6835 53061
rect 6891 53005 6977 53061
rect 7033 53005 7119 53061
rect 7175 53005 7261 53061
rect 7317 53005 7403 53061
rect 7459 53005 7545 53061
rect 7601 53005 7687 53061
rect 7743 53005 7829 53061
rect 7885 53005 7971 53061
rect 8027 53005 8113 53061
rect 8169 53005 8255 53061
rect 8311 53005 8397 53061
rect 8453 53005 8539 53061
rect 8595 53005 8681 53061
rect 8737 53005 8823 53061
rect 8879 53005 8965 53061
rect 9021 53005 9107 53061
rect 9163 53005 9249 53061
rect 9305 53005 9391 53061
rect 9447 53005 9533 53061
rect 9589 53005 9675 53061
rect 9731 53005 9817 53061
rect 9873 53005 9959 53061
rect 10015 53005 10101 53061
rect 10157 53005 10243 53061
rect 10299 53005 10385 53061
rect 10441 53005 10527 53061
rect 10583 53005 10669 53061
rect 10725 53005 10811 53061
rect 10867 53005 10953 53061
rect 11009 53005 11095 53061
rect 11151 53005 11237 53061
rect 11293 53005 11379 53061
rect 11435 53005 11521 53061
rect 11577 53005 11663 53061
rect 11719 53005 11805 53061
rect 11861 53005 11947 53061
rect 12003 53005 12089 53061
rect 12145 53005 12231 53061
rect 12287 53005 12373 53061
rect 12429 53005 12515 53061
rect 12571 53005 12657 53061
rect 12713 53005 12799 53061
rect 12855 53005 12941 53061
rect 12997 53005 13083 53061
rect 13139 53005 13225 53061
rect 13281 53005 13367 53061
rect 13423 53005 13509 53061
rect 13565 53005 13651 53061
rect 13707 53005 13793 53061
rect 13849 53005 13935 53061
rect 13991 53005 14077 53061
rect 14133 53005 14219 53061
rect 14275 53005 14361 53061
rect 14417 53005 14503 53061
rect 14559 53005 14645 53061
rect 14701 53005 14787 53061
rect 14843 53005 14853 53061
rect 151 52919 14853 53005
rect 151 52863 161 52919
rect 217 52863 303 52919
rect 359 52863 445 52919
rect 501 52863 587 52919
rect 643 52863 729 52919
rect 785 52863 871 52919
rect 927 52863 1013 52919
rect 1069 52863 1155 52919
rect 1211 52863 1297 52919
rect 1353 52863 1439 52919
rect 1495 52863 1581 52919
rect 1637 52863 1723 52919
rect 1779 52863 1865 52919
rect 1921 52863 2007 52919
rect 2063 52863 2149 52919
rect 2205 52863 2291 52919
rect 2347 52863 2433 52919
rect 2489 52863 2575 52919
rect 2631 52863 2717 52919
rect 2773 52863 2859 52919
rect 2915 52863 3001 52919
rect 3057 52863 3143 52919
rect 3199 52863 3285 52919
rect 3341 52863 3427 52919
rect 3483 52863 3569 52919
rect 3625 52863 3711 52919
rect 3767 52863 3853 52919
rect 3909 52863 3995 52919
rect 4051 52863 4137 52919
rect 4193 52863 4279 52919
rect 4335 52863 4421 52919
rect 4477 52863 4563 52919
rect 4619 52863 4705 52919
rect 4761 52863 4847 52919
rect 4903 52863 4989 52919
rect 5045 52863 5131 52919
rect 5187 52863 5273 52919
rect 5329 52863 5415 52919
rect 5471 52863 5557 52919
rect 5613 52863 5699 52919
rect 5755 52863 5841 52919
rect 5897 52863 5983 52919
rect 6039 52863 6125 52919
rect 6181 52863 6267 52919
rect 6323 52863 6409 52919
rect 6465 52863 6551 52919
rect 6607 52863 6693 52919
rect 6749 52863 6835 52919
rect 6891 52863 6977 52919
rect 7033 52863 7119 52919
rect 7175 52863 7261 52919
rect 7317 52863 7403 52919
rect 7459 52863 7545 52919
rect 7601 52863 7687 52919
rect 7743 52863 7829 52919
rect 7885 52863 7971 52919
rect 8027 52863 8113 52919
rect 8169 52863 8255 52919
rect 8311 52863 8397 52919
rect 8453 52863 8539 52919
rect 8595 52863 8681 52919
rect 8737 52863 8823 52919
rect 8879 52863 8965 52919
rect 9021 52863 9107 52919
rect 9163 52863 9249 52919
rect 9305 52863 9391 52919
rect 9447 52863 9533 52919
rect 9589 52863 9675 52919
rect 9731 52863 9817 52919
rect 9873 52863 9959 52919
rect 10015 52863 10101 52919
rect 10157 52863 10243 52919
rect 10299 52863 10385 52919
rect 10441 52863 10527 52919
rect 10583 52863 10669 52919
rect 10725 52863 10811 52919
rect 10867 52863 10953 52919
rect 11009 52863 11095 52919
rect 11151 52863 11237 52919
rect 11293 52863 11379 52919
rect 11435 52863 11521 52919
rect 11577 52863 11663 52919
rect 11719 52863 11805 52919
rect 11861 52863 11947 52919
rect 12003 52863 12089 52919
rect 12145 52863 12231 52919
rect 12287 52863 12373 52919
rect 12429 52863 12515 52919
rect 12571 52863 12657 52919
rect 12713 52863 12799 52919
rect 12855 52863 12941 52919
rect 12997 52863 13083 52919
rect 13139 52863 13225 52919
rect 13281 52863 13367 52919
rect 13423 52863 13509 52919
rect 13565 52863 13651 52919
rect 13707 52863 13793 52919
rect 13849 52863 13935 52919
rect 13991 52863 14077 52919
rect 14133 52863 14219 52919
rect 14275 52863 14361 52919
rect 14417 52863 14503 52919
rect 14559 52863 14645 52919
rect 14701 52863 14787 52919
rect 14843 52863 14853 52919
rect 151 52777 14853 52863
rect 151 52721 161 52777
rect 217 52721 303 52777
rect 359 52721 445 52777
rect 501 52721 587 52777
rect 643 52721 729 52777
rect 785 52721 871 52777
rect 927 52721 1013 52777
rect 1069 52721 1155 52777
rect 1211 52721 1297 52777
rect 1353 52721 1439 52777
rect 1495 52721 1581 52777
rect 1637 52721 1723 52777
rect 1779 52721 1865 52777
rect 1921 52721 2007 52777
rect 2063 52721 2149 52777
rect 2205 52721 2291 52777
rect 2347 52721 2433 52777
rect 2489 52721 2575 52777
rect 2631 52721 2717 52777
rect 2773 52721 2859 52777
rect 2915 52721 3001 52777
rect 3057 52721 3143 52777
rect 3199 52721 3285 52777
rect 3341 52721 3427 52777
rect 3483 52721 3569 52777
rect 3625 52721 3711 52777
rect 3767 52721 3853 52777
rect 3909 52721 3995 52777
rect 4051 52721 4137 52777
rect 4193 52721 4279 52777
rect 4335 52721 4421 52777
rect 4477 52721 4563 52777
rect 4619 52721 4705 52777
rect 4761 52721 4847 52777
rect 4903 52721 4989 52777
rect 5045 52721 5131 52777
rect 5187 52721 5273 52777
rect 5329 52721 5415 52777
rect 5471 52721 5557 52777
rect 5613 52721 5699 52777
rect 5755 52721 5841 52777
rect 5897 52721 5983 52777
rect 6039 52721 6125 52777
rect 6181 52721 6267 52777
rect 6323 52721 6409 52777
rect 6465 52721 6551 52777
rect 6607 52721 6693 52777
rect 6749 52721 6835 52777
rect 6891 52721 6977 52777
rect 7033 52721 7119 52777
rect 7175 52721 7261 52777
rect 7317 52721 7403 52777
rect 7459 52721 7545 52777
rect 7601 52721 7687 52777
rect 7743 52721 7829 52777
rect 7885 52721 7971 52777
rect 8027 52721 8113 52777
rect 8169 52721 8255 52777
rect 8311 52721 8397 52777
rect 8453 52721 8539 52777
rect 8595 52721 8681 52777
rect 8737 52721 8823 52777
rect 8879 52721 8965 52777
rect 9021 52721 9107 52777
rect 9163 52721 9249 52777
rect 9305 52721 9391 52777
rect 9447 52721 9533 52777
rect 9589 52721 9675 52777
rect 9731 52721 9817 52777
rect 9873 52721 9959 52777
rect 10015 52721 10101 52777
rect 10157 52721 10243 52777
rect 10299 52721 10385 52777
rect 10441 52721 10527 52777
rect 10583 52721 10669 52777
rect 10725 52721 10811 52777
rect 10867 52721 10953 52777
rect 11009 52721 11095 52777
rect 11151 52721 11237 52777
rect 11293 52721 11379 52777
rect 11435 52721 11521 52777
rect 11577 52721 11663 52777
rect 11719 52721 11805 52777
rect 11861 52721 11947 52777
rect 12003 52721 12089 52777
rect 12145 52721 12231 52777
rect 12287 52721 12373 52777
rect 12429 52721 12515 52777
rect 12571 52721 12657 52777
rect 12713 52721 12799 52777
rect 12855 52721 12941 52777
rect 12997 52721 13083 52777
rect 13139 52721 13225 52777
rect 13281 52721 13367 52777
rect 13423 52721 13509 52777
rect 13565 52721 13651 52777
rect 13707 52721 13793 52777
rect 13849 52721 13935 52777
rect 13991 52721 14077 52777
rect 14133 52721 14219 52777
rect 14275 52721 14361 52777
rect 14417 52721 14503 52777
rect 14559 52721 14645 52777
rect 14701 52721 14787 52777
rect 14843 52721 14853 52777
rect 151 52635 14853 52721
rect 151 52579 161 52635
rect 217 52579 303 52635
rect 359 52579 445 52635
rect 501 52579 587 52635
rect 643 52579 729 52635
rect 785 52579 871 52635
rect 927 52579 1013 52635
rect 1069 52579 1155 52635
rect 1211 52579 1297 52635
rect 1353 52579 1439 52635
rect 1495 52579 1581 52635
rect 1637 52579 1723 52635
rect 1779 52579 1865 52635
rect 1921 52579 2007 52635
rect 2063 52579 2149 52635
rect 2205 52579 2291 52635
rect 2347 52579 2433 52635
rect 2489 52579 2575 52635
rect 2631 52579 2717 52635
rect 2773 52579 2859 52635
rect 2915 52579 3001 52635
rect 3057 52579 3143 52635
rect 3199 52579 3285 52635
rect 3341 52579 3427 52635
rect 3483 52579 3569 52635
rect 3625 52579 3711 52635
rect 3767 52579 3853 52635
rect 3909 52579 3995 52635
rect 4051 52579 4137 52635
rect 4193 52579 4279 52635
rect 4335 52579 4421 52635
rect 4477 52579 4563 52635
rect 4619 52579 4705 52635
rect 4761 52579 4847 52635
rect 4903 52579 4989 52635
rect 5045 52579 5131 52635
rect 5187 52579 5273 52635
rect 5329 52579 5415 52635
rect 5471 52579 5557 52635
rect 5613 52579 5699 52635
rect 5755 52579 5841 52635
rect 5897 52579 5983 52635
rect 6039 52579 6125 52635
rect 6181 52579 6267 52635
rect 6323 52579 6409 52635
rect 6465 52579 6551 52635
rect 6607 52579 6693 52635
rect 6749 52579 6835 52635
rect 6891 52579 6977 52635
rect 7033 52579 7119 52635
rect 7175 52579 7261 52635
rect 7317 52579 7403 52635
rect 7459 52579 7545 52635
rect 7601 52579 7687 52635
rect 7743 52579 7829 52635
rect 7885 52579 7971 52635
rect 8027 52579 8113 52635
rect 8169 52579 8255 52635
rect 8311 52579 8397 52635
rect 8453 52579 8539 52635
rect 8595 52579 8681 52635
rect 8737 52579 8823 52635
rect 8879 52579 8965 52635
rect 9021 52579 9107 52635
rect 9163 52579 9249 52635
rect 9305 52579 9391 52635
rect 9447 52579 9533 52635
rect 9589 52579 9675 52635
rect 9731 52579 9817 52635
rect 9873 52579 9959 52635
rect 10015 52579 10101 52635
rect 10157 52579 10243 52635
rect 10299 52579 10385 52635
rect 10441 52579 10527 52635
rect 10583 52579 10669 52635
rect 10725 52579 10811 52635
rect 10867 52579 10953 52635
rect 11009 52579 11095 52635
rect 11151 52579 11237 52635
rect 11293 52579 11379 52635
rect 11435 52579 11521 52635
rect 11577 52579 11663 52635
rect 11719 52579 11805 52635
rect 11861 52579 11947 52635
rect 12003 52579 12089 52635
rect 12145 52579 12231 52635
rect 12287 52579 12373 52635
rect 12429 52579 12515 52635
rect 12571 52579 12657 52635
rect 12713 52579 12799 52635
rect 12855 52579 12941 52635
rect 12997 52579 13083 52635
rect 13139 52579 13225 52635
rect 13281 52579 13367 52635
rect 13423 52579 13509 52635
rect 13565 52579 13651 52635
rect 13707 52579 13793 52635
rect 13849 52579 13935 52635
rect 13991 52579 14077 52635
rect 14133 52579 14219 52635
rect 14275 52579 14361 52635
rect 14417 52579 14503 52635
rect 14559 52579 14645 52635
rect 14701 52579 14787 52635
rect 14843 52579 14853 52635
rect 151 52493 14853 52579
rect 151 52437 161 52493
rect 217 52437 303 52493
rect 359 52437 445 52493
rect 501 52437 587 52493
rect 643 52437 729 52493
rect 785 52437 871 52493
rect 927 52437 1013 52493
rect 1069 52437 1155 52493
rect 1211 52437 1297 52493
rect 1353 52437 1439 52493
rect 1495 52437 1581 52493
rect 1637 52437 1723 52493
rect 1779 52437 1865 52493
rect 1921 52437 2007 52493
rect 2063 52437 2149 52493
rect 2205 52437 2291 52493
rect 2347 52437 2433 52493
rect 2489 52437 2575 52493
rect 2631 52437 2717 52493
rect 2773 52437 2859 52493
rect 2915 52437 3001 52493
rect 3057 52437 3143 52493
rect 3199 52437 3285 52493
rect 3341 52437 3427 52493
rect 3483 52437 3569 52493
rect 3625 52437 3711 52493
rect 3767 52437 3853 52493
rect 3909 52437 3995 52493
rect 4051 52437 4137 52493
rect 4193 52437 4279 52493
rect 4335 52437 4421 52493
rect 4477 52437 4563 52493
rect 4619 52437 4705 52493
rect 4761 52437 4847 52493
rect 4903 52437 4989 52493
rect 5045 52437 5131 52493
rect 5187 52437 5273 52493
rect 5329 52437 5415 52493
rect 5471 52437 5557 52493
rect 5613 52437 5699 52493
rect 5755 52437 5841 52493
rect 5897 52437 5983 52493
rect 6039 52437 6125 52493
rect 6181 52437 6267 52493
rect 6323 52437 6409 52493
rect 6465 52437 6551 52493
rect 6607 52437 6693 52493
rect 6749 52437 6835 52493
rect 6891 52437 6977 52493
rect 7033 52437 7119 52493
rect 7175 52437 7261 52493
rect 7317 52437 7403 52493
rect 7459 52437 7545 52493
rect 7601 52437 7687 52493
rect 7743 52437 7829 52493
rect 7885 52437 7971 52493
rect 8027 52437 8113 52493
rect 8169 52437 8255 52493
rect 8311 52437 8397 52493
rect 8453 52437 8539 52493
rect 8595 52437 8681 52493
rect 8737 52437 8823 52493
rect 8879 52437 8965 52493
rect 9021 52437 9107 52493
rect 9163 52437 9249 52493
rect 9305 52437 9391 52493
rect 9447 52437 9533 52493
rect 9589 52437 9675 52493
rect 9731 52437 9817 52493
rect 9873 52437 9959 52493
rect 10015 52437 10101 52493
rect 10157 52437 10243 52493
rect 10299 52437 10385 52493
rect 10441 52437 10527 52493
rect 10583 52437 10669 52493
rect 10725 52437 10811 52493
rect 10867 52437 10953 52493
rect 11009 52437 11095 52493
rect 11151 52437 11237 52493
rect 11293 52437 11379 52493
rect 11435 52437 11521 52493
rect 11577 52437 11663 52493
rect 11719 52437 11805 52493
rect 11861 52437 11947 52493
rect 12003 52437 12089 52493
rect 12145 52437 12231 52493
rect 12287 52437 12373 52493
rect 12429 52437 12515 52493
rect 12571 52437 12657 52493
rect 12713 52437 12799 52493
rect 12855 52437 12941 52493
rect 12997 52437 13083 52493
rect 13139 52437 13225 52493
rect 13281 52437 13367 52493
rect 13423 52437 13509 52493
rect 13565 52437 13651 52493
rect 13707 52437 13793 52493
rect 13849 52437 13935 52493
rect 13991 52437 14077 52493
rect 14133 52437 14219 52493
rect 14275 52437 14361 52493
rect 14417 52437 14503 52493
rect 14559 52437 14645 52493
rect 14701 52437 14787 52493
rect 14843 52437 14853 52493
rect 151 52427 14853 52437
rect 151 52163 14853 52173
rect 151 52107 161 52163
rect 217 52107 303 52163
rect 359 52107 445 52163
rect 501 52107 587 52163
rect 643 52107 729 52163
rect 785 52107 871 52163
rect 927 52107 1013 52163
rect 1069 52107 1155 52163
rect 1211 52107 1297 52163
rect 1353 52107 1439 52163
rect 1495 52107 1581 52163
rect 1637 52107 1723 52163
rect 1779 52107 1865 52163
rect 1921 52107 2007 52163
rect 2063 52107 2149 52163
rect 2205 52107 2291 52163
rect 2347 52107 2433 52163
rect 2489 52107 2575 52163
rect 2631 52107 2717 52163
rect 2773 52107 2859 52163
rect 2915 52107 3001 52163
rect 3057 52107 3143 52163
rect 3199 52107 3285 52163
rect 3341 52107 3427 52163
rect 3483 52107 3569 52163
rect 3625 52107 3711 52163
rect 3767 52107 3853 52163
rect 3909 52107 3995 52163
rect 4051 52107 4137 52163
rect 4193 52107 4279 52163
rect 4335 52107 4421 52163
rect 4477 52107 4563 52163
rect 4619 52107 4705 52163
rect 4761 52107 4847 52163
rect 4903 52107 4989 52163
rect 5045 52107 5131 52163
rect 5187 52107 5273 52163
rect 5329 52107 5415 52163
rect 5471 52107 5557 52163
rect 5613 52107 5699 52163
rect 5755 52107 5841 52163
rect 5897 52107 5983 52163
rect 6039 52107 6125 52163
rect 6181 52107 6267 52163
rect 6323 52107 6409 52163
rect 6465 52107 6551 52163
rect 6607 52107 6693 52163
rect 6749 52107 6835 52163
rect 6891 52107 6977 52163
rect 7033 52107 7119 52163
rect 7175 52107 7261 52163
rect 7317 52107 7403 52163
rect 7459 52107 7545 52163
rect 7601 52107 7687 52163
rect 7743 52107 7829 52163
rect 7885 52107 7971 52163
rect 8027 52107 8113 52163
rect 8169 52107 8255 52163
rect 8311 52107 8397 52163
rect 8453 52107 8539 52163
rect 8595 52107 8681 52163
rect 8737 52107 8823 52163
rect 8879 52107 8965 52163
rect 9021 52107 9107 52163
rect 9163 52107 9249 52163
rect 9305 52107 9391 52163
rect 9447 52107 9533 52163
rect 9589 52107 9675 52163
rect 9731 52107 9817 52163
rect 9873 52107 9959 52163
rect 10015 52107 10101 52163
rect 10157 52107 10243 52163
rect 10299 52107 10385 52163
rect 10441 52107 10527 52163
rect 10583 52107 10669 52163
rect 10725 52107 10811 52163
rect 10867 52107 10953 52163
rect 11009 52107 11095 52163
rect 11151 52107 11237 52163
rect 11293 52107 11379 52163
rect 11435 52107 11521 52163
rect 11577 52107 11663 52163
rect 11719 52107 11805 52163
rect 11861 52107 11947 52163
rect 12003 52107 12089 52163
rect 12145 52107 12231 52163
rect 12287 52107 12373 52163
rect 12429 52107 12515 52163
rect 12571 52107 12657 52163
rect 12713 52107 12799 52163
rect 12855 52107 12941 52163
rect 12997 52107 13083 52163
rect 13139 52107 13225 52163
rect 13281 52107 13367 52163
rect 13423 52107 13509 52163
rect 13565 52107 13651 52163
rect 13707 52107 13793 52163
rect 13849 52107 13935 52163
rect 13991 52107 14077 52163
rect 14133 52107 14219 52163
rect 14275 52107 14361 52163
rect 14417 52107 14503 52163
rect 14559 52107 14645 52163
rect 14701 52107 14787 52163
rect 14843 52107 14853 52163
rect 151 52021 14853 52107
rect 151 51965 161 52021
rect 217 51965 303 52021
rect 359 51965 445 52021
rect 501 51965 587 52021
rect 643 51965 729 52021
rect 785 51965 871 52021
rect 927 51965 1013 52021
rect 1069 51965 1155 52021
rect 1211 51965 1297 52021
rect 1353 51965 1439 52021
rect 1495 51965 1581 52021
rect 1637 51965 1723 52021
rect 1779 51965 1865 52021
rect 1921 51965 2007 52021
rect 2063 51965 2149 52021
rect 2205 51965 2291 52021
rect 2347 51965 2433 52021
rect 2489 51965 2575 52021
rect 2631 51965 2717 52021
rect 2773 51965 2859 52021
rect 2915 51965 3001 52021
rect 3057 51965 3143 52021
rect 3199 51965 3285 52021
rect 3341 51965 3427 52021
rect 3483 51965 3569 52021
rect 3625 51965 3711 52021
rect 3767 51965 3853 52021
rect 3909 51965 3995 52021
rect 4051 51965 4137 52021
rect 4193 51965 4279 52021
rect 4335 51965 4421 52021
rect 4477 51965 4563 52021
rect 4619 51965 4705 52021
rect 4761 51965 4847 52021
rect 4903 51965 4989 52021
rect 5045 51965 5131 52021
rect 5187 51965 5273 52021
rect 5329 51965 5415 52021
rect 5471 51965 5557 52021
rect 5613 51965 5699 52021
rect 5755 51965 5841 52021
rect 5897 51965 5983 52021
rect 6039 51965 6125 52021
rect 6181 51965 6267 52021
rect 6323 51965 6409 52021
rect 6465 51965 6551 52021
rect 6607 51965 6693 52021
rect 6749 51965 6835 52021
rect 6891 51965 6977 52021
rect 7033 51965 7119 52021
rect 7175 51965 7261 52021
rect 7317 51965 7403 52021
rect 7459 51965 7545 52021
rect 7601 51965 7687 52021
rect 7743 51965 7829 52021
rect 7885 51965 7971 52021
rect 8027 51965 8113 52021
rect 8169 51965 8255 52021
rect 8311 51965 8397 52021
rect 8453 51965 8539 52021
rect 8595 51965 8681 52021
rect 8737 51965 8823 52021
rect 8879 51965 8965 52021
rect 9021 51965 9107 52021
rect 9163 51965 9249 52021
rect 9305 51965 9391 52021
rect 9447 51965 9533 52021
rect 9589 51965 9675 52021
rect 9731 51965 9817 52021
rect 9873 51965 9959 52021
rect 10015 51965 10101 52021
rect 10157 51965 10243 52021
rect 10299 51965 10385 52021
rect 10441 51965 10527 52021
rect 10583 51965 10669 52021
rect 10725 51965 10811 52021
rect 10867 51965 10953 52021
rect 11009 51965 11095 52021
rect 11151 51965 11237 52021
rect 11293 51965 11379 52021
rect 11435 51965 11521 52021
rect 11577 51965 11663 52021
rect 11719 51965 11805 52021
rect 11861 51965 11947 52021
rect 12003 51965 12089 52021
rect 12145 51965 12231 52021
rect 12287 51965 12373 52021
rect 12429 51965 12515 52021
rect 12571 51965 12657 52021
rect 12713 51965 12799 52021
rect 12855 51965 12941 52021
rect 12997 51965 13083 52021
rect 13139 51965 13225 52021
rect 13281 51965 13367 52021
rect 13423 51965 13509 52021
rect 13565 51965 13651 52021
rect 13707 51965 13793 52021
rect 13849 51965 13935 52021
rect 13991 51965 14077 52021
rect 14133 51965 14219 52021
rect 14275 51965 14361 52021
rect 14417 51965 14503 52021
rect 14559 51965 14645 52021
rect 14701 51965 14787 52021
rect 14843 51965 14853 52021
rect 151 51879 14853 51965
rect 151 51823 161 51879
rect 217 51823 303 51879
rect 359 51823 445 51879
rect 501 51823 587 51879
rect 643 51823 729 51879
rect 785 51823 871 51879
rect 927 51823 1013 51879
rect 1069 51823 1155 51879
rect 1211 51823 1297 51879
rect 1353 51823 1439 51879
rect 1495 51823 1581 51879
rect 1637 51823 1723 51879
rect 1779 51823 1865 51879
rect 1921 51823 2007 51879
rect 2063 51823 2149 51879
rect 2205 51823 2291 51879
rect 2347 51823 2433 51879
rect 2489 51823 2575 51879
rect 2631 51823 2717 51879
rect 2773 51823 2859 51879
rect 2915 51823 3001 51879
rect 3057 51823 3143 51879
rect 3199 51823 3285 51879
rect 3341 51823 3427 51879
rect 3483 51823 3569 51879
rect 3625 51823 3711 51879
rect 3767 51823 3853 51879
rect 3909 51823 3995 51879
rect 4051 51823 4137 51879
rect 4193 51823 4279 51879
rect 4335 51823 4421 51879
rect 4477 51823 4563 51879
rect 4619 51823 4705 51879
rect 4761 51823 4847 51879
rect 4903 51823 4989 51879
rect 5045 51823 5131 51879
rect 5187 51823 5273 51879
rect 5329 51823 5415 51879
rect 5471 51823 5557 51879
rect 5613 51823 5699 51879
rect 5755 51823 5841 51879
rect 5897 51823 5983 51879
rect 6039 51823 6125 51879
rect 6181 51823 6267 51879
rect 6323 51823 6409 51879
rect 6465 51823 6551 51879
rect 6607 51823 6693 51879
rect 6749 51823 6835 51879
rect 6891 51823 6977 51879
rect 7033 51823 7119 51879
rect 7175 51823 7261 51879
rect 7317 51823 7403 51879
rect 7459 51823 7545 51879
rect 7601 51823 7687 51879
rect 7743 51823 7829 51879
rect 7885 51823 7971 51879
rect 8027 51823 8113 51879
rect 8169 51823 8255 51879
rect 8311 51823 8397 51879
rect 8453 51823 8539 51879
rect 8595 51823 8681 51879
rect 8737 51823 8823 51879
rect 8879 51823 8965 51879
rect 9021 51823 9107 51879
rect 9163 51823 9249 51879
rect 9305 51823 9391 51879
rect 9447 51823 9533 51879
rect 9589 51823 9675 51879
rect 9731 51823 9817 51879
rect 9873 51823 9959 51879
rect 10015 51823 10101 51879
rect 10157 51823 10243 51879
rect 10299 51823 10385 51879
rect 10441 51823 10527 51879
rect 10583 51823 10669 51879
rect 10725 51823 10811 51879
rect 10867 51823 10953 51879
rect 11009 51823 11095 51879
rect 11151 51823 11237 51879
rect 11293 51823 11379 51879
rect 11435 51823 11521 51879
rect 11577 51823 11663 51879
rect 11719 51823 11805 51879
rect 11861 51823 11947 51879
rect 12003 51823 12089 51879
rect 12145 51823 12231 51879
rect 12287 51823 12373 51879
rect 12429 51823 12515 51879
rect 12571 51823 12657 51879
rect 12713 51823 12799 51879
rect 12855 51823 12941 51879
rect 12997 51823 13083 51879
rect 13139 51823 13225 51879
rect 13281 51823 13367 51879
rect 13423 51823 13509 51879
rect 13565 51823 13651 51879
rect 13707 51823 13793 51879
rect 13849 51823 13935 51879
rect 13991 51823 14077 51879
rect 14133 51823 14219 51879
rect 14275 51823 14361 51879
rect 14417 51823 14503 51879
rect 14559 51823 14645 51879
rect 14701 51823 14787 51879
rect 14843 51823 14853 51879
rect 151 51737 14853 51823
rect 151 51681 161 51737
rect 217 51681 303 51737
rect 359 51681 445 51737
rect 501 51681 587 51737
rect 643 51681 729 51737
rect 785 51681 871 51737
rect 927 51681 1013 51737
rect 1069 51681 1155 51737
rect 1211 51681 1297 51737
rect 1353 51681 1439 51737
rect 1495 51681 1581 51737
rect 1637 51681 1723 51737
rect 1779 51681 1865 51737
rect 1921 51681 2007 51737
rect 2063 51681 2149 51737
rect 2205 51681 2291 51737
rect 2347 51681 2433 51737
rect 2489 51681 2575 51737
rect 2631 51681 2717 51737
rect 2773 51681 2859 51737
rect 2915 51681 3001 51737
rect 3057 51681 3143 51737
rect 3199 51681 3285 51737
rect 3341 51681 3427 51737
rect 3483 51681 3569 51737
rect 3625 51681 3711 51737
rect 3767 51681 3853 51737
rect 3909 51681 3995 51737
rect 4051 51681 4137 51737
rect 4193 51681 4279 51737
rect 4335 51681 4421 51737
rect 4477 51681 4563 51737
rect 4619 51681 4705 51737
rect 4761 51681 4847 51737
rect 4903 51681 4989 51737
rect 5045 51681 5131 51737
rect 5187 51681 5273 51737
rect 5329 51681 5415 51737
rect 5471 51681 5557 51737
rect 5613 51681 5699 51737
rect 5755 51681 5841 51737
rect 5897 51681 5983 51737
rect 6039 51681 6125 51737
rect 6181 51681 6267 51737
rect 6323 51681 6409 51737
rect 6465 51681 6551 51737
rect 6607 51681 6693 51737
rect 6749 51681 6835 51737
rect 6891 51681 6977 51737
rect 7033 51681 7119 51737
rect 7175 51681 7261 51737
rect 7317 51681 7403 51737
rect 7459 51681 7545 51737
rect 7601 51681 7687 51737
rect 7743 51681 7829 51737
rect 7885 51681 7971 51737
rect 8027 51681 8113 51737
rect 8169 51681 8255 51737
rect 8311 51681 8397 51737
rect 8453 51681 8539 51737
rect 8595 51681 8681 51737
rect 8737 51681 8823 51737
rect 8879 51681 8965 51737
rect 9021 51681 9107 51737
rect 9163 51681 9249 51737
rect 9305 51681 9391 51737
rect 9447 51681 9533 51737
rect 9589 51681 9675 51737
rect 9731 51681 9817 51737
rect 9873 51681 9959 51737
rect 10015 51681 10101 51737
rect 10157 51681 10243 51737
rect 10299 51681 10385 51737
rect 10441 51681 10527 51737
rect 10583 51681 10669 51737
rect 10725 51681 10811 51737
rect 10867 51681 10953 51737
rect 11009 51681 11095 51737
rect 11151 51681 11237 51737
rect 11293 51681 11379 51737
rect 11435 51681 11521 51737
rect 11577 51681 11663 51737
rect 11719 51681 11805 51737
rect 11861 51681 11947 51737
rect 12003 51681 12089 51737
rect 12145 51681 12231 51737
rect 12287 51681 12373 51737
rect 12429 51681 12515 51737
rect 12571 51681 12657 51737
rect 12713 51681 12799 51737
rect 12855 51681 12941 51737
rect 12997 51681 13083 51737
rect 13139 51681 13225 51737
rect 13281 51681 13367 51737
rect 13423 51681 13509 51737
rect 13565 51681 13651 51737
rect 13707 51681 13793 51737
rect 13849 51681 13935 51737
rect 13991 51681 14077 51737
rect 14133 51681 14219 51737
rect 14275 51681 14361 51737
rect 14417 51681 14503 51737
rect 14559 51681 14645 51737
rect 14701 51681 14787 51737
rect 14843 51681 14853 51737
rect 151 51595 14853 51681
rect 151 51539 161 51595
rect 217 51539 303 51595
rect 359 51539 445 51595
rect 501 51539 587 51595
rect 643 51539 729 51595
rect 785 51539 871 51595
rect 927 51539 1013 51595
rect 1069 51539 1155 51595
rect 1211 51539 1297 51595
rect 1353 51539 1439 51595
rect 1495 51539 1581 51595
rect 1637 51539 1723 51595
rect 1779 51539 1865 51595
rect 1921 51539 2007 51595
rect 2063 51539 2149 51595
rect 2205 51539 2291 51595
rect 2347 51539 2433 51595
rect 2489 51539 2575 51595
rect 2631 51539 2717 51595
rect 2773 51539 2859 51595
rect 2915 51539 3001 51595
rect 3057 51539 3143 51595
rect 3199 51539 3285 51595
rect 3341 51539 3427 51595
rect 3483 51539 3569 51595
rect 3625 51539 3711 51595
rect 3767 51539 3853 51595
rect 3909 51539 3995 51595
rect 4051 51539 4137 51595
rect 4193 51539 4279 51595
rect 4335 51539 4421 51595
rect 4477 51539 4563 51595
rect 4619 51539 4705 51595
rect 4761 51539 4847 51595
rect 4903 51539 4989 51595
rect 5045 51539 5131 51595
rect 5187 51539 5273 51595
rect 5329 51539 5415 51595
rect 5471 51539 5557 51595
rect 5613 51539 5699 51595
rect 5755 51539 5841 51595
rect 5897 51539 5983 51595
rect 6039 51539 6125 51595
rect 6181 51539 6267 51595
rect 6323 51539 6409 51595
rect 6465 51539 6551 51595
rect 6607 51539 6693 51595
rect 6749 51539 6835 51595
rect 6891 51539 6977 51595
rect 7033 51539 7119 51595
rect 7175 51539 7261 51595
rect 7317 51539 7403 51595
rect 7459 51539 7545 51595
rect 7601 51539 7687 51595
rect 7743 51539 7829 51595
rect 7885 51539 7971 51595
rect 8027 51539 8113 51595
rect 8169 51539 8255 51595
rect 8311 51539 8397 51595
rect 8453 51539 8539 51595
rect 8595 51539 8681 51595
rect 8737 51539 8823 51595
rect 8879 51539 8965 51595
rect 9021 51539 9107 51595
rect 9163 51539 9249 51595
rect 9305 51539 9391 51595
rect 9447 51539 9533 51595
rect 9589 51539 9675 51595
rect 9731 51539 9817 51595
rect 9873 51539 9959 51595
rect 10015 51539 10101 51595
rect 10157 51539 10243 51595
rect 10299 51539 10385 51595
rect 10441 51539 10527 51595
rect 10583 51539 10669 51595
rect 10725 51539 10811 51595
rect 10867 51539 10953 51595
rect 11009 51539 11095 51595
rect 11151 51539 11237 51595
rect 11293 51539 11379 51595
rect 11435 51539 11521 51595
rect 11577 51539 11663 51595
rect 11719 51539 11805 51595
rect 11861 51539 11947 51595
rect 12003 51539 12089 51595
rect 12145 51539 12231 51595
rect 12287 51539 12373 51595
rect 12429 51539 12515 51595
rect 12571 51539 12657 51595
rect 12713 51539 12799 51595
rect 12855 51539 12941 51595
rect 12997 51539 13083 51595
rect 13139 51539 13225 51595
rect 13281 51539 13367 51595
rect 13423 51539 13509 51595
rect 13565 51539 13651 51595
rect 13707 51539 13793 51595
rect 13849 51539 13935 51595
rect 13991 51539 14077 51595
rect 14133 51539 14219 51595
rect 14275 51539 14361 51595
rect 14417 51539 14503 51595
rect 14559 51539 14645 51595
rect 14701 51539 14787 51595
rect 14843 51539 14853 51595
rect 151 51453 14853 51539
rect 151 51397 161 51453
rect 217 51397 303 51453
rect 359 51397 445 51453
rect 501 51397 587 51453
rect 643 51397 729 51453
rect 785 51397 871 51453
rect 927 51397 1013 51453
rect 1069 51397 1155 51453
rect 1211 51397 1297 51453
rect 1353 51397 1439 51453
rect 1495 51397 1581 51453
rect 1637 51397 1723 51453
rect 1779 51397 1865 51453
rect 1921 51397 2007 51453
rect 2063 51397 2149 51453
rect 2205 51397 2291 51453
rect 2347 51397 2433 51453
rect 2489 51397 2575 51453
rect 2631 51397 2717 51453
rect 2773 51397 2859 51453
rect 2915 51397 3001 51453
rect 3057 51397 3143 51453
rect 3199 51397 3285 51453
rect 3341 51397 3427 51453
rect 3483 51397 3569 51453
rect 3625 51397 3711 51453
rect 3767 51397 3853 51453
rect 3909 51397 3995 51453
rect 4051 51397 4137 51453
rect 4193 51397 4279 51453
rect 4335 51397 4421 51453
rect 4477 51397 4563 51453
rect 4619 51397 4705 51453
rect 4761 51397 4847 51453
rect 4903 51397 4989 51453
rect 5045 51397 5131 51453
rect 5187 51397 5273 51453
rect 5329 51397 5415 51453
rect 5471 51397 5557 51453
rect 5613 51397 5699 51453
rect 5755 51397 5841 51453
rect 5897 51397 5983 51453
rect 6039 51397 6125 51453
rect 6181 51397 6267 51453
rect 6323 51397 6409 51453
rect 6465 51397 6551 51453
rect 6607 51397 6693 51453
rect 6749 51397 6835 51453
rect 6891 51397 6977 51453
rect 7033 51397 7119 51453
rect 7175 51397 7261 51453
rect 7317 51397 7403 51453
rect 7459 51397 7545 51453
rect 7601 51397 7687 51453
rect 7743 51397 7829 51453
rect 7885 51397 7971 51453
rect 8027 51397 8113 51453
rect 8169 51397 8255 51453
rect 8311 51397 8397 51453
rect 8453 51397 8539 51453
rect 8595 51397 8681 51453
rect 8737 51397 8823 51453
rect 8879 51397 8965 51453
rect 9021 51397 9107 51453
rect 9163 51397 9249 51453
rect 9305 51397 9391 51453
rect 9447 51397 9533 51453
rect 9589 51397 9675 51453
rect 9731 51397 9817 51453
rect 9873 51397 9959 51453
rect 10015 51397 10101 51453
rect 10157 51397 10243 51453
rect 10299 51397 10385 51453
rect 10441 51397 10527 51453
rect 10583 51397 10669 51453
rect 10725 51397 10811 51453
rect 10867 51397 10953 51453
rect 11009 51397 11095 51453
rect 11151 51397 11237 51453
rect 11293 51397 11379 51453
rect 11435 51397 11521 51453
rect 11577 51397 11663 51453
rect 11719 51397 11805 51453
rect 11861 51397 11947 51453
rect 12003 51397 12089 51453
rect 12145 51397 12231 51453
rect 12287 51397 12373 51453
rect 12429 51397 12515 51453
rect 12571 51397 12657 51453
rect 12713 51397 12799 51453
rect 12855 51397 12941 51453
rect 12997 51397 13083 51453
rect 13139 51397 13225 51453
rect 13281 51397 13367 51453
rect 13423 51397 13509 51453
rect 13565 51397 13651 51453
rect 13707 51397 13793 51453
rect 13849 51397 13935 51453
rect 13991 51397 14077 51453
rect 14133 51397 14219 51453
rect 14275 51397 14361 51453
rect 14417 51397 14503 51453
rect 14559 51397 14645 51453
rect 14701 51397 14787 51453
rect 14843 51397 14853 51453
rect 151 51311 14853 51397
rect 151 51255 161 51311
rect 217 51255 303 51311
rect 359 51255 445 51311
rect 501 51255 587 51311
rect 643 51255 729 51311
rect 785 51255 871 51311
rect 927 51255 1013 51311
rect 1069 51255 1155 51311
rect 1211 51255 1297 51311
rect 1353 51255 1439 51311
rect 1495 51255 1581 51311
rect 1637 51255 1723 51311
rect 1779 51255 1865 51311
rect 1921 51255 2007 51311
rect 2063 51255 2149 51311
rect 2205 51255 2291 51311
rect 2347 51255 2433 51311
rect 2489 51255 2575 51311
rect 2631 51255 2717 51311
rect 2773 51255 2859 51311
rect 2915 51255 3001 51311
rect 3057 51255 3143 51311
rect 3199 51255 3285 51311
rect 3341 51255 3427 51311
rect 3483 51255 3569 51311
rect 3625 51255 3711 51311
rect 3767 51255 3853 51311
rect 3909 51255 3995 51311
rect 4051 51255 4137 51311
rect 4193 51255 4279 51311
rect 4335 51255 4421 51311
rect 4477 51255 4563 51311
rect 4619 51255 4705 51311
rect 4761 51255 4847 51311
rect 4903 51255 4989 51311
rect 5045 51255 5131 51311
rect 5187 51255 5273 51311
rect 5329 51255 5415 51311
rect 5471 51255 5557 51311
rect 5613 51255 5699 51311
rect 5755 51255 5841 51311
rect 5897 51255 5983 51311
rect 6039 51255 6125 51311
rect 6181 51255 6267 51311
rect 6323 51255 6409 51311
rect 6465 51255 6551 51311
rect 6607 51255 6693 51311
rect 6749 51255 6835 51311
rect 6891 51255 6977 51311
rect 7033 51255 7119 51311
rect 7175 51255 7261 51311
rect 7317 51255 7403 51311
rect 7459 51255 7545 51311
rect 7601 51255 7687 51311
rect 7743 51255 7829 51311
rect 7885 51255 7971 51311
rect 8027 51255 8113 51311
rect 8169 51255 8255 51311
rect 8311 51255 8397 51311
rect 8453 51255 8539 51311
rect 8595 51255 8681 51311
rect 8737 51255 8823 51311
rect 8879 51255 8965 51311
rect 9021 51255 9107 51311
rect 9163 51255 9249 51311
rect 9305 51255 9391 51311
rect 9447 51255 9533 51311
rect 9589 51255 9675 51311
rect 9731 51255 9817 51311
rect 9873 51255 9959 51311
rect 10015 51255 10101 51311
rect 10157 51255 10243 51311
rect 10299 51255 10385 51311
rect 10441 51255 10527 51311
rect 10583 51255 10669 51311
rect 10725 51255 10811 51311
rect 10867 51255 10953 51311
rect 11009 51255 11095 51311
rect 11151 51255 11237 51311
rect 11293 51255 11379 51311
rect 11435 51255 11521 51311
rect 11577 51255 11663 51311
rect 11719 51255 11805 51311
rect 11861 51255 11947 51311
rect 12003 51255 12089 51311
rect 12145 51255 12231 51311
rect 12287 51255 12373 51311
rect 12429 51255 12515 51311
rect 12571 51255 12657 51311
rect 12713 51255 12799 51311
rect 12855 51255 12941 51311
rect 12997 51255 13083 51311
rect 13139 51255 13225 51311
rect 13281 51255 13367 51311
rect 13423 51255 13509 51311
rect 13565 51255 13651 51311
rect 13707 51255 13793 51311
rect 13849 51255 13935 51311
rect 13991 51255 14077 51311
rect 14133 51255 14219 51311
rect 14275 51255 14361 51311
rect 14417 51255 14503 51311
rect 14559 51255 14645 51311
rect 14701 51255 14787 51311
rect 14843 51255 14853 51311
rect 151 51169 14853 51255
rect 151 51113 161 51169
rect 217 51113 303 51169
rect 359 51113 445 51169
rect 501 51113 587 51169
rect 643 51113 729 51169
rect 785 51113 871 51169
rect 927 51113 1013 51169
rect 1069 51113 1155 51169
rect 1211 51113 1297 51169
rect 1353 51113 1439 51169
rect 1495 51113 1581 51169
rect 1637 51113 1723 51169
rect 1779 51113 1865 51169
rect 1921 51113 2007 51169
rect 2063 51113 2149 51169
rect 2205 51113 2291 51169
rect 2347 51113 2433 51169
rect 2489 51113 2575 51169
rect 2631 51113 2717 51169
rect 2773 51113 2859 51169
rect 2915 51113 3001 51169
rect 3057 51113 3143 51169
rect 3199 51113 3285 51169
rect 3341 51113 3427 51169
rect 3483 51113 3569 51169
rect 3625 51113 3711 51169
rect 3767 51113 3853 51169
rect 3909 51113 3995 51169
rect 4051 51113 4137 51169
rect 4193 51113 4279 51169
rect 4335 51113 4421 51169
rect 4477 51113 4563 51169
rect 4619 51113 4705 51169
rect 4761 51113 4847 51169
rect 4903 51113 4989 51169
rect 5045 51113 5131 51169
rect 5187 51113 5273 51169
rect 5329 51113 5415 51169
rect 5471 51113 5557 51169
rect 5613 51113 5699 51169
rect 5755 51113 5841 51169
rect 5897 51113 5983 51169
rect 6039 51113 6125 51169
rect 6181 51113 6267 51169
rect 6323 51113 6409 51169
rect 6465 51113 6551 51169
rect 6607 51113 6693 51169
rect 6749 51113 6835 51169
rect 6891 51113 6977 51169
rect 7033 51113 7119 51169
rect 7175 51113 7261 51169
rect 7317 51113 7403 51169
rect 7459 51113 7545 51169
rect 7601 51113 7687 51169
rect 7743 51113 7829 51169
rect 7885 51113 7971 51169
rect 8027 51113 8113 51169
rect 8169 51113 8255 51169
rect 8311 51113 8397 51169
rect 8453 51113 8539 51169
rect 8595 51113 8681 51169
rect 8737 51113 8823 51169
rect 8879 51113 8965 51169
rect 9021 51113 9107 51169
rect 9163 51113 9249 51169
rect 9305 51113 9391 51169
rect 9447 51113 9533 51169
rect 9589 51113 9675 51169
rect 9731 51113 9817 51169
rect 9873 51113 9959 51169
rect 10015 51113 10101 51169
rect 10157 51113 10243 51169
rect 10299 51113 10385 51169
rect 10441 51113 10527 51169
rect 10583 51113 10669 51169
rect 10725 51113 10811 51169
rect 10867 51113 10953 51169
rect 11009 51113 11095 51169
rect 11151 51113 11237 51169
rect 11293 51113 11379 51169
rect 11435 51113 11521 51169
rect 11577 51113 11663 51169
rect 11719 51113 11805 51169
rect 11861 51113 11947 51169
rect 12003 51113 12089 51169
rect 12145 51113 12231 51169
rect 12287 51113 12373 51169
rect 12429 51113 12515 51169
rect 12571 51113 12657 51169
rect 12713 51113 12799 51169
rect 12855 51113 12941 51169
rect 12997 51113 13083 51169
rect 13139 51113 13225 51169
rect 13281 51113 13367 51169
rect 13423 51113 13509 51169
rect 13565 51113 13651 51169
rect 13707 51113 13793 51169
rect 13849 51113 13935 51169
rect 13991 51113 14077 51169
rect 14133 51113 14219 51169
rect 14275 51113 14361 51169
rect 14417 51113 14503 51169
rect 14559 51113 14645 51169
rect 14701 51113 14787 51169
rect 14843 51113 14853 51169
rect 151 51027 14853 51113
rect 151 50971 161 51027
rect 217 50971 303 51027
rect 359 50971 445 51027
rect 501 50971 587 51027
rect 643 50971 729 51027
rect 785 50971 871 51027
rect 927 50971 1013 51027
rect 1069 50971 1155 51027
rect 1211 50971 1297 51027
rect 1353 50971 1439 51027
rect 1495 50971 1581 51027
rect 1637 50971 1723 51027
rect 1779 50971 1865 51027
rect 1921 50971 2007 51027
rect 2063 50971 2149 51027
rect 2205 50971 2291 51027
rect 2347 50971 2433 51027
rect 2489 50971 2575 51027
rect 2631 50971 2717 51027
rect 2773 50971 2859 51027
rect 2915 50971 3001 51027
rect 3057 50971 3143 51027
rect 3199 50971 3285 51027
rect 3341 50971 3427 51027
rect 3483 50971 3569 51027
rect 3625 50971 3711 51027
rect 3767 50971 3853 51027
rect 3909 50971 3995 51027
rect 4051 50971 4137 51027
rect 4193 50971 4279 51027
rect 4335 50971 4421 51027
rect 4477 50971 4563 51027
rect 4619 50971 4705 51027
rect 4761 50971 4847 51027
rect 4903 50971 4989 51027
rect 5045 50971 5131 51027
rect 5187 50971 5273 51027
rect 5329 50971 5415 51027
rect 5471 50971 5557 51027
rect 5613 50971 5699 51027
rect 5755 50971 5841 51027
rect 5897 50971 5983 51027
rect 6039 50971 6125 51027
rect 6181 50971 6267 51027
rect 6323 50971 6409 51027
rect 6465 50971 6551 51027
rect 6607 50971 6693 51027
rect 6749 50971 6835 51027
rect 6891 50971 6977 51027
rect 7033 50971 7119 51027
rect 7175 50971 7261 51027
rect 7317 50971 7403 51027
rect 7459 50971 7545 51027
rect 7601 50971 7687 51027
rect 7743 50971 7829 51027
rect 7885 50971 7971 51027
rect 8027 50971 8113 51027
rect 8169 50971 8255 51027
rect 8311 50971 8397 51027
rect 8453 50971 8539 51027
rect 8595 50971 8681 51027
rect 8737 50971 8823 51027
rect 8879 50971 8965 51027
rect 9021 50971 9107 51027
rect 9163 50971 9249 51027
rect 9305 50971 9391 51027
rect 9447 50971 9533 51027
rect 9589 50971 9675 51027
rect 9731 50971 9817 51027
rect 9873 50971 9959 51027
rect 10015 50971 10101 51027
rect 10157 50971 10243 51027
rect 10299 50971 10385 51027
rect 10441 50971 10527 51027
rect 10583 50971 10669 51027
rect 10725 50971 10811 51027
rect 10867 50971 10953 51027
rect 11009 50971 11095 51027
rect 11151 50971 11237 51027
rect 11293 50971 11379 51027
rect 11435 50971 11521 51027
rect 11577 50971 11663 51027
rect 11719 50971 11805 51027
rect 11861 50971 11947 51027
rect 12003 50971 12089 51027
rect 12145 50971 12231 51027
rect 12287 50971 12373 51027
rect 12429 50971 12515 51027
rect 12571 50971 12657 51027
rect 12713 50971 12799 51027
rect 12855 50971 12941 51027
rect 12997 50971 13083 51027
rect 13139 50971 13225 51027
rect 13281 50971 13367 51027
rect 13423 50971 13509 51027
rect 13565 50971 13651 51027
rect 13707 50971 13793 51027
rect 13849 50971 13935 51027
rect 13991 50971 14077 51027
rect 14133 50971 14219 51027
rect 14275 50971 14361 51027
rect 14417 50971 14503 51027
rect 14559 50971 14645 51027
rect 14701 50971 14787 51027
rect 14843 50971 14853 51027
rect 151 50885 14853 50971
rect 151 50829 161 50885
rect 217 50829 303 50885
rect 359 50829 445 50885
rect 501 50829 587 50885
rect 643 50829 729 50885
rect 785 50829 871 50885
rect 927 50829 1013 50885
rect 1069 50829 1155 50885
rect 1211 50829 1297 50885
rect 1353 50829 1439 50885
rect 1495 50829 1581 50885
rect 1637 50829 1723 50885
rect 1779 50829 1865 50885
rect 1921 50829 2007 50885
rect 2063 50829 2149 50885
rect 2205 50829 2291 50885
rect 2347 50829 2433 50885
rect 2489 50829 2575 50885
rect 2631 50829 2717 50885
rect 2773 50829 2859 50885
rect 2915 50829 3001 50885
rect 3057 50829 3143 50885
rect 3199 50829 3285 50885
rect 3341 50829 3427 50885
rect 3483 50829 3569 50885
rect 3625 50829 3711 50885
rect 3767 50829 3853 50885
rect 3909 50829 3995 50885
rect 4051 50829 4137 50885
rect 4193 50829 4279 50885
rect 4335 50829 4421 50885
rect 4477 50829 4563 50885
rect 4619 50829 4705 50885
rect 4761 50829 4847 50885
rect 4903 50829 4989 50885
rect 5045 50829 5131 50885
rect 5187 50829 5273 50885
rect 5329 50829 5415 50885
rect 5471 50829 5557 50885
rect 5613 50829 5699 50885
rect 5755 50829 5841 50885
rect 5897 50829 5983 50885
rect 6039 50829 6125 50885
rect 6181 50829 6267 50885
rect 6323 50829 6409 50885
rect 6465 50829 6551 50885
rect 6607 50829 6693 50885
rect 6749 50829 6835 50885
rect 6891 50829 6977 50885
rect 7033 50829 7119 50885
rect 7175 50829 7261 50885
rect 7317 50829 7403 50885
rect 7459 50829 7545 50885
rect 7601 50829 7687 50885
rect 7743 50829 7829 50885
rect 7885 50829 7971 50885
rect 8027 50829 8113 50885
rect 8169 50829 8255 50885
rect 8311 50829 8397 50885
rect 8453 50829 8539 50885
rect 8595 50829 8681 50885
rect 8737 50829 8823 50885
rect 8879 50829 8965 50885
rect 9021 50829 9107 50885
rect 9163 50829 9249 50885
rect 9305 50829 9391 50885
rect 9447 50829 9533 50885
rect 9589 50829 9675 50885
rect 9731 50829 9817 50885
rect 9873 50829 9959 50885
rect 10015 50829 10101 50885
rect 10157 50829 10243 50885
rect 10299 50829 10385 50885
rect 10441 50829 10527 50885
rect 10583 50829 10669 50885
rect 10725 50829 10811 50885
rect 10867 50829 10953 50885
rect 11009 50829 11095 50885
rect 11151 50829 11237 50885
rect 11293 50829 11379 50885
rect 11435 50829 11521 50885
rect 11577 50829 11663 50885
rect 11719 50829 11805 50885
rect 11861 50829 11947 50885
rect 12003 50829 12089 50885
rect 12145 50829 12231 50885
rect 12287 50829 12373 50885
rect 12429 50829 12515 50885
rect 12571 50829 12657 50885
rect 12713 50829 12799 50885
rect 12855 50829 12941 50885
rect 12997 50829 13083 50885
rect 13139 50829 13225 50885
rect 13281 50829 13367 50885
rect 13423 50829 13509 50885
rect 13565 50829 13651 50885
rect 13707 50829 13793 50885
rect 13849 50829 13935 50885
rect 13991 50829 14077 50885
rect 14133 50829 14219 50885
rect 14275 50829 14361 50885
rect 14417 50829 14503 50885
rect 14559 50829 14645 50885
rect 14701 50829 14787 50885
rect 14843 50829 14853 50885
rect 151 50819 14853 50829
rect 151 50563 14853 50573
rect 151 50507 161 50563
rect 217 50507 303 50563
rect 359 50507 445 50563
rect 501 50507 587 50563
rect 643 50507 729 50563
rect 785 50507 871 50563
rect 927 50507 1013 50563
rect 1069 50507 1155 50563
rect 1211 50507 1297 50563
rect 1353 50507 1439 50563
rect 1495 50507 1581 50563
rect 1637 50507 1723 50563
rect 1779 50507 1865 50563
rect 1921 50507 2007 50563
rect 2063 50507 2149 50563
rect 2205 50507 2291 50563
rect 2347 50507 2433 50563
rect 2489 50507 2575 50563
rect 2631 50507 2717 50563
rect 2773 50507 2859 50563
rect 2915 50507 3001 50563
rect 3057 50507 3143 50563
rect 3199 50507 3285 50563
rect 3341 50507 3427 50563
rect 3483 50507 3569 50563
rect 3625 50507 3711 50563
rect 3767 50507 3853 50563
rect 3909 50507 3995 50563
rect 4051 50507 4137 50563
rect 4193 50507 4279 50563
rect 4335 50507 4421 50563
rect 4477 50507 4563 50563
rect 4619 50507 4705 50563
rect 4761 50507 4847 50563
rect 4903 50507 4989 50563
rect 5045 50507 5131 50563
rect 5187 50507 5273 50563
rect 5329 50507 5415 50563
rect 5471 50507 5557 50563
rect 5613 50507 5699 50563
rect 5755 50507 5841 50563
rect 5897 50507 5983 50563
rect 6039 50507 6125 50563
rect 6181 50507 6267 50563
rect 6323 50507 6409 50563
rect 6465 50507 6551 50563
rect 6607 50507 6693 50563
rect 6749 50507 6835 50563
rect 6891 50507 6977 50563
rect 7033 50507 7119 50563
rect 7175 50507 7261 50563
rect 7317 50507 7403 50563
rect 7459 50507 7545 50563
rect 7601 50507 7687 50563
rect 7743 50507 7829 50563
rect 7885 50507 7971 50563
rect 8027 50507 8113 50563
rect 8169 50507 8255 50563
rect 8311 50507 8397 50563
rect 8453 50507 8539 50563
rect 8595 50507 8681 50563
rect 8737 50507 8823 50563
rect 8879 50507 8965 50563
rect 9021 50507 9107 50563
rect 9163 50507 9249 50563
rect 9305 50507 9391 50563
rect 9447 50507 9533 50563
rect 9589 50507 9675 50563
rect 9731 50507 9817 50563
rect 9873 50507 9959 50563
rect 10015 50507 10101 50563
rect 10157 50507 10243 50563
rect 10299 50507 10385 50563
rect 10441 50507 10527 50563
rect 10583 50507 10669 50563
rect 10725 50507 10811 50563
rect 10867 50507 10953 50563
rect 11009 50507 11095 50563
rect 11151 50507 11237 50563
rect 11293 50507 11379 50563
rect 11435 50507 11521 50563
rect 11577 50507 11663 50563
rect 11719 50507 11805 50563
rect 11861 50507 11947 50563
rect 12003 50507 12089 50563
rect 12145 50507 12231 50563
rect 12287 50507 12373 50563
rect 12429 50507 12515 50563
rect 12571 50507 12657 50563
rect 12713 50507 12799 50563
rect 12855 50507 12941 50563
rect 12997 50507 13083 50563
rect 13139 50507 13225 50563
rect 13281 50507 13367 50563
rect 13423 50507 13509 50563
rect 13565 50507 13651 50563
rect 13707 50507 13793 50563
rect 13849 50507 13935 50563
rect 13991 50507 14077 50563
rect 14133 50507 14219 50563
rect 14275 50507 14361 50563
rect 14417 50507 14503 50563
rect 14559 50507 14645 50563
rect 14701 50507 14787 50563
rect 14843 50507 14853 50563
rect 151 50421 14853 50507
rect 151 50365 161 50421
rect 217 50365 303 50421
rect 359 50365 445 50421
rect 501 50365 587 50421
rect 643 50365 729 50421
rect 785 50365 871 50421
rect 927 50365 1013 50421
rect 1069 50365 1155 50421
rect 1211 50365 1297 50421
rect 1353 50365 1439 50421
rect 1495 50365 1581 50421
rect 1637 50365 1723 50421
rect 1779 50365 1865 50421
rect 1921 50365 2007 50421
rect 2063 50365 2149 50421
rect 2205 50365 2291 50421
rect 2347 50365 2433 50421
rect 2489 50365 2575 50421
rect 2631 50365 2717 50421
rect 2773 50365 2859 50421
rect 2915 50365 3001 50421
rect 3057 50365 3143 50421
rect 3199 50365 3285 50421
rect 3341 50365 3427 50421
rect 3483 50365 3569 50421
rect 3625 50365 3711 50421
rect 3767 50365 3853 50421
rect 3909 50365 3995 50421
rect 4051 50365 4137 50421
rect 4193 50365 4279 50421
rect 4335 50365 4421 50421
rect 4477 50365 4563 50421
rect 4619 50365 4705 50421
rect 4761 50365 4847 50421
rect 4903 50365 4989 50421
rect 5045 50365 5131 50421
rect 5187 50365 5273 50421
rect 5329 50365 5415 50421
rect 5471 50365 5557 50421
rect 5613 50365 5699 50421
rect 5755 50365 5841 50421
rect 5897 50365 5983 50421
rect 6039 50365 6125 50421
rect 6181 50365 6267 50421
rect 6323 50365 6409 50421
rect 6465 50365 6551 50421
rect 6607 50365 6693 50421
rect 6749 50365 6835 50421
rect 6891 50365 6977 50421
rect 7033 50365 7119 50421
rect 7175 50365 7261 50421
rect 7317 50365 7403 50421
rect 7459 50365 7545 50421
rect 7601 50365 7687 50421
rect 7743 50365 7829 50421
rect 7885 50365 7971 50421
rect 8027 50365 8113 50421
rect 8169 50365 8255 50421
rect 8311 50365 8397 50421
rect 8453 50365 8539 50421
rect 8595 50365 8681 50421
rect 8737 50365 8823 50421
rect 8879 50365 8965 50421
rect 9021 50365 9107 50421
rect 9163 50365 9249 50421
rect 9305 50365 9391 50421
rect 9447 50365 9533 50421
rect 9589 50365 9675 50421
rect 9731 50365 9817 50421
rect 9873 50365 9959 50421
rect 10015 50365 10101 50421
rect 10157 50365 10243 50421
rect 10299 50365 10385 50421
rect 10441 50365 10527 50421
rect 10583 50365 10669 50421
rect 10725 50365 10811 50421
rect 10867 50365 10953 50421
rect 11009 50365 11095 50421
rect 11151 50365 11237 50421
rect 11293 50365 11379 50421
rect 11435 50365 11521 50421
rect 11577 50365 11663 50421
rect 11719 50365 11805 50421
rect 11861 50365 11947 50421
rect 12003 50365 12089 50421
rect 12145 50365 12231 50421
rect 12287 50365 12373 50421
rect 12429 50365 12515 50421
rect 12571 50365 12657 50421
rect 12713 50365 12799 50421
rect 12855 50365 12941 50421
rect 12997 50365 13083 50421
rect 13139 50365 13225 50421
rect 13281 50365 13367 50421
rect 13423 50365 13509 50421
rect 13565 50365 13651 50421
rect 13707 50365 13793 50421
rect 13849 50365 13935 50421
rect 13991 50365 14077 50421
rect 14133 50365 14219 50421
rect 14275 50365 14361 50421
rect 14417 50365 14503 50421
rect 14559 50365 14645 50421
rect 14701 50365 14787 50421
rect 14843 50365 14853 50421
rect 151 50279 14853 50365
rect 151 50223 161 50279
rect 217 50223 303 50279
rect 359 50223 445 50279
rect 501 50223 587 50279
rect 643 50223 729 50279
rect 785 50223 871 50279
rect 927 50223 1013 50279
rect 1069 50223 1155 50279
rect 1211 50223 1297 50279
rect 1353 50223 1439 50279
rect 1495 50223 1581 50279
rect 1637 50223 1723 50279
rect 1779 50223 1865 50279
rect 1921 50223 2007 50279
rect 2063 50223 2149 50279
rect 2205 50223 2291 50279
rect 2347 50223 2433 50279
rect 2489 50223 2575 50279
rect 2631 50223 2717 50279
rect 2773 50223 2859 50279
rect 2915 50223 3001 50279
rect 3057 50223 3143 50279
rect 3199 50223 3285 50279
rect 3341 50223 3427 50279
rect 3483 50223 3569 50279
rect 3625 50223 3711 50279
rect 3767 50223 3853 50279
rect 3909 50223 3995 50279
rect 4051 50223 4137 50279
rect 4193 50223 4279 50279
rect 4335 50223 4421 50279
rect 4477 50223 4563 50279
rect 4619 50223 4705 50279
rect 4761 50223 4847 50279
rect 4903 50223 4989 50279
rect 5045 50223 5131 50279
rect 5187 50223 5273 50279
rect 5329 50223 5415 50279
rect 5471 50223 5557 50279
rect 5613 50223 5699 50279
rect 5755 50223 5841 50279
rect 5897 50223 5983 50279
rect 6039 50223 6125 50279
rect 6181 50223 6267 50279
rect 6323 50223 6409 50279
rect 6465 50223 6551 50279
rect 6607 50223 6693 50279
rect 6749 50223 6835 50279
rect 6891 50223 6977 50279
rect 7033 50223 7119 50279
rect 7175 50223 7261 50279
rect 7317 50223 7403 50279
rect 7459 50223 7545 50279
rect 7601 50223 7687 50279
rect 7743 50223 7829 50279
rect 7885 50223 7971 50279
rect 8027 50223 8113 50279
rect 8169 50223 8255 50279
rect 8311 50223 8397 50279
rect 8453 50223 8539 50279
rect 8595 50223 8681 50279
rect 8737 50223 8823 50279
rect 8879 50223 8965 50279
rect 9021 50223 9107 50279
rect 9163 50223 9249 50279
rect 9305 50223 9391 50279
rect 9447 50223 9533 50279
rect 9589 50223 9675 50279
rect 9731 50223 9817 50279
rect 9873 50223 9959 50279
rect 10015 50223 10101 50279
rect 10157 50223 10243 50279
rect 10299 50223 10385 50279
rect 10441 50223 10527 50279
rect 10583 50223 10669 50279
rect 10725 50223 10811 50279
rect 10867 50223 10953 50279
rect 11009 50223 11095 50279
rect 11151 50223 11237 50279
rect 11293 50223 11379 50279
rect 11435 50223 11521 50279
rect 11577 50223 11663 50279
rect 11719 50223 11805 50279
rect 11861 50223 11947 50279
rect 12003 50223 12089 50279
rect 12145 50223 12231 50279
rect 12287 50223 12373 50279
rect 12429 50223 12515 50279
rect 12571 50223 12657 50279
rect 12713 50223 12799 50279
rect 12855 50223 12941 50279
rect 12997 50223 13083 50279
rect 13139 50223 13225 50279
rect 13281 50223 13367 50279
rect 13423 50223 13509 50279
rect 13565 50223 13651 50279
rect 13707 50223 13793 50279
rect 13849 50223 13935 50279
rect 13991 50223 14077 50279
rect 14133 50223 14219 50279
rect 14275 50223 14361 50279
rect 14417 50223 14503 50279
rect 14559 50223 14645 50279
rect 14701 50223 14787 50279
rect 14843 50223 14853 50279
rect 151 50137 14853 50223
rect 151 50081 161 50137
rect 217 50081 303 50137
rect 359 50081 445 50137
rect 501 50081 587 50137
rect 643 50081 729 50137
rect 785 50081 871 50137
rect 927 50081 1013 50137
rect 1069 50081 1155 50137
rect 1211 50081 1297 50137
rect 1353 50081 1439 50137
rect 1495 50081 1581 50137
rect 1637 50081 1723 50137
rect 1779 50081 1865 50137
rect 1921 50081 2007 50137
rect 2063 50081 2149 50137
rect 2205 50081 2291 50137
rect 2347 50081 2433 50137
rect 2489 50081 2575 50137
rect 2631 50081 2717 50137
rect 2773 50081 2859 50137
rect 2915 50081 3001 50137
rect 3057 50081 3143 50137
rect 3199 50081 3285 50137
rect 3341 50081 3427 50137
rect 3483 50081 3569 50137
rect 3625 50081 3711 50137
rect 3767 50081 3853 50137
rect 3909 50081 3995 50137
rect 4051 50081 4137 50137
rect 4193 50081 4279 50137
rect 4335 50081 4421 50137
rect 4477 50081 4563 50137
rect 4619 50081 4705 50137
rect 4761 50081 4847 50137
rect 4903 50081 4989 50137
rect 5045 50081 5131 50137
rect 5187 50081 5273 50137
rect 5329 50081 5415 50137
rect 5471 50081 5557 50137
rect 5613 50081 5699 50137
rect 5755 50081 5841 50137
rect 5897 50081 5983 50137
rect 6039 50081 6125 50137
rect 6181 50081 6267 50137
rect 6323 50081 6409 50137
rect 6465 50081 6551 50137
rect 6607 50081 6693 50137
rect 6749 50081 6835 50137
rect 6891 50081 6977 50137
rect 7033 50081 7119 50137
rect 7175 50081 7261 50137
rect 7317 50081 7403 50137
rect 7459 50081 7545 50137
rect 7601 50081 7687 50137
rect 7743 50081 7829 50137
rect 7885 50081 7971 50137
rect 8027 50081 8113 50137
rect 8169 50081 8255 50137
rect 8311 50081 8397 50137
rect 8453 50081 8539 50137
rect 8595 50081 8681 50137
rect 8737 50081 8823 50137
rect 8879 50081 8965 50137
rect 9021 50081 9107 50137
rect 9163 50081 9249 50137
rect 9305 50081 9391 50137
rect 9447 50081 9533 50137
rect 9589 50081 9675 50137
rect 9731 50081 9817 50137
rect 9873 50081 9959 50137
rect 10015 50081 10101 50137
rect 10157 50081 10243 50137
rect 10299 50081 10385 50137
rect 10441 50081 10527 50137
rect 10583 50081 10669 50137
rect 10725 50081 10811 50137
rect 10867 50081 10953 50137
rect 11009 50081 11095 50137
rect 11151 50081 11237 50137
rect 11293 50081 11379 50137
rect 11435 50081 11521 50137
rect 11577 50081 11663 50137
rect 11719 50081 11805 50137
rect 11861 50081 11947 50137
rect 12003 50081 12089 50137
rect 12145 50081 12231 50137
rect 12287 50081 12373 50137
rect 12429 50081 12515 50137
rect 12571 50081 12657 50137
rect 12713 50081 12799 50137
rect 12855 50081 12941 50137
rect 12997 50081 13083 50137
rect 13139 50081 13225 50137
rect 13281 50081 13367 50137
rect 13423 50081 13509 50137
rect 13565 50081 13651 50137
rect 13707 50081 13793 50137
rect 13849 50081 13935 50137
rect 13991 50081 14077 50137
rect 14133 50081 14219 50137
rect 14275 50081 14361 50137
rect 14417 50081 14503 50137
rect 14559 50081 14645 50137
rect 14701 50081 14787 50137
rect 14843 50081 14853 50137
rect 151 49995 14853 50081
rect 151 49939 161 49995
rect 217 49939 303 49995
rect 359 49939 445 49995
rect 501 49939 587 49995
rect 643 49939 729 49995
rect 785 49939 871 49995
rect 927 49939 1013 49995
rect 1069 49939 1155 49995
rect 1211 49939 1297 49995
rect 1353 49939 1439 49995
rect 1495 49939 1581 49995
rect 1637 49939 1723 49995
rect 1779 49939 1865 49995
rect 1921 49939 2007 49995
rect 2063 49939 2149 49995
rect 2205 49939 2291 49995
rect 2347 49939 2433 49995
rect 2489 49939 2575 49995
rect 2631 49939 2717 49995
rect 2773 49939 2859 49995
rect 2915 49939 3001 49995
rect 3057 49939 3143 49995
rect 3199 49939 3285 49995
rect 3341 49939 3427 49995
rect 3483 49939 3569 49995
rect 3625 49939 3711 49995
rect 3767 49939 3853 49995
rect 3909 49939 3995 49995
rect 4051 49939 4137 49995
rect 4193 49939 4279 49995
rect 4335 49939 4421 49995
rect 4477 49939 4563 49995
rect 4619 49939 4705 49995
rect 4761 49939 4847 49995
rect 4903 49939 4989 49995
rect 5045 49939 5131 49995
rect 5187 49939 5273 49995
rect 5329 49939 5415 49995
rect 5471 49939 5557 49995
rect 5613 49939 5699 49995
rect 5755 49939 5841 49995
rect 5897 49939 5983 49995
rect 6039 49939 6125 49995
rect 6181 49939 6267 49995
rect 6323 49939 6409 49995
rect 6465 49939 6551 49995
rect 6607 49939 6693 49995
rect 6749 49939 6835 49995
rect 6891 49939 6977 49995
rect 7033 49939 7119 49995
rect 7175 49939 7261 49995
rect 7317 49939 7403 49995
rect 7459 49939 7545 49995
rect 7601 49939 7687 49995
rect 7743 49939 7829 49995
rect 7885 49939 7971 49995
rect 8027 49939 8113 49995
rect 8169 49939 8255 49995
rect 8311 49939 8397 49995
rect 8453 49939 8539 49995
rect 8595 49939 8681 49995
rect 8737 49939 8823 49995
rect 8879 49939 8965 49995
rect 9021 49939 9107 49995
rect 9163 49939 9249 49995
rect 9305 49939 9391 49995
rect 9447 49939 9533 49995
rect 9589 49939 9675 49995
rect 9731 49939 9817 49995
rect 9873 49939 9959 49995
rect 10015 49939 10101 49995
rect 10157 49939 10243 49995
rect 10299 49939 10385 49995
rect 10441 49939 10527 49995
rect 10583 49939 10669 49995
rect 10725 49939 10811 49995
rect 10867 49939 10953 49995
rect 11009 49939 11095 49995
rect 11151 49939 11237 49995
rect 11293 49939 11379 49995
rect 11435 49939 11521 49995
rect 11577 49939 11663 49995
rect 11719 49939 11805 49995
rect 11861 49939 11947 49995
rect 12003 49939 12089 49995
rect 12145 49939 12231 49995
rect 12287 49939 12373 49995
rect 12429 49939 12515 49995
rect 12571 49939 12657 49995
rect 12713 49939 12799 49995
rect 12855 49939 12941 49995
rect 12997 49939 13083 49995
rect 13139 49939 13225 49995
rect 13281 49939 13367 49995
rect 13423 49939 13509 49995
rect 13565 49939 13651 49995
rect 13707 49939 13793 49995
rect 13849 49939 13935 49995
rect 13991 49939 14077 49995
rect 14133 49939 14219 49995
rect 14275 49939 14361 49995
rect 14417 49939 14503 49995
rect 14559 49939 14645 49995
rect 14701 49939 14787 49995
rect 14843 49939 14853 49995
rect 151 49853 14853 49939
rect 151 49797 161 49853
rect 217 49797 303 49853
rect 359 49797 445 49853
rect 501 49797 587 49853
rect 643 49797 729 49853
rect 785 49797 871 49853
rect 927 49797 1013 49853
rect 1069 49797 1155 49853
rect 1211 49797 1297 49853
rect 1353 49797 1439 49853
rect 1495 49797 1581 49853
rect 1637 49797 1723 49853
rect 1779 49797 1865 49853
rect 1921 49797 2007 49853
rect 2063 49797 2149 49853
rect 2205 49797 2291 49853
rect 2347 49797 2433 49853
rect 2489 49797 2575 49853
rect 2631 49797 2717 49853
rect 2773 49797 2859 49853
rect 2915 49797 3001 49853
rect 3057 49797 3143 49853
rect 3199 49797 3285 49853
rect 3341 49797 3427 49853
rect 3483 49797 3569 49853
rect 3625 49797 3711 49853
rect 3767 49797 3853 49853
rect 3909 49797 3995 49853
rect 4051 49797 4137 49853
rect 4193 49797 4279 49853
rect 4335 49797 4421 49853
rect 4477 49797 4563 49853
rect 4619 49797 4705 49853
rect 4761 49797 4847 49853
rect 4903 49797 4989 49853
rect 5045 49797 5131 49853
rect 5187 49797 5273 49853
rect 5329 49797 5415 49853
rect 5471 49797 5557 49853
rect 5613 49797 5699 49853
rect 5755 49797 5841 49853
rect 5897 49797 5983 49853
rect 6039 49797 6125 49853
rect 6181 49797 6267 49853
rect 6323 49797 6409 49853
rect 6465 49797 6551 49853
rect 6607 49797 6693 49853
rect 6749 49797 6835 49853
rect 6891 49797 6977 49853
rect 7033 49797 7119 49853
rect 7175 49797 7261 49853
rect 7317 49797 7403 49853
rect 7459 49797 7545 49853
rect 7601 49797 7687 49853
rect 7743 49797 7829 49853
rect 7885 49797 7971 49853
rect 8027 49797 8113 49853
rect 8169 49797 8255 49853
rect 8311 49797 8397 49853
rect 8453 49797 8539 49853
rect 8595 49797 8681 49853
rect 8737 49797 8823 49853
rect 8879 49797 8965 49853
rect 9021 49797 9107 49853
rect 9163 49797 9249 49853
rect 9305 49797 9391 49853
rect 9447 49797 9533 49853
rect 9589 49797 9675 49853
rect 9731 49797 9817 49853
rect 9873 49797 9959 49853
rect 10015 49797 10101 49853
rect 10157 49797 10243 49853
rect 10299 49797 10385 49853
rect 10441 49797 10527 49853
rect 10583 49797 10669 49853
rect 10725 49797 10811 49853
rect 10867 49797 10953 49853
rect 11009 49797 11095 49853
rect 11151 49797 11237 49853
rect 11293 49797 11379 49853
rect 11435 49797 11521 49853
rect 11577 49797 11663 49853
rect 11719 49797 11805 49853
rect 11861 49797 11947 49853
rect 12003 49797 12089 49853
rect 12145 49797 12231 49853
rect 12287 49797 12373 49853
rect 12429 49797 12515 49853
rect 12571 49797 12657 49853
rect 12713 49797 12799 49853
rect 12855 49797 12941 49853
rect 12997 49797 13083 49853
rect 13139 49797 13225 49853
rect 13281 49797 13367 49853
rect 13423 49797 13509 49853
rect 13565 49797 13651 49853
rect 13707 49797 13793 49853
rect 13849 49797 13935 49853
rect 13991 49797 14077 49853
rect 14133 49797 14219 49853
rect 14275 49797 14361 49853
rect 14417 49797 14503 49853
rect 14559 49797 14645 49853
rect 14701 49797 14787 49853
rect 14843 49797 14853 49853
rect 151 49711 14853 49797
rect 151 49655 161 49711
rect 217 49655 303 49711
rect 359 49655 445 49711
rect 501 49655 587 49711
rect 643 49655 729 49711
rect 785 49655 871 49711
rect 927 49655 1013 49711
rect 1069 49655 1155 49711
rect 1211 49655 1297 49711
rect 1353 49655 1439 49711
rect 1495 49655 1581 49711
rect 1637 49655 1723 49711
rect 1779 49655 1865 49711
rect 1921 49655 2007 49711
rect 2063 49655 2149 49711
rect 2205 49655 2291 49711
rect 2347 49655 2433 49711
rect 2489 49655 2575 49711
rect 2631 49655 2717 49711
rect 2773 49655 2859 49711
rect 2915 49655 3001 49711
rect 3057 49655 3143 49711
rect 3199 49655 3285 49711
rect 3341 49655 3427 49711
rect 3483 49655 3569 49711
rect 3625 49655 3711 49711
rect 3767 49655 3853 49711
rect 3909 49655 3995 49711
rect 4051 49655 4137 49711
rect 4193 49655 4279 49711
rect 4335 49655 4421 49711
rect 4477 49655 4563 49711
rect 4619 49655 4705 49711
rect 4761 49655 4847 49711
rect 4903 49655 4989 49711
rect 5045 49655 5131 49711
rect 5187 49655 5273 49711
rect 5329 49655 5415 49711
rect 5471 49655 5557 49711
rect 5613 49655 5699 49711
rect 5755 49655 5841 49711
rect 5897 49655 5983 49711
rect 6039 49655 6125 49711
rect 6181 49655 6267 49711
rect 6323 49655 6409 49711
rect 6465 49655 6551 49711
rect 6607 49655 6693 49711
rect 6749 49655 6835 49711
rect 6891 49655 6977 49711
rect 7033 49655 7119 49711
rect 7175 49655 7261 49711
rect 7317 49655 7403 49711
rect 7459 49655 7545 49711
rect 7601 49655 7687 49711
rect 7743 49655 7829 49711
rect 7885 49655 7971 49711
rect 8027 49655 8113 49711
rect 8169 49655 8255 49711
rect 8311 49655 8397 49711
rect 8453 49655 8539 49711
rect 8595 49655 8681 49711
rect 8737 49655 8823 49711
rect 8879 49655 8965 49711
rect 9021 49655 9107 49711
rect 9163 49655 9249 49711
rect 9305 49655 9391 49711
rect 9447 49655 9533 49711
rect 9589 49655 9675 49711
rect 9731 49655 9817 49711
rect 9873 49655 9959 49711
rect 10015 49655 10101 49711
rect 10157 49655 10243 49711
rect 10299 49655 10385 49711
rect 10441 49655 10527 49711
rect 10583 49655 10669 49711
rect 10725 49655 10811 49711
rect 10867 49655 10953 49711
rect 11009 49655 11095 49711
rect 11151 49655 11237 49711
rect 11293 49655 11379 49711
rect 11435 49655 11521 49711
rect 11577 49655 11663 49711
rect 11719 49655 11805 49711
rect 11861 49655 11947 49711
rect 12003 49655 12089 49711
rect 12145 49655 12231 49711
rect 12287 49655 12373 49711
rect 12429 49655 12515 49711
rect 12571 49655 12657 49711
rect 12713 49655 12799 49711
rect 12855 49655 12941 49711
rect 12997 49655 13083 49711
rect 13139 49655 13225 49711
rect 13281 49655 13367 49711
rect 13423 49655 13509 49711
rect 13565 49655 13651 49711
rect 13707 49655 13793 49711
rect 13849 49655 13935 49711
rect 13991 49655 14077 49711
rect 14133 49655 14219 49711
rect 14275 49655 14361 49711
rect 14417 49655 14503 49711
rect 14559 49655 14645 49711
rect 14701 49655 14787 49711
rect 14843 49655 14853 49711
rect 151 49569 14853 49655
rect 151 49513 161 49569
rect 217 49513 303 49569
rect 359 49513 445 49569
rect 501 49513 587 49569
rect 643 49513 729 49569
rect 785 49513 871 49569
rect 927 49513 1013 49569
rect 1069 49513 1155 49569
rect 1211 49513 1297 49569
rect 1353 49513 1439 49569
rect 1495 49513 1581 49569
rect 1637 49513 1723 49569
rect 1779 49513 1865 49569
rect 1921 49513 2007 49569
rect 2063 49513 2149 49569
rect 2205 49513 2291 49569
rect 2347 49513 2433 49569
rect 2489 49513 2575 49569
rect 2631 49513 2717 49569
rect 2773 49513 2859 49569
rect 2915 49513 3001 49569
rect 3057 49513 3143 49569
rect 3199 49513 3285 49569
rect 3341 49513 3427 49569
rect 3483 49513 3569 49569
rect 3625 49513 3711 49569
rect 3767 49513 3853 49569
rect 3909 49513 3995 49569
rect 4051 49513 4137 49569
rect 4193 49513 4279 49569
rect 4335 49513 4421 49569
rect 4477 49513 4563 49569
rect 4619 49513 4705 49569
rect 4761 49513 4847 49569
rect 4903 49513 4989 49569
rect 5045 49513 5131 49569
rect 5187 49513 5273 49569
rect 5329 49513 5415 49569
rect 5471 49513 5557 49569
rect 5613 49513 5699 49569
rect 5755 49513 5841 49569
rect 5897 49513 5983 49569
rect 6039 49513 6125 49569
rect 6181 49513 6267 49569
rect 6323 49513 6409 49569
rect 6465 49513 6551 49569
rect 6607 49513 6693 49569
rect 6749 49513 6835 49569
rect 6891 49513 6977 49569
rect 7033 49513 7119 49569
rect 7175 49513 7261 49569
rect 7317 49513 7403 49569
rect 7459 49513 7545 49569
rect 7601 49513 7687 49569
rect 7743 49513 7829 49569
rect 7885 49513 7971 49569
rect 8027 49513 8113 49569
rect 8169 49513 8255 49569
rect 8311 49513 8397 49569
rect 8453 49513 8539 49569
rect 8595 49513 8681 49569
rect 8737 49513 8823 49569
rect 8879 49513 8965 49569
rect 9021 49513 9107 49569
rect 9163 49513 9249 49569
rect 9305 49513 9391 49569
rect 9447 49513 9533 49569
rect 9589 49513 9675 49569
rect 9731 49513 9817 49569
rect 9873 49513 9959 49569
rect 10015 49513 10101 49569
rect 10157 49513 10243 49569
rect 10299 49513 10385 49569
rect 10441 49513 10527 49569
rect 10583 49513 10669 49569
rect 10725 49513 10811 49569
rect 10867 49513 10953 49569
rect 11009 49513 11095 49569
rect 11151 49513 11237 49569
rect 11293 49513 11379 49569
rect 11435 49513 11521 49569
rect 11577 49513 11663 49569
rect 11719 49513 11805 49569
rect 11861 49513 11947 49569
rect 12003 49513 12089 49569
rect 12145 49513 12231 49569
rect 12287 49513 12373 49569
rect 12429 49513 12515 49569
rect 12571 49513 12657 49569
rect 12713 49513 12799 49569
rect 12855 49513 12941 49569
rect 12997 49513 13083 49569
rect 13139 49513 13225 49569
rect 13281 49513 13367 49569
rect 13423 49513 13509 49569
rect 13565 49513 13651 49569
rect 13707 49513 13793 49569
rect 13849 49513 13935 49569
rect 13991 49513 14077 49569
rect 14133 49513 14219 49569
rect 14275 49513 14361 49569
rect 14417 49513 14503 49569
rect 14559 49513 14645 49569
rect 14701 49513 14787 49569
rect 14843 49513 14853 49569
rect 151 49427 14853 49513
rect 151 49371 161 49427
rect 217 49371 303 49427
rect 359 49371 445 49427
rect 501 49371 587 49427
rect 643 49371 729 49427
rect 785 49371 871 49427
rect 927 49371 1013 49427
rect 1069 49371 1155 49427
rect 1211 49371 1297 49427
rect 1353 49371 1439 49427
rect 1495 49371 1581 49427
rect 1637 49371 1723 49427
rect 1779 49371 1865 49427
rect 1921 49371 2007 49427
rect 2063 49371 2149 49427
rect 2205 49371 2291 49427
rect 2347 49371 2433 49427
rect 2489 49371 2575 49427
rect 2631 49371 2717 49427
rect 2773 49371 2859 49427
rect 2915 49371 3001 49427
rect 3057 49371 3143 49427
rect 3199 49371 3285 49427
rect 3341 49371 3427 49427
rect 3483 49371 3569 49427
rect 3625 49371 3711 49427
rect 3767 49371 3853 49427
rect 3909 49371 3995 49427
rect 4051 49371 4137 49427
rect 4193 49371 4279 49427
rect 4335 49371 4421 49427
rect 4477 49371 4563 49427
rect 4619 49371 4705 49427
rect 4761 49371 4847 49427
rect 4903 49371 4989 49427
rect 5045 49371 5131 49427
rect 5187 49371 5273 49427
rect 5329 49371 5415 49427
rect 5471 49371 5557 49427
rect 5613 49371 5699 49427
rect 5755 49371 5841 49427
rect 5897 49371 5983 49427
rect 6039 49371 6125 49427
rect 6181 49371 6267 49427
rect 6323 49371 6409 49427
rect 6465 49371 6551 49427
rect 6607 49371 6693 49427
rect 6749 49371 6835 49427
rect 6891 49371 6977 49427
rect 7033 49371 7119 49427
rect 7175 49371 7261 49427
rect 7317 49371 7403 49427
rect 7459 49371 7545 49427
rect 7601 49371 7687 49427
rect 7743 49371 7829 49427
rect 7885 49371 7971 49427
rect 8027 49371 8113 49427
rect 8169 49371 8255 49427
rect 8311 49371 8397 49427
rect 8453 49371 8539 49427
rect 8595 49371 8681 49427
rect 8737 49371 8823 49427
rect 8879 49371 8965 49427
rect 9021 49371 9107 49427
rect 9163 49371 9249 49427
rect 9305 49371 9391 49427
rect 9447 49371 9533 49427
rect 9589 49371 9675 49427
rect 9731 49371 9817 49427
rect 9873 49371 9959 49427
rect 10015 49371 10101 49427
rect 10157 49371 10243 49427
rect 10299 49371 10385 49427
rect 10441 49371 10527 49427
rect 10583 49371 10669 49427
rect 10725 49371 10811 49427
rect 10867 49371 10953 49427
rect 11009 49371 11095 49427
rect 11151 49371 11237 49427
rect 11293 49371 11379 49427
rect 11435 49371 11521 49427
rect 11577 49371 11663 49427
rect 11719 49371 11805 49427
rect 11861 49371 11947 49427
rect 12003 49371 12089 49427
rect 12145 49371 12231 49427
rect 12287 49371 12373 49427
rect 12429 49371 12515 49427
rect 12571 49371 12657 49427
rect 12713 49371 12799 49427
rect 12855 49371 12941 49427
rect 12997 49371 13083 49427
rect 13139 49371 13225 49427
rect 13281 49371 13367 49427
rect 13423 49371 13509 49427
rect 13565 49371 13651 49427
rect 13707 49371 13793 49427
rect 13849 49371 13935 49427
rect 13991 49371 14077 49427
rect 14133 49371 14219 49427
rect 14275 49371 14361 49427
rect 14417 49371 14503 49427
rect 14559 49371 14645 49427
rect 14701 49371 14787 49427
rect 14843 49371 14853 49427
rect 151 49285 14853 49371
rect 151 49229 161 49285
rect 217 49229 303 49285
rect 359 49229 445 49285
rect 501 49229 587 49285
rect 643 49229 729 49285
rect 785 49229 871 49285
rect 927 49229 1013 49285
rect 1069 49229 1155 49285
rect 1211 49229 1297 49285
rect 1353 49229 1439 49285
rect 1495 49229 1581 49285
rect 1637 49229 1723 49285
rect 1779 49229 1865 49285
rect 1921 49229 2007 49285
rect 2063 49229 2149 49285
rect 2205 49229 2291 49285
rect 2347 49229 2433 49285
rect 2489 49229 2575 49285
rect 2631 49229 2717 49285
rect 2773 49229 2859 49285
rect 2915 49229 3001 49285
rect 3057 49229 3143 49285
rect 3199 49229 3285 49285
rect 3341 49229 3427 49285
rect 3483 49229 3569 49285
rect 3625 49229 3711 49285
rect 3767 49229 3853 49285
rect 3909 49229 3995 49285
rect 4051 49229 4137 49285
rect 4193 49229 4279 49285
rect 4335 49229 4421 49285
rect 4477 49229 4563 49285
rect 4619 49229 4705 49285
rect 4761 49229 4847 49285
rect 4903 49229 4989 49285
rect 5045 49229 5131 49285
rect 5187 49229 5273 49285
rect 5329 49229 5415 49285
rect 5471 49229 5557 49285
rect 5613 49229 5699 49285
rect 5755 49229 5841 49285
rect 5897 49229 5983 49285
rect 6039 49229 6125 49285
rect 6181 49229 6267 49285
rect 6323 49229 6409 49285
rect 6465 49229 6551 49285
rect 6607 49229 6693 49285
rect 6749 49229 6835 49285
rect 6891 49229 6977 49285
rect 7033 49229 7119 49285
rect 7175 49229 7261 49285
rect 7317 49229 7403 49285
rect 7459 49229 7545 49285
rect 7601 49229 7687 49285
rect 7743 49229 7829 49285
rect 7885 49229 7971 49285
rect 8027 49229 8113 49285
rect 8169 49229 8255 49285
rect 8311 49229 8397 49285
rect 8453 49229 8539 49285
rect 8595 49229 8681 49285
rect 8737 49229 8823 49285
rect 8879 49229 8965 49285
rect 9021 49229 9107 49285
rect 9163 49229 9249 49285
rect 9305 49229 9391 49285
rect 9447 49229 9533 49285
rect 9589 49229 9675 49285
rect 9731 49229 9817 49285
rect 9873 49229 9959 49285
rect 10015 49229 10101 49285
rect 10157 49229 10243 49285
rect 10299 49229 10385 49285
rect 10441 49229 10527 49285
rect 10583 49229 10669 49285
rect 10725 49229 10811 49285
rect 10867 49229 10953 49285
rect 11009 49229 11095 49285
rect 11151 49229 11237 49285
rect 11293 49229 11379 49285
rect 11435 49229 11521 49285
rect 11577 49229 11663 49285
rect 11719 49229 11805 49285
rect 11861 49229 11947 49285
rect 12003 49229 12089 49285
rect 12145 49229 12231 49285
rect 12287 49229 12373 49285
rect 12429 49229 12515 49285
rect 12571 49229 12657 49285
rect 12713 49229 12799 49285
rect 12855 49229 12941 49285
rect 12997 49229 13083 49285
rect 13139 49229 13225 49285
rect 13281 49229 13367 49285
rect 13423 49229 13509 49285
rect 13565 49229 13651 49285
rect 13707 49229 13793 49285
rect 13849 49229 13935 49285
rect 13991 49229 14077 49285
rect 14133 49229 14219 49285
rect 14275 49229 14361 49285
rect 14417 49229 14503 49285
rect 14559 49229 14645 49285
rect 14701 49229 14787 49285
rect 14843 49229 14853 49285
rect 151 49219 14853 49229
rect 151 48941 14853 48951
rect 151 48885 161 48941
rect 217 48885 303 48941
rect 359 48885 445 48941
rect 501 48885 587 48941
rect 643 48885 729 48941
rect 785 48885 871 48941
rect 927 48885 1013 48941
rect 1069 48885 1155 48941
rect 1211 48885 1297 48941
rect 1353 48885 1439 48941
rect 1495 48885 1581 48941
rect 1637 48885 1723 48941
rect 1779 48885 1865 48941
rect 1921 48885 2007 48941
rect 2063 48885 2149 48941
rect 2205 48885 2291 48941
rect 2347 48885 2433 48941
rect 2489 48885 2575 48941
rect 2631 48885 2717 48941
rect 2773 48885 2859 48941
rect 2915 48885 3001 48941
rect 3057 48885 3143 48941
rect 3199 48885 3285 48941
rect 3341 48885 3427 48941
rect 3483 48885 3569 48941
rect 3625 48885 3711 48941
rect 3767 48885 3853 48941
rect 3909 48885 3995 48941
rect 4051 48885 4137 48941
rect 4193 48885 4279 48941
rect 4335 48885 4421 48941
rect 4477 48885 4563 48941
rect 4619 48885 4705 48941
rect 4761 48885 4847 48941
rect 4903 48885 4989 48941
rect 5045 48885 5131 48941
rect 5187 48885 5273 48941
rect 5329 48885 5415 48941
rect 5471 48885 5557 48941
rect 5613 48885 5699 48941
rect 5755 48885 5841 48941
rect 5897 48885 5983 48941
rect 6039 48885 6125 48941
rect 6181 48885 6267 48941
rect 6323 48885 6409 48941
rect 6465 48885 6551 48941
rect 6607 48885 6693 48941
rect 6749 48885 6835 48941
rect 6891 48885 6977 48941
rect 7033 48885 7119 48941
rect 7175 48885 7261 48941
rect 7317 48885 7403 48941
rect 7459 48885 7545 48941
rect 7601 48885 7687 48941
rect 7743 48885 7829 48941
rect 7885 48885 7971 48941
rect 8027 48885 8113 48941
rect 8169 48885 8255 48941
rect 8311 48885 8397 48941
rect 8453 48885 8539 48941
rect 8595 48885 8681 48941
rect 8737 48885 8823 48941
rect 8879 48885 8965 48941
rect 9021 48885 9107 48941
rect 9163 48885 9249 48941
rect 9305 48885 9391 48941
rect 9447 48885 9533 48941
rect 9589 48885 9675 48941
rect 9731 48885 9817 48941
rect 9873 48885 9959 48941
rect 10015 48885 10101 48941
rect 10157 48885 10243 48941
rect 10299 48885 10385 48941
rect 10441 48885 10527 48941
rect 10583 48885 10669 48941
rect 10725 48885 10811 48941
rect 10867 48885 10953 48941
rect 11009 48885 11095 48941
rect 11151 48885 11237 48941
rect 11293 48885 11379 48941
rect 11435 48885 11521 48941
rect 11577 48885 11663 48941
rect 11719 48885 11805 48941
rect 11861 48885 11947 48941
rect 12003 48885 12089 48941
rect 12145 48885 12231 48941
rect 12287 48885 12373 48941
rect 12429 48885 12515 48941
rect 12571 48885 12657 48941
rect 12713 48885 12799 48941
rect 12855 48885 12941 48941
rect 12997 48885 13083 48941
rect 13139 48885 13225 48941
rect 13281 48885 13367 48941
rect 13423 48885 13509 48941
rect 13565 48885 13651 48941
rect 13707 48885 13793 48941
rect 13849 48885 13935 48941
rect 13991 48885 14077 48941
rect 14133 48885 14219 48941
rect 14275 48885 14361 48941
rect 14417 48885 14503 48941
rect 14559 48885 14645 48941
rect 14701 48885 14787 48941
rect 14843 48885 14853 48941
rect 151 48799 14853 48885
rect 151 48743 161 48799
rect 217 48743 303 48799
rect 359 48743 445 48799
rect 501 48743 587 48799
rect 643 48743 729 48799
rect 785 48743 871 48799
rect 927 48743 1013 48799
rect 1069 48743 1155 48799
rect 1211 48743 1297 48799
rect 1353 48743 1439 48799
rect 1495 48743 1581 48799
rect 1637 48743 1723 48799
rect 1779 48743 1865 48799
rect 1921 48743 2007 48799
rect 2063 48743 2149 48799
rect 2205 48743 2291 48799
rect 2347 48743 2433 48799
rect 2489 48743 2575 48799
rect 2631 48743 2717 48799
rect 2773 48743 2859 48799
rect 2915 48743 3001 48799
rect 3057 48743 3143 48799
rect 3199 48743 3285 48799
rect 3341 48743 3427 48799
rect 3483 48743 3569 48799
rect 3625 48743 3711 48799
rect 3767 48743 3853 48799
rect 3909 48743 3995 48799
rect 4051 48743 4137 48799
rect 4193 48743 4279 48799
rect 4335 48743 4421 48799
rect 4477 48743 4563 48799
rect 4619 48743 4705 48799
rect 4761 48743 4847 48799
rect 4903 48743 4989 48799
rect 5045 48743 5131 48799
rect 5187 48743 5273 48799
rect 5329 48743 5415 48799
rect 5471 48743 5557 48799
rect 5613 48743 5699 48799
rect 5755 48743 5841 48799
rect 5897 48743 5983 48799
rect 6039 48743 6125 48799
rect 6181 48743 6267 48799
rect 6323 48743 6409 48799
rect 6465 48743 6551 48799
rect 6607 48743 6693 48799
rect 6749 48743 6835 48799
rect 6891 48743 6977 48799
rect 7033 48743 7119 48799
rect 7175 48743 7261 48799
rect 7317 48743 7403 48799
rect 7459 48743 7545 48799
rect 7601 48743 7687 48799
rect 7743 48743 7829 48799
rect 7885 48743 7971 48799
rect 8027 48743 8113 48799
rect 8169 48743 8255 48799
rect 8311 48743 8397 48799
rect 8453 48743 8539 48799
rect 8595 48743 8681 48799
rect 8737 48743 8823 48799
rect 8879 48743 8965 48799
rect 9021 48743 9107 48799
rect 9163 48743 9249 48799
rect 9305 48743 9391 48799
rect 9447 48743 9533 48799
rect 9589 48743 9675 48799
rect 9731 48743 9817 48799
rect 9873 48743 9959 48799
rect 10015 48743 10101 48799
rect 10157 48743 10243 48799
rect 10299 48743 10385 48799
rect 10441 48743 10527 48799
rect 10583 48743 10669 48799
rect 10725 48743 10811 48799
rect 10867 48743 10953 48799
rect 11009 48743 11095 48799
rect 11151 48743 11237 48799
rect 11293 48743 11379 48799
rect 11435 48743 11521 48799
rect 11577 48743 11663 48799
rect 11719 48743 11805 48799
rect 11861 48743 11947 48799
rect 12003 48743 12089 48799
rect 12145 48743 12231 48799
rect 12287 48743 12373 48799
rect 12429 48743 12515 48799
rect 12571 48743 12657 48799
rect 12713 48743 12799 48799
rect 12855 48743 12941 48799
rect 12997 48743 13083 48799
rect 13139 48743 13225 48799
rect 13281 48743 13367 48799
rect 13423 48743 13509 48799
rect 13565 48743 13651 48799
rect 13707 48743 13793 48799
rect 13849 48743 13935 48799
rect 13991 48743 14077 48799
rect 14133 48743 14219 48799
rect 14275 48743 14361 48799
rect 14417 48743 14503 48799
rect 14559 48743 14645 48799
rect 14701 48743 14787 48799
rect 14843 48743 14853 48799
rect 151 48657 14853 48743
rect 151 48601 161 48657
rect 217 48601 303 48657
rect 359 48601 445 48657
rect 501 48601 587 48657
rect 643 48601 729 48657
rect 785 48601 871 48657
rect 927 48601 1013 48657
rect 1069 48601 1155 48657
rect 1211 48601 1297 48657
rect 1353 48601 1439 48657
rect 1495 48601 1581 48657
rect 1637 48601 1723 48657
rect 1779 48601 1865 48657
rect 1921 48601 2007 48657
rect 2063 48601 2149 48657
rect 2205 48601 2291 48657
rect 2347 48601 2433 48657
rect 2489 48601 2575 48657
rect 2631 48601 2717 48657
rect 2773 48601 2859 48657
rect 2915 48601 3001 48657
rect 3057 48601 3143 48657
rect 3199 48601 3285 48657
rect 3341 48601 3427 48657
rect 3483 48601 3569 48657
rect 3625 48601 3711 48657
rect 3767 48601 3853 48657
rect 3909 48601 3995 48657
rect 4051 48601 4137 48657
rect 4193 48601 4279 48657
rect 4335 48601 4421 48657
rect 4477 48601 4563 48657
rect 4619 48601 4705 48657
rect 4761 48601 4847 48657
rect 4903 48601 4989 48657
rect 5045 48601 5131 48657
rect 5187 48601 5273 48657
rect 5329 48601 5415 48657
rect 5471 48601 5557 48657
rect 5613 48601 5699 48657
rect 5755 48601 5841 48657
rect 5897 48601 5983 48657
rect 6039 48601 6125 48657
rect 6181 48601 6267 48657
rect 6323 48601 6409 48657
rect 6465 48601 6551 48657
rect 6607 48601 6693 48657
rect 6749 48601 6835 48657
rect 6891 48601 6977 48657
rect 7033 48601 7119 48657
rect 7175 48601 7261 48657
rect 7317 48601 7403 48657
rect 7459 48601 7545 48657
rect 7601 48601 7687 48657
rect 7743 48601 7829 48657
rect 7885 48601 7971 48657
rect 8027 48601 8113 48657
rect 8169 48601 8255 48657
rect 8311 48601 8397 48657
rect 8453 48601 8539 48657
rect 8595 48601 8681 48657
rect 8737 48601 8823 48657
rect 8879 48601 8965 48657
rect 9021 48601 9107 48657
rect 9163 48601 9249 48657
rect 9305 48601 9391 48657
rect 9447 48601 9533 48657
rect 9589 48601 9675 48657
rect 9731 48601 9817 48657
rect 9873 48601 9959 48657
rect 10015 48601 10101 48657
rect 10157 48601 10243 48657
rect 10299 48601 10385 48657
rect 10441 48601 10527 48657
rect 10583 48601 10669 48657
rect 10725 48601 10811 48657
rect 10867 48601 10953 48657
rect 11009 48601 11095 48657
rect 11151 48601 11237 48657
rect 11293 48601 11379 48657
rect 11435 48601 11521 48657
rect 11577 48601 11663 48657
rect 11719 48601 11805 48657
rect 11861 48601 11947 48657
rect 12003 48601 12089 48657
rect 12145 48601 12231 48657
rect 12287 48601 12373 48657
rect 12429 48601 12515 48657
rect 12571 48601 12657 48657
rect 12713 48601 12799 48657
rect 12855 48601 12941 48657
rect 12997 48601 13083 48657
rect 13139 48601 13225 48657
rect 13281 48601 13367 48657
rect 13423 48601 13509 48657
rect 13565 48601 13651 48657
rect 13707 48601 13793 48657
rect 13849 48601 13935 48657
rect 13991 48601 14077 48657
rect 14133 48601 14219 48657
rect 14275 48601 14361 48657
rect 14417 48601 14503 48657
rect 14559 48601 14645 48657
rect 14701 48601 14787 48657
rect 14843 48601 14853 48657
rect 151 48515 14853 48601
rect 151 48459 161 48515
rect 217 48459 303 48515
rect 359 48459 445 48515
rect 501 48459 587 48515
rect 643 48459 729 48515
rect 785 48459 871 48515
rect 927 48459 1013 48515
rect 1069 48459 1155 48515
rect 1211 48459 1297 48515
rect 1353 48459 1439 48515
rect 1495 48459 1581 48515
rect 1637 48459 1723 48515
rect 1779 48459 1865 48515
rect 1921 48459 2007 48515
rect 2063 48459 2149 48515
rect 2205 48459 2291 48515
rect 2347 48459 2433 48515
rect 2489 48459 2575 48515
rect 2631 48459 2717 48515
rect 2773 48459 2859 48515
rect 2915 48459 3001 48515
rect 3057 48459 3143 48515
rect 3199 48459 3285 48515
rect 3341 48459 3427 48515
rect 3483 48459 3569 48515
rect 3625 48459 3711 48515
rect 3767 48459 3853 48515
rect 3909 48459 3995 48515
rect 4051 48459 4137 48515
rect 4193 48459 4279 48515
rect 4335 48459 4421 48515
rect 4477 48459 4563 48515
rect 4619 48459 4705 48515
rect 4761 48459 4847 48515
rect 4903 48459 4989 48515
rect 5045 48459 5131 48515
rect 5187 48459 5273 48515
rect 5329 48459 5415 48515
rect 5471 48459 5557 48515
rect 5613 48459 5699 48515
rect 5755 48459 5841 48515
rect 5897 48459 5983 48515
rect 6039 48459 6125 48515
rect 6181 48459 6267 48515
rect 6323 48459 6409 48515
rect 6465 48459 6551 48515
rect 6607 48459 6693 48515
rect 6749 48459 6835 48515
rect 6891 48459 6977 48515
rect 7033 48459 7119 48515
rect 7175 48459 7261 48515
rect 7317 48459 7403 48515
rect 7459 48459 7545 48515
rect 7601 48459 7687 48515
rect 7743 48459 7829 48515
rect 7885 48459 7971 48515
rect 8027 48459 8113 48515
rect 8169 48459 8255 48515
rect 8311 48459 8397 48515
rect 8453 48459 8539 48515
rect 8595 48459 8681 48515
rect 8737 48459 8823 48515
rect 8879 48459 8965 48515
rect 9021 48459 9107 48515
rect 9163 48459 9249 48515
rect 9305 48459 9391 48515
rect 9447 48459 9533 48515
rect 9589 48459 9675 48515
rect 9731 48459 9817 48515
rect 9873 48459 9959 48515
rect 10015 48459 10101 48515
rect 10157 48459 10243 48515
rect 10299 48459 10385 48515
rect 10441 48459 10527 48515
rect 10583 48459 10669 48515
rect 10725 48459 10811 48515
rect 10867 48459 10953 48515
rect 11009 48459 11095 48515
rect 11151 48459 11237 48515
rect 11293 48459 11379 48515
rect 11435 48459 11521 48515
rect 11577 48459 11663 48515
rect 11719 48459 11805 48515
rect 11861 48459 11947 48515
rect 12003 48459 12089 48515
rect 12145 48459 12231 48515
rect 12287 48459 12373 48515
rect 12429 48459 12515 48515
rect 12571 48459 12657 48515
rect 12713 48459 12799 48515
rect 12855 48459 12941 48515
rect 12997 48459 13083 48515
rect 13139 48459 13225 48515
rect 13281 48459 13367 48515
rect 13423 48459 13509 48515
rect 13565 48459 13651 48515
rect 13707 48459 13793 48515
rect 13849 48459 13935 48515
rect 13991 48459 14077 48515
rect 14133 48459 14219 48515
rect 14275 48459 14361 48515
rect 14417 48459 14503 48515
rect 14559 48459 14645 48515
rect 14701 48459 14787 48515
rect 14843 48459 14853 48515
rect 151 48373 14853 48459
rect 151 48317 161 48373
rect 217 48317 303 48373
rect 359 48317 445 48373
rect 501 48317 587 48373
rect 643 48317 729 48373
rect 785 48317 871 48373
rect 927 48317 1013 48373
rect 1069 48317 1155 48373
rect 1211 48317 1297 48373
rect 1353 48317 1439 48373
rect 1495 48317 1581 48373
rect 1637 48317 1723 48373
rect 1779 48317 1865 48373
rect 1921 48317 2007 48373
rect 2063 48317 2149 48373
rect 2205 48317 2291 48373
rect 2347 48317 2433 48373
rect 2489 48317 2575 48373
rect 2631 48317 2717 48373
rect 2773 48317 2859 48373
rect 2915 48317 3001 48373
rect 3057 48317 3143 48373
rect 3199 48317 3285 48373
rect 3341 48317 3427 48373
rect 3483 48317 3569 48373
rect 3625 48317 3711 48373
rect 3767 48317 3853 48373
rect 3909 48317 3995 48373
rect 4051 48317 4137 48373
rect 4193 48317 4279 48373
rect 4335 48317 4421 48373
rect 4477 48317 4563 48373
rect 4619 48317 4705 48373
rect 4761 48317 4847 48373
rect 4903 48317 4989 48373
rect 5045 48317 5131 48373
rect 5187 48317 5273 48373
rect 5329 48317 5415 48373
rect 5471 48317 5557 48373
rect 5613 48317 5699 48373
rect 5755 48317 5841 48373
rect 5897 48317 5983 48373
rect 6039 48317 6125 48373
rect 6181 48317 6267 48373
rect 6323 48317 6409 48373
rect 6465 48317 6551 48373
rect 6607 48317 6693 48373
rect 6749 48317 6835 48373
rect 6891 48317 6977 48373
rect 7033 48317 7119 48373
rect 7175 48317 7261 48373
rect 7317 48317 7403 48373
rect 7459 48317 7545 48373
rect 7601 48317 7687 48373
rect 7743 48317 7829 48373
rect 7885 48317 7971 48373
rect 8027 48317 8113 48373
rect 8169 48317 8255 48373
rect 8311 48317 8397 48373
rect 8453 48317 8539 48373
rect 8595 48317 8681 48373
rect 8737 48317 8823 48373
rect 8879 48317 8965 48373
rect 9021 48317 9107 48373
rect 9163 48317 9249 48373
rect 9305 48317 9391 48373
rect 9447 48317 9533 48373
rect 9589 48317 9675 48373
rect 9731 48317 9817 48373
rect 9873 48317 9959 48373
rect 10015 48317 10101 48373
rect 10157 48317 10243 48373
rect 10299 48317 10385 48373
rect 10441 48317 10527 48373
rect 10583 48317 10669 48373
rect 10725 48317 10811 48373
rect 10867 48317 10953 48373
rect 11009 48317 11095 48373
rect 11151 48317 11237 48373
rect 11293 48317 11379 48373
rect 11435 48317 11521 48373
rect 11577 48317 11663 48373
rect 11719 48317 11805 48373
rect 11861 48317 11947 48373
rect 12003 48317 12089 48373
rect 12145 48317 12231 48373
rect 12287 48317 12373 48373
rect 12429 48317 12515 48373
rect 12571 48317 12657 48373
rect 12713 48317 12799 48373
rect 12855 48317 12941 48373
rect 12997 48317 13083 48373
rect 13139 48317 13225 48373
rect 13281 48317 13367 48373
rect 13423 48317 13509 48373
rect 13565 48317 13651 48373
rect 13707 48317 13793 48373
rect 13849 48317 13935 48373
rect 13991 48317 14077 48373
rect 14133 48317 14219 48373
rect 14275 48317 14361 48373
rect 14417 48317 14503 48373
rect 14559 48317 14645 48373
rect 14701 48317 14787 48373
rect 14843 48317 14853 48373
rect 151 48231 14853 48317
rect 151 48175 161 48231
rect 217 48175 303 48231
rect 359 48175 445 48231
rect 501 48175 587 48231
rect 643 48175 729 48231
rect 785 48175 871 48231
rect 927 48175 1013 48231
rect 1069 48175 1155 48231
rect 1211 48175 1297 48231
rect 1353 48175 1439 48231
rect 1495 48175 1581 48231
rect 1637 48175 1723 48231
rect 1779 48175 1865 48231
rect 1921 48175 2007 48231
rect 2063 48175 2149 48231
rect 2205 48175 2291 48231
rect 2347 48175 2433 48231
rect 2489 48175 2575 48231
rect 2631 48175 2717 48231
rect 2773 48175 2859 48231
rect 2915 48175 3001 48231
rect 3057 48175 3143 48231
rect 3199 48175 3285 48231
rect 3341 48175 3427 48231
rect 3483 48175 3569 48231
rect 3625 48175 3711 48231
rect 3767 48175 3853 48231
rect 3909 48175 3995 48231
rect 4051 48175 4137 48231
rect 4193 48175 4279 48231
rect 4335 48175 4421 48231
rect 4477 48175 4563 48231
rect 4619 48175 4705 48231
rect 4761 48175 4847 48231
rect 4903 48175 4989 48231
rect 5045 48175 5131 48231
rect 5187 48175 5273 48231
rect 5329 48175 5415 48231
rect 5471 48175 5557 48231
rect 5613 48175 5699 48231
rect 5755 48175 5841 48231
rect 5897 48175 5983 48231
rect 6039 48175 6125 48231
rect 6181 48175 6267 48231
rect 6323 48175 6409 48231
rect 6465 48175 6551 48231
rect 6607 48175 6693 48231
rect 6749 48175 6835 48231
rect 6891 48175 6977 48231
rect 7033 48175 7119 48231
rect 7175 48175 7261 48231
rect 7317 48175 7403 48231
rect 7459 48175 7545 48231
rect 7601 48175 7687 48231
rect 7743 48175 7829 48231
rect 7885 48175 7971 48231
rect 8027 48175 8113 48231
rect 8169 48175 8255 48231
rect 8311 48175 8397 48231
rect 8453 48175 8539 48231
rect 8595 48175 8681 48231
rect 8737 48175 8823 48231
rect 8879 48175 8965 48231
rect 9021 48175 9107 48231
rect 9163 48175 9249 48231
rect 9305 48175 9391 48231
rect 9447 48175 9533 48231
rect 9589 48175 9675 48231
rect 9731 48175 9817 48231
rect 9873 48175 9959 48231
rect 10015 48175 10101 48231
rect 10157 48175 10243 48231
rect 10299 48175 10385 48231
rect 10441 48175 10527 48231
rect 10583 48175 10669 48231
rect 10725 48175 10811 48231
rect 10867 48175 10953 48231
rect 11009 48175 11095 48231
rect 11151 48175 11237 48231
rect 11293 48175 11379 48231
rect 11435 48175 11521 48231
rect 11577 48175 11663 48231
rect 11719 48175 11805 48231
rect 11861 48175 11947 48231
rect 12003 48175 12089 48231
rect 12145 48175 12231 48231
rect 12287 48175 12373 48231
rect 12429 48175 12515 48231
rect 12571 48175 12657 48231
rect 12713 48175 12799 48231
rect 12855 48175 12941 48231
rect 12997 48175 13083 48231
rect 13139 48175 13225 48231
rect 13281 48175 13367 48231
rect 13423 48175 13509 48231
rect 13565 48175 13651 48231
rect 13707 48175 13793 48231
rect 13849 48175 13935 48231
rect 13991 48175 14077 48231
rect 14133 48175 14219 48231
rect 14275 48175 14361 48231
rect 14417 48175 14503 48231
rect 14559 48175 14645 48231
rect 14701 48175 14787 48231
rect 14843 48175 14853 48231
rect 151 48089 14853 48175
rect 151 48033 161 48089
rect 217 48033 303 48089
rect 359 48033 445 48089
rect 501 48033 587 48089
rect 643 48033 729 48089
rect 785 48033 871 48089
rect 927 48033 1013 48089
rect 1069 48033 1155 48089
rect 1211 48033 1297 48089
rect 1353 48033 1439 48089
rect 1495 48033 1581 48089
rect 1637 48033 1723 48089
rect 1779 48033 1865 48089
rect 1921 48033 2007 48089
rect 2063 48033 2149 48089
rect 2205 48033 2291 48089
rect 2347 48033 2433 48089
rect 2489 48033 2575 48089
rect 2631 48033 2717 48089
rect 2773 48033 2859 48089
rect 2915 48033 3001 48089
rect 3057 48033 3143 48089
rect 3199 48033 3285 48089
rect 3341 48033 3427 48089
rect 3483 48033 3569 48089
rect 3625 48033 3711 48089
rect 3767 48033 3853 48089
rect 3909 48033 3995 48089
rect 4051 48033 4137 48089
rect 4193 48033 4279 48089
rect 4335 48033 4421 48089
rect 4477 48033 4563 48089
rect 4619 48033 4705 48089
rect 4761 48033 4847 48089
rect 4903 48033 4989 48089
rect 5045 48033 5131 48089
rect 5187 48033 5273 48089
rect 5329 48033 5415 48089
rect 5471 48033 5557 48089
rect 5613 48033 5699 48089
rect 5755 48033 5841 48089
rect 5897 48033 5983 48089
rect 6039 48033 6125 48089
rect 6181 48033 6267 48089
rect 6323 48033 6409 48089
rect 6465 48033 6551 48089
rect 6607 48033 6693 48089
rect 6749 48033 6835 48089
rect 6891 48033 6977 48089
rect 7033 48033 7119 48089
rect 7175 48033 7261 48089
rect 7317 48033 7403 48089
rect 7459 48033 7545 48089
rect 7601 48033 7687 48089
rect 7743 48033 7829 48089
rect 7885 48033 7971 48089
rect 8027 48033 8113 48089
rect 8169 48033 8255 48089
rect 8311 48033 8397 48089
rect 8453 48033 8539 48089
rect 8595 48033 8681 48089
rect 8737 48033 8823 48089
rect 8879 48033 8965 48089
rect 9021 48033 9107 48089
rect 9163 48033 9249 48089
rect 9305 48033 9391 48089
rect 9447 48033 9533 48089
rect 9589 48033 9675 48089
rect 9731 48033 9817 48089
rect 9873 48033 9959 48089
rect 10015 48033 10101 48089
rect 10157 48033 10243 48089
rect 10299 48033 10385 48089
rect 10441 48033 10527 48089
rect 10583 48033 10669 48089
rect 10725 48033 10811 48089
rect 10867 48033 10953 48089
rect 11009 48033 11095 48089
rect 11151 48033 11237 48089
rect 11293 48033 11379 48089
rect 11435 48033 11521 48089
rect 11577 48033 11663 48089
rect 11719 48033 11805 48089
rect 11861 48033 11947 48089
rect 12003 48033 12089 48089
rect 12145 48033 12231 48089
rect 12287 48033 12373 48089
rect 12429 48033 12515 48089
rect 12571 48033 12657 48089
rect 12713 48033 12799 48089
rect 12855 48033 12941 48089
rect 12997 48033 13083 48089
rect 13139 48033 13225 48089
rect 13281 48033 13367 48089
rect 13423 48033 13509 48089
rect 13565 48033 13651 48089
rect 13707 48033 13793 48089
rect 13849 48033 13935 48089
rect 13991 48033 14077 48089
rect 14133 48033 14219 48089
rect 14275 48033 14361 48089
rect 14417 48033 14503 48089
rect 14559 48033 14645 48089
rect 14701 48033 14787 48089
rect 14843 48033 14853 48089
rect 151 47947 14853 48033
rect 151 47891 161 47947
rect 217 47891 303 47947
rect 359 47891 445 47947
rect 501 47891 587 47947
rect 643 47891 729 47947
rect 785 47891 871 47947
rect 927 47891 1013 47947
rect 1069 47891 1155 47947
rect 1211 47891 1297 47947
rect 1353 47891 1439 47947
rect 1495 47891 1581 47947
rect 1637 47891 1723 47947
rect 1779 47891 1865 47947
rect 1921 47891 2007 47947
rect 2063 47891 2149 47947
rect 2205 47891 2291 47947
rect 2347 47891 2433 47947
rect 2489 47891 2575 47947
rect 2631 47891 2717 47947
rect 2773 47891 2859 47947
rect 2915 47891 3001 47947
rect 3057 47891 3143 47947
rect 3199 47891 3285 47947
rect 3341 47891 3427 47947
rect 3483 47891 3569 47947
rect 3625 47891 3711 47947
rect 3767 47891 3853 47947
rect 3909 47891 3995 47947
rect 4051 47891 4137 47947
rect 4193 47891 4279 47947
rect 4335 47891 4421 47947
rect 4477 47891 4563 47947
rect 4619 47891 4705 47947
rect 4761 47891 4847 47947
rect 4903 47891 4989 47947
rect 5045 47891 5131 47947
rect 5187 47891 5273 47947
rect 5329 47891 5415 47947
rect 5471 47891 5557 47947
rect 5613 47891 5699 47947
rect 5755 47891 5841 47947
rect 5897 47891 5983 47947
rect 6039 47891 6125 47947
rect 6181 47891 6267 47947
rect 6323 47891 6409 47947
rect 6465 47891 6551 47947
rect 6607 47891 6693 47947
rect 6749 47891 6835 47947
rect 6891 47891 6977 47947
rect 7033 47891 7119 47947
rect 7175 47891 7261 47947
rect 7317 47891 7403 47947
rect 7459 47891 7545 47947
rect 7601 47891 7687 47947
rect 7743 47891 7829 47947
rect 7885 47891 7971 47947
rect 8027 47891 8113 47947
rect 8169 47891 8255 47947
rect 8311 47891 8397 47947
rect 8453 47891 8539 47947
rect 8595 47891 8681 47947
rect 8737 47891 8823 47947
rect 8879 47891 8965 47947
rect 9021 47891 9107 47947
rect 9163 47891 9249 47947
rect 9305 47891 9391 47947
rect 9447 47891 9533 47947
rect 9589 47891 9675 47947
rect 9731 47891 9817 47947
rect 9873 47891 9959 47947
rect 10015 47891 10101 47947
rect 10157 47891 10243 47947
rect 10299 47891 10385 47947
rect 10441 47891 10527 47947
rect 10583 47891 10669 47947
rect 10725 47891 10811 47947
rect 10867 47891 10953 47947
rect 11009 47891 11095 47947
rect 11151 47891 11237 47947
rect 11293 47891 11379 47947
rect 11435 47891 11521 47947
rect 11577 47891 11663 47947
rect 11719 47891 11805 47947
rect 11861 47891 11947 47947
rect 12003 47891 12089 47947
rect 12145 47891 12231 47947
rect 12287 47891 12373 47947
rect 12429 47891 12515 47947
rect 12571 47891 12657 47947
rect 12713 47891 12799 47947
rect 12855 47891 12941 47947
rect 12997 47891 13083 47947
rect 13139 47891 13225 47947
rect 13281 47891 13367 47947
rect 13423 47891 13509 47947
rect 13565 47891 13651 47947
rect 13707 47891 13793 47947
rect 13849 47891 13935 47947
rect 13991 47891 14077 47947
rect 14133 47891 14219 47947
rect 14275 47891 14361 47947
rect 14417 47891 14503 47947
rect 14559 47891 14645 47947
rect 14701 47891 14787 47947
rect 14843 47891 14853 47947
rect 151 47805 14853 47891
rect 151 47749 161 47805
rect 217 47749 303 47805
rect 359 47749 445 47805
rect 501 47749 587 47805
rect 643 47749 729 47805
rect 785 47749 871 47805
rect 927 47749 1013 47805
rect 1069 47749 1155 47805
rect 1211 47749 1297 47805
rect 1353 47749 1439 47805
rect 1495 47749 1581 47805
rect 1637 47749 1723 47805
rect 1779 47749 1865 47805
rect 1921 47749 2007 47805
rect 2063 47749 2149 47805
rect 2205 47749 2291 47805
rect 2347 47749 2433 47805
rect 2489 47749 2575 47805
rect 2631 47749 2717 47805
rect 2773 47749 2859 47805
rect 2915 47749 3001 47805
rect 3057 47749 3143 47805
rect 3199 47749 3285 47805
rect 3341 47749 3427 47805
rect 3483 47749 3569 47805
rect 3625 47749 3711 47805
rect 3767 47749 3853 47805
rect 3909 47749 3995 47805
rect 4051 47749 4137 47805
rect 4193 47749 4279 47805
rect 4335 47749 4421 47805
rect 4477 47749 4563 47805
rect 4619 47749 4705 47805
rect 4761 47749 4847 47805
rect 4903 47749 4989 47805
rect 5045 47749 5131 47805
rect 5187 47749 5273 47805
rect 5329 47749 5415 47805
rect 5471 47749 5557 47805
rect 5613 47749 5699 47805
rect 5755 47749 5841 47805
rect 5897 47749 5983 47805
rect 6039 47749 6125 47805
rect 6181 47749 6267 47805
rect 6323 47749 6409 47805
rect 6465 47749 6551 47805
rect 6607 47749 6693 47805
rect 6749 47749 6835 47805
rect 6891 47749 6977 47805
rect 7033 47749 7119 47805
rect 7175 47749 7261 47805
rect 7317 47749 7403 47805
rect 7459 47749 7545 47805
rect 7601 47749 7687 47805
rect 7743 47749 7829 47805
rect 7885 47749 7971 47805
rect 8027 47749 8113 47805
rect 8169 47749 8255 47805
rect 8311 47749 8397 47805
rect 8453 47749 8539 47805
rect 8595 47749 8681 47805
rect 8737 47749 8823 47805
rect 8879 47749 8965 47805
rect 9021 47749 9107 47805
rect 9163 47749 9249 47805
rect 9305 47749 9391 47805
rect 9447 47749 9533 47805
rect 9589 47749 9675 47805
rect 9731 47749 9817 47805
rect 9873 47749 9959 47805
rect 10015 47749 10101 47805
rect 10157 47749 10243 47805
rect 10299 47749 10385 47805
rect 10441 47749 10527 47805
rect 10583 47749 10669 47805
rect 10725 47749 10811 47805
rect 10867 47749 10953 47805
rect 11009 47749 11095 47805
rect 11151 47749 11237 47805
rect 11293 47749 11379 47805
rect 11435 47749 11521 47805
rect 11577 47749 11663 47805
rect 11719 47749 11805 47805
rect 11861 47749 11947 47805
rect 12003 47749 12089 47805
rect 12145 47749 12231 47805
rect 12287 47749 12373 47805
rect 12429 47749 12515 47805
rect 12571 47749 12657 47805
rect 12713 47749 12799 47805
rect 12855 47749 12941 47805
rect 12997 47749 13083 47805
rect 13139 47749 13225 47805
rect 13281 47749 13367 47805
rect 13423 47749 13509 47805
rect 13565 47749 13651 47805
rect 13707 47749 13793 47805
rect 13849 47749 13935 47805
rect 13991 47749 14077 47805
rect 14133 47749 14219 47805
rect 14275 47749 14361 47805
rect 14417 47749 14503 47805
rect 14559 47749 14645 47805
rect 14701 47749 14787 47805
rect 14843 47749 14853 47805
rect 151 47663 14853 47749
rect 151 47607 161 47663
rect 217 47607 303 47663
rect 359 47607 445 47663
rect 501 47607 587 47663
rect 643 47607 729 47663
rect 785 47607 871 47663
rect 927 47607 1013 47663
rect 1069 47607 1155 47663
rect 1211 47607 1297 47663
rect 1353 47607 1439 47663
rect 1495 47607 1581 47663
rect 1637 47607 1723 47663
rect 1779 47607 1865 47663
rect 1921 47607 2007 47663
rect 2063 47607 2149 47663
rect 2205 47607 2291 47663
rect 2347 47607 2433 47663
rect 2489 47607 2575 47663
rect 2631 47607 2717 47663
rect 2773 47607 2859 47663
rect 2915 47607 3001 47663
rect 3057 47607 3143 47663
rect 3199 47607 3285 47663
rect 3341 47607 3427 47663
rect 3483 47607 3569 47663
rect 3625 47607 3711 47663
rect 3767 47607 3853 47663
rect 3909 47607 3995 47663
rect 4051 47607 4137 47663
rect 4193 47607 4279 47663
rect 4335 47607 4421 47663
rect 4477 47607 4563 47663
rect 4619 47607 4705 47663
rect 4761 47607 4847 47663
rect 4903 47607 4989 47663
rect 5045 47607 5131 47663
rect 5187 47607 5273 47663
rect 5329 47607 5415 47663
rect 5471 47607 5557 47663
rect 5613 47607 5699 47663
rect 5755 47607 5841 47663
rect 5897 47607 5983 47663
rect 6039 47607 6125 47663
rect 6181 47607 6267 47663
rect 6323 47607 6409 47663
rect 6465 47607 6551 47663
rect 6607 47607 6693 47663
rect 6749 47607 6835 47663
rect 6891 47607 6977 47663
rect 7033 47607 7119 47663
rect 7175 47607 7261 47663
rect 7317 47607 7403 47663
rect 7459 47607 7545 47663
rect 7601 47607 7687 47663
rect 7743 47607 7829 47663
rect 7885 47607 7971 47663
rect 8027 47607 8113 47663
rect 8169 47607 8255 47663
rect 8311 47607 8397 47663
rect 8453 47607 8539 47663
rect 8595 47607 8681 47663
rect 8737 47607 8823 47663
rect 8879 47607 8965 47663
rect 9021 47607 9107 47663
rect 9163 47607 9249 47663
rect 9305 47607 9391 47663
rect 9447 47607 9533 47663
rect 9589 47607 9675 47663
rect 9731 47607 9817 47663
rect 9873 47607 9959 47663
rect 10015 47607 10101 47663
rect 10157 47607 10243 47663
rect 10299 47607 10385 47663
rect 10441 47607 10527 47663
rect 10583 47607 10669 47663
rect 10725 47607 10811 47663
rect 10867 47607 10953 47663
rect 11009 47607 11095 47663
rect 11151 47607 11237 47663
rect 11293 47607 11379 47663
rect 11435 47607 11521 47663
rect 11577 47607 11663 47663
rect 11719 47607 11805 47663
rect 11861 47607 11947 47663
rect 12003 47607 12089 47663
rect 12145 47607 12231 47663
rect 12287 47607 12373 47663
rect 12429 47607 12515 47663
rect 12571 47607 12657 47663
rect 12713 47607 12799 47663
rect 12855 47607 12941 47663
rect 12997 47607 13083 47663
rect 13139 47607 13225 47663
rect 13281 47607 13367 47663
rect 13423 47607 13509 47663
rect 13565 47607 13651 47663
rect 13707 47607 13793 47663
rect 13849 47607 13935 47663
rect 13991 47607 14077 47663
rect 14133 47607 14219 47663
rect 14275 47607 14361 47663
rect 14417 47607 14503 47663
rect 14559 47607 14645 47663
rect 14701 47607 14787 47663
rect 14843 47607 14853 47663
rect 151 47521 14853 47607
rect 151 47465 161 47521
rect 217 47465 303 47521
rect 359 47465 445 47521
rect 501 47465 587 47521
rect 643 47465 729 47521
rect 785 47465 871 47521
rect 927 47465 1013 47521
rect 1069 47465 1155 47521
rect 1211 47465 1297 47521
rect 1353 47465 1439 47521
rect 1495 47465 1581 47521
rect 1637 47465 1723 47521
rect 1779 47465 1865 47521
rect 1921 47465 2007 47521
rect 2063 47465 2149 47521
rect 2205 47465 2291 47521
rect 2347 47465 2433 47521
rect 2489 47465 2575 47521
rect 2631 47465 2717 47521
rect 2773 47465 2859 47521
rect 2915 47465 3001 47521
rect 3057 47465 3143 47521
rect 3199 47465 3285 47521
rect 3341 47465 3427 47521
rect 3483 47465 3569 47521
rect 3625 47465 3711 47521
rect 3767 47465 3853 47521
rect 3909 47465 3995 47521
rect 4051 47465 4137 47521
rect 4193 47465 4279 47521
rect 4335 47465 4421 47521
rect 4477 47465 4563 47521
rect 4619 47465 4705 47521
rect 4761 47465 4847 47521
rect 4903 47465 4989 47521
rect 5045 47465 5131 47521
rect 5187 47465 5273 47521
rect 5329 47465 5415 47521
rect 5471 47465 5557 47521
rect 5613 47465 5699 47521
rect 5755 47465 5841 47521
rect 5897 47465 5983 47521
rect 6039 47465 6125 47521
rect 6181 47465 6267 47521
rect 6323 47465 6409 47521
rect 6465 47465 6551 47521
rect 6607 47465 6693 47521
rect 6749 47465 6835 47521
rect 6891 47465 6977 47521
rect 7033 47465 7119 47521
rect 7175 47465 7261 47521
rect 7317 47465 7403 47521
rect 7459 47465 7545 47521
rect 7601 47465 7687 47521
rect 7743 47465 7829 47521
rect 7885 47465 7971 47521
rect 8027 47465 8113 47521
rect 8169 47465 8255 47521
rect 8311 47465 8397 47521
rect 8453 47465 8539 47521
rect 8595 47465 8681 47521
rect 8737 47465 8823 47521
rect 8879 47465 8965 47521
rect 9021 47465 9107 47521
rect 9163 47465 9249 47521
rect 9305 47465 9391 47521
rect 9447 47465 9533 47521
rect 9589 47465 9675 47521
rect 9731 47465 9817 47521
rect 9873 47465 9959 47521
rect 10015 47465 10101 47521
rect 10157 47465 10243 47521
rect 10299 47465 10385 47521
rect 10441 47465 10527 47521
rect 10583 47465 10669 47521
rect 10725 47465 10811 47521
rect 10867 47465 10953 47521
rect 11009 47465 11095 47521
rect 11151 47465 11237 47521
rect 11293 47465 11379 47521
rect 11435 47465 11521 47521
rect 11577 47465 11663 47521
rect 11719 47465 11805 47521
rect 11861 47465 11947 47521
rect 12003 47465 12089 47521
rect 12145 47465 12231 47521
rect 12287 47465 12373 47521
rect 12429 47465 12515 47521
rect 12571 47465 12657 47521
rect 12713 47465 12799 47521
rect 12855 47465 12941 47521
rect 12997 47465 13083 47521
rect 13139 47465 13225 47521
rect 13281 47465 13367 47521
rect 13423 47465 13509 47521
rect 13565 47465 13651 47521
rect 13707 47465 13793 47521
rect 13849 47465 13935 47521
rect 13991 47465 14077 47521
rect 14133 47465 14219 47521
rect 14275 47465 14361 47521
rect 14417 47465 14503 47521
rect 14559 47465 14645 47521
rect 14701 47465 14787 47521
rect 14843 47465 14853 47521
rect 151 47379 14853 47465
rect 151 47323 161 47379
rect 217 47323 303 47379
rect 359 47323 445 47379
rect 501 47323 587 47379
rect 643 47323 729 47379
rect 785 47323 871 47379
rect 927 47323 1013 47379
rect 1069 47323 1155 47379
rect 1211 47323 1297 47379
rect 1353 47323 1439 47379
rect 1495 47323 1581 47379
rect 1637 47323 1723 47379
rect 1779 47323 1865 47379
rect 1921 47323 2007 47379
rect 2063 47323 2149 47379
rect 2205 47323 2291 47379
rect 2347 47323 2433 47379
rect 2489 47323 2575 47379
rect 2631 47323 2717 47379
rect 2773 47323 2859 47379
rect 2915 47323 3001 47379
rect 3057 47323 3143 47379
rect 3199 47323 3285 47379
rect 3341 47323 3427 47379
rect 3483 47323 3569 47379
rect 3625 47323 3711 47379
rect 3767 47323 3853 47379
rect 3909 47323 3995 47379
rect 4051 47323 4137 47379
rect 4193 47323 4279 47379
rect 4335 47323 4421 47379
rect 4477 47323 4563 47379
rect 4619 47323 4705 47379
rect 4761 47323 4847 47379
rect 4903 47323 4989 47379
rect 5045 47323 5131 47379
rect 5187 47323 5273 47379
rect 5329 47323 5415 47379
rect 5471 47323 5557 47379
rect 5613 47323 5699 47379
rect 5755 47323 5841 47379
rect 5897 47323 5983 47379
rect 6039 47323 6125 47379
rect 6181 47323 6267 47379
rect 6323 47323 6409 47379
rect 6465 47323 6551 47379
rect 6607 47323 6693 47379
rect 6749 47323 6835 47379
rect 6891 47323 6977 47379
rect 7033 47323 7119 47379
rect 7175 47323 7261 47379
rect 7317 47323 7403 47379
rect 7459 47323 7545 47379
rect 7601 47323 7687 47379
rect 7743 47323 7829 47379
rect 7885 47323 7971 47379
rect 8027 47323 8113 47379
rect 8169 47323 8255 47379
rect 8311 47323 8397 47379
rect 8453 47323 8539 47379
rect 8595 47323 8681 47379
rect 8737 47323 8823 47379
rect 8879 47323 8965 47379
rect 9021 47323 9107 47379
rect 9163 47323 9249 47379
rect 9305 47323 9391 47379
rect 9447 47323 9533 47379
rect 9589 47323 9675 47379
rect 9731 47323 9817 47379
rect 9873 47323 9959 47379
rect 10015 47323 10101 47379
rect 10157 47323 10243 47379
rect 10299 47323 10385 47379
rect 10441 47323 10527 47379
rect 10583 47323 10669 47379
rect 10725 47323 10811 47379
rect 10867 47323 10953 47379
rect 11009 47323 11095 47379
rect 11151 47323 11237 47379
rect 11293 47323 11379 47379
rect 11435 47323 11521 47379
rect 11577 47323 11663 47379
rect 11719 47323 11805 47379
rect 11861 47323 11947 47379
rect 12003 47323 12089 47379
rect 12145 47323 12231 47379
rect 12287 47323 12373 47379
rect 12429 47323 12515 47379
rect 12571 47323 12657 47379
rect 12713 47323 12799 47379
rect 12855 47323 12941 47379
rect 12997 47323 13083 47379
rect 13139 47323 13225 47379
rect 13281 47323 13367 47379
rect 13423 47323 13509 47379
rect 13565 47323 13651 47379
rect 13707 47323 13793 47379
rect 13849 47323 13935 47379
rect 13991 47323 14077 47379
rect 14133 47323 14219 47379
rect 14275 47323 14361 47379
rect 14417 47323 14503 47379
rect 14559 47323 14645 47379
rect 14701 47323 14787 47379
rect 14843 47323 14853 47379
rect 151 47237 14853 47323
rect 151 47181 161 47237
rect 217 47181 303 47237
rect 359 47181 445 47237
rect 501 47181 587 47237
rect 643 47181 729 47237
rect 785 47181 871 47237
rect 927 47181 1013 47237
rect 1069 47181 1155 47237
rect 1211 47181 1297 47237
rect 1353 47181 1439 47237
rect 1495 47181 1581 47237
rect 1637 47181 1723 47237
rect 1779 47181 1865 47237
rect 1921 47181 2007 47237
rect 2063 47181 2149 47237
rect 2205 47181 2291 47237
rect 2347 47181 2433 47237
rect 2489 47181 2575 47237
rect 2631 47181 2717 47237
rect 2773 47181 2859 47237
rect 2915 47181 3001 47237
rect 3057 47181 3143 47237
rect 3199 47181 3285 47237
rect 3341 47181 3427 47237
rect 3483 47181 3569 47237
rect 3625 47181 3711 47237
rect 3767 47181 3853 47237
rect 3909 47181 3995 47237
rect 4051 47181 4137 47237
rect 4193 47181 4279 47237
rect 4335 47181 4421 47237
rect 4477 47181 4563 47237
rect 4619 47181 4705 47237
rect 4761 47181 4847 47237
rect 4903 47181 4989 47237
rect 5045 47181 5131 47237
rect 5187 47181 5273 47237
rect 5329 47181 5415 47237
rect 5471 47181 5557 47237
rect 5613 47181 5699 47237
rect 5755 47181 5841 47237
rect 5897 47181 5983 47237
rect 6039 47181 6125 47237
rect 6181 47181 6267 47237
rect 6323 47181 6409 47237
rect 6465 47181 6551 47237
rect 6607 47181 6693 47237
rect 6749 47181 6835 47237
rect 6891 47181 6977 47237
rect 7033 47181 7119 47237
rect 7175 47181 7261 47237
rect 7317 47181 7403 47237
rect 7459 47181 7545 47237
rect 7601 47181 7687 47237
rect 7743 47181 7829 47237
rect 7885 47181 7971 47237
rect 8027 47181 8113 47237
rect 8169 47181 8255 47237
rect 8311 47181 8397 47237
rect 8453 47181 8539 47237
rect 8595 47181 8681 47237
rect 8737 47181 8823 47237
rect 8879 47181 8965 47237
rect 9021 47181 9107 47237
rect 9163 47181 9249 47237
rect 9305 47181 9391 47237
rect 9447 47181 9533 47237
rect 9589 47181 9675 47237
rect 9731 47181 9817 47237
rect 9873 47181 9959 47237
rect 10015 47181 10101 47237
rect 10157 47181 10243 47237
rect 10299 47181 10385 47237
rect 10441 47181 10527 47237
rect 10583 47181 10669 47237
rect 10725 47181 10811 47237
rect 10867 47181 10953 47237
rect 11009 47181 11095 47237
rect 11151 47181 11237 47237
rect 11293 47181 11379 47237
rect 11435 47181 11521 47237
rect 11577 47181 11663 47237
rect 11719 47181 11805 47237
rect 11861 47181 11947 47237
rect 12003 47181 12089 47237
rect 12145 47181 12231 47237
rect 12287 47181 12373 47237
rect 12429 47181 12515 47237
rect 12571 47181 12657 47237
rect 12713 47181 12799 47237
rect 12855 47181 12941 47237
rect 12997 47181 13083 47237
rect 13139 47181 13225 47237
rect 13281 47181 13367 47237
rect 13423 47181 13509 47237
rect 13565 47181 13651 47237
rect 13707 47181 13793 47237
rect 13849 47181 13935 47237
rect 13991 47181 14077 47237
rect 14133 47181 14219 47237
rect 14275 47181 14361 47237
rect 14417 47181 14503 47237
rect 14559 47181 14645 47237
rect 14701 47181 14787 47237
rect 14843 47181 14853 47237
rect 151 47095 14853 47181
rect 151 47039 161 47095
rect 217 47039 303 47095
rect 359 47039 445 47095
rect 501 47039 587 47095
rect 643 47039 729 47095
rect 785 47039 871 47095
rect 927 47039 1013 47095
rect 1069 47039 1155 47095
rect 1211 47039 1297 47095
rect 1353 47039 1439 47095
rect 1495 47039 1581 47095
rect 1637 47039 1723 47095
rect 1779 47039 1865 47095
rect 1921 47039 2007 47095
rect 2063 47039 2149 47095
rect 2205 47039 2291 47095
rect 2347 47039 2433 47095
rect 2489 47039 2575 47095
rect 2631 47039 2717 47095
rect 2773 47039 2859 47095
rect 2915 47039 3001 47095
rect 3057 47039 3143 47095
rect 3199 47039 3285 47095
rect 3341 47039 3427 47095
rect 3483 47039 3569 47095
rect 3625 47039 3711 47095
rect 3767 47039 3853 47095
rect 3909 47039 3995 47095
rect 4051 47039 4137 47095
rect 4193 47039 4279 47095
rect 4335 47039 4421 47095
rect 4477 47039 4563 47095
rect 4619 47039 4705 47095
rect 4761 47039 4847 47095
rect 4903 47039 4989 47095
rect 5045 47039 5131 47095
rect 5187 47039 5273 47095
rect 5329 47039 5415 47095
rect 5471 47039 5557 47095
rect 5613 47039 5699 47095
rect 5755 47039 5841 47095
rect 5897 47039 5983 47095
rect 6039 47039 6125 47095
rect 6181 47039 6267 47095
rect 6323 47039 6409 47095
rect 6465 47039 6551 47095
rect 6607 47039 6693 47095
rect 6749 47039 6835 47095
rect 6891 47039 6977 47095
rect 7033 47039 7119 47095
rect 7175 47039 7261 47095
rect 7317 47039 7403 47095
rect 7459 47039 7545 47095
rect 7601 47039 7687 47095
rect 7743 47039 7829 47095
rect 7885 47039 7971 47095
rect 8027 47039 8113 47095
rect 8169 47039 8255 47095
rect 8311 47039 8397 47095
rect 8453 47039 8539 47095
rect 8595 47039 8681 47095
rect 8737 47039 8823 47095
rect 8879 47039 8965 47095
rect 9021 47039 9107 47095
rect 9163 47039 9249 47095
rect 9305 47039 9391 47095
rect 9447 47039 9533 47095
rect 9589 47039 9675 47095
rect 9731 47039 9817 47095
rect 9873 47039 9959 47095
rect 10015 47039 10101 47095
rect 10157 47039 10243 47095
rect 10299 47039 10385 47095
rect 10441 47039 10527 47095
rect 10583 47039 10669 47095
rect 10725 47039 10811 47095
rect 10867 47039 10953 47095
rect 11009 47039 11095 47095
rect 11151 47039 11237 47095
rect 11293 47039 11379 47095
rect 11435 47039 11521 47095
rect 11577 47039 11663 47095
rect 11719 47039 11805 47095
rect 11861 47039 11947 47095
rect 12003 47039 12089 47095
rect 12145 47039 12231 47095
rect 12287 47039 12373 47095
rect 12429 47039 12515 47095
rect 12571 47039 12657 47095
rect 12713 47039 12799 47095
rect 12855 47039 12941 47095
rect 12997 47039 13083 47095
rect 13139 47039 13225 47095
rect 13281 47039 13367 47095
rect 13423 47039 13509 47095
rect 13565 47039 13651 47095
rect 13707 47039 13793 47095
rect 13849 47039 13935 47095
rect 13991 47039 14077 47095
rect 14133 47039 14219 47095
rect 14275 47039 14361 47095
rect 14417 47039 14503 47095
rect 14559 47039 14645 47095
rect 14701 47039 14787 47095
rect 14843 47039 14853 47095
rect 151 46953 14853 47039
rect 151 46897 161 46953
rect 217 46897 303 46953
rect 359 46897 445 46953
rect 501 46897 587 46953
rect 643 46897 729 46953
rect 785 46897 871 46953
rect 927 46897 1013 46953
rect 1069 46897 1155 46953
rect 1211 46897 1297 46953
rect 1353 46897 1439 46953
rect 1495 46897 1581 46953
rect 1637 46897 1723 46953
rect 1779 46897 1865 46953
rect 1921 46897 2007 46953
rect 2063 46897 2149 46953
rect 2205 46897 2291 46953
rect 2347 46897 2433 46953
rect 2489 46897 2575 46953
rect 2631 46897 2717 46953
rect 2773 46897 2859 46953
rect 2915 46897 3001 46953
rect 3057 46897 3143 46953
rect 3199 46897 3285 46953
rect 3341 46897 3427 46953
rect 3483 46897 3569 46953
rect 3625 46897 3711 46953
rect 3767 46897 3853 46953
rect 3909 46897 3995 46953
rect 4051 46897 4137 46953
rect 4193 46897 4279 46953
rect 4335 46897 4421 46953
rect 4477 46897 4563 46953
rect 4619 46897 4705 46953
rect 4761 46897 4847 46953
rect 4903 46897 4989 46953
rect 5045 46897 5131 46953
rect 5187 46897 5273 46953
rect 5329 46897 5415 46953
rect 5471 46897 5557 46953
rect 5613 46897 5699 46953
rect 5755 46897 5841 46953
rect 5897 46897 5983 46953
rect 6039 46897 6125 46953
rect 6181 46897 6267 46953
rect 6323 46897 6409 46953
rect 6465 46897 6551 46953
rect 6607 46897 6693 46953
rect 6749 46897 6835 46953
rect 6891 46897 6977 46953
rect 7033 46897 7119 46953
rect 7175 46897 7261 46953
rect 7317 46897 7403 46953
rect 7459 46897 7545 46953
rect 7601 46897 7687 46953
rect 7743 46897 7829 46953
rect 7885 46897 7971 46953
rect 8027 46897 8113 46953
rect 8169 46897 8255 46953
rect 8311 46897 8397 46953
rect 8453 46897 8539 46953
rect 8595 46897 8681 46953
rect 8737 46897 8823 46953
rect 8879 46897 8965 46953
rect 9021 46897 9107 46953
rect 9163 46897 9249 46953
rect 9305 46897 9391 46953
rect 9447 46897 9533 46953
rect 9589 46897 9675 46953
rect 9731 46897 9817 46953
rect 9873 46897 9959 46953
rect 10015 46897 10101 46953
rect 10157 46897 10243 46953
rect 10299 46897 10385 46953
rect 10441 46897 10527 46953
rect 10583 46897 10669 46953
rect 10725 46897 10811 46953
rect 10867 46897 10953 46953
rect 11009 46897 11095 46953
rect 11151 46897 11237 46953
rect 11293 46897 11379 46953
rect 11435 46897 11521 46953
rect 11577 46897 11663 46953
rect 11719 46897 11805 46953
rect 11861 46897 11947 46953
rect 12003 46897 12089 46953
rect 12145 46897 12231 46953
rect 12287 46897 12373 46953
rect 12429 46897 12515 46953
rect 12571 46897 12657 46953
rect 12713 46897 12799 46953
rect 12855 46897 12941 46953
rect 12997 46897 13083 46953
rect 13139 46897 13225 46953
rect 13281 46897 13367 46953
rect 13423 46897 13509 46953
rect 13565 46897 13651 46953
rect 13707 46897 13793 46953
rect 13849 46897 13935 46953
rect 13991 46897 14077 46953
rect 14133 46897 14219 46953
rect 14275 46897 14361 46953
rect 14417 46897 14503 46953
rect 14559 46897 14645 46953
rect 14701 46897 14787 46953
rect 14843 46897 14853 46953
rect 151 46811 14853 46897
rect 151 46755 161 46811
rect 217 46755 303 46811
rect 359 46755 445 46811
rect 501 46755 587 46811
rect 643 46755 729 46811
rect 785 46755 871 46811
rect 927 46755 1013 46811
rect 1069 46755 1155 46811
rect 1211 46755 1297 46811
rect 1353 46755 1439 46811
rect 1495 46755 1581 46811
rect 1637 46755 1723 46811
rect 1779 46755 1865 46811
rect 1921 46755 2007 46811
rect 2063 46755 2149 46811
rect 2205 46755 2291 46811
rect 2347 46755 2433 46811
rect 2489 46755 2575 46811
rect 2631 46755 2717 46811
rect 2773 46755 2859 46811
rect 2915 46755 3001 46811
rect 3057 46755 3143 46811
rect 3199 46755 3285 46811
rect 3341 46755 3427 46811
rect 3483 46755 3569 46811
rect 3625 46755 3711 46811
rect 3767 46755 3853 46811
rect 3909 46755 3995 46811
rect 4051 46755 4137 46811
rect 4193 46755 4279 46811
rect 4335 46755 4421 46811
rect 4477 46755 4563 46811
rect 4619 46755 4705 46811
rect 4761 46755 4847 46811
rect 4903 46755 4989 46811
rect 5045 46755 5131 46811
rect 5187 46755 5273 46811
rect 5329 46755 5415 46811
rect 5471 46755 5557 46811
rect 5613 46755 5699 46811
rect 5755 46755 5841 46811
rect 5897 46755 5983 46811
rect 6039 46755 6125 46811
rect 6181 46755 6267 46811
rect 6323 46755 6409 46811
rect 6465 46755 6551 46811
rect 6607 46755 6693 46811
rect 6749 46755 6835 46811
rect 6891 46755 6977 46811
rect 7033 46755 7119 46811
rect 7175 46755 7261 46811
rect 7317 46755 7403 46811
rect 7459 46755 7545 46811
rect 7601 46755 7687 46811
rect 7743 46755 7829 46811
rect 7885 46755 7971 46811
rect 8027 46755 8113 46811
rect 8169 46755 8255 46811
rect 8311 46755 8397 46811
rect 8453 46755 8539 46811
rect 8595 46755 8681 46811
rect 8737 46755 8823 46811
rect 8879 46755 8965 46811
rect 9021 46755 9107 46811
rect 9163 46755 9249 46811
rect 9305 46755 9391 46811
rect 9447 46755 9533 46811
rect 9589 46755 9675 46811
rect 9731 46755 9817 46811
rect 9873 46755 9959 46811
rect 10015 46755 10101 46811
rect 10157 46755 10243 46811
rect 10299 46755 10385 46811
rect 10441 46755 10527 46811
rect 10583 46755 10669 46811
rect 10725 46755 10811 46811
rect 10867 46755 10953 46811
rect 11009 46755 11095 46811
rect 11151 46755 11237 46811
rect 11293 46755 11379 46811
rect 11435 46755 11521 46811
rect 11577 46755 11663 46811
rect 11719 46755 11805 46811
rect 11861 46755 11947 46811
rect 12003 46755 12089 46811
rect 12145 46755 12231 46811
rect 12287 46755 12373 46811
rect 12429 46755 12515 46811
rect 12571 46755 12657 46811
rect 12713 46755 12799 46811
rect 12855 46755 12941 46811
rect 12997 46755 13083 46811
rect 13139 46755 13225 46811
rect 13281 46755 13367 46811
rect 13423 46755 13509 46811
rect 13565 46755 13651 46811
rect 13707 46755 13793 46811
rect 13849 46755 13935 46811
rect 13991 46755 14077 46811
rect 14133 46755 14219 46811
rect 14275 46755 14361 46811
rect 14417 46755 14503 46811
rect 14559 46755 14645 46811
rect 14701 46755 14787 46811
rect 14843 46755 14853 46811
rect 151 46669 14853 46755
rect 151 46613 161 46669
rect 217 46613 303 46669
rect 359 46613 445 46669
rect 501 46613 587 46669
rect 643 46613 729 46669
rect 785 46613 871 46669
rect 927 46613 1013 46669
rect 1069 46613 1155 46669
rect 1211 46613 1297 46669
rect 1353 46613 1439 46669
rect 1495 46613 1581 46669
rect 1637 46613 1723 46669
rect 1779 46613 1865 46669
rect 1921 46613 2007 46669
rect 2063 46613 2149 46669
rect 2205 46613 2291 46669
rect 2347 46613 2433 46669
rect 2489 46613 2575 46669
rect 2631 46613 2717 46669
rect 2773 46613 2859 46669
rect 2915 46613 3001 46669
rect 3057 46613 3143 46669
rect 3199 46613 3285 46669
rect 3341 46613 3427 46669
rect 3483 46613 3569 46669
rect 3625 46613 3711 46669
rect 3767 46613 3853 46669
rect 3909 46613 3995 46669
rect 4051 46613 4137 46669
rect 4193 46613 4279 46669
rect 4335 46613 4421 46669
rect 4477 46613 4563 46669
rect 4619 46613 4705 46669
rect 4761 46613 4847 46669
rect 4903 46613 4989 46669
rect 5045 46613 5131 46669
rect 5187 46613 5273 46669
rect 5329 46613 5415 46669
rect 5471 46613 5557 46669
rect 5613 46613 5699 46669
rect 5755 46613 5841 46669
rect 5897 46613 5983 46669
rect 6039 46613 6125 46669
rect 6181 46613 6267 46669
rect 6323 46613 6409 46669
rect 6465 46613 6551 46669
rect 6607 46613 6693 46669
rect 6749 46613 6835 46669
rect 6891 46613 6977 46669
rect 7033 46613 7119 46669
rect 7175 46613 7261 46669
rect 7317 46613 7403 46669
rect 7459 46613 7545 46669
rect 7601 46613 7687 46669
rect 7743 46613 7829 46669
rect 7885 46613 7971 46669
rect 8027 46613 8113 46669
rect 8169 46613 8255 46669
rect 8311 46613 8397 46669
rect 8453 46613 8539 46669
rect 8595 46613 8681 46669
rect 8737 46613 8823 46669
rect 8879 46613 8965 46669
rect 9021 46613 9107 46669
rect 9163 46613 9249 46669
rect 9305 46613 9391 46669
rect 9447 46613 9533 46669
rect 9589 46613 9675 46669
rect 9731 46613 9817 46669
rect 9873 46613 9959 46669
rect 10015 46613 10101 46669
rect 10157 46613 10243 46669
rect 10299 46613 10385 46669
rect 10441 46613 10527 46669
rect 10583 46613 10669 46669
rect 10725 46613 10811 46669
rect 10867 46613 10953 46669
rect 11009 46613 11095 46669
rect 11151 46613 11237 46669
rect 11293 46613 11379 46669
rect 11435 46613 11521 46669
rect 11577 46613 11663 46669
rect 11719 46613 11805 46669
rect 11861 46613 11947 46669
rect 12003 46613 12089 46669
rect 12145 46613 12231 46669
rect 12287 46613 12373 46669
rect 12429 46613 12515 46669
rect 12571 46613 12657 46669
rect 12713 46613 12799 46669
rect 12855 46613 12941 46669
rect 12997 46613 13083 46669
rect 13139 46613 13225 46669
rect 13281 46613 13367 46669
rect 13423 46613 13509 46669
rect 13565 46613 13651 46669
rect 13707 46613 13793 46669
rect 13849 46613 13935 46669
rect 13991 46613 14077 46669
rect 14133 46613 14219 46669
rect 14275 46613 14361 46669
rect 14417 46613 14503 46669
rect 14559 46613 14645 46669
rect 14701 46613 14787 46669
rect 14843 46613 14853 46669
rect 151 46527 14853 46613
rect 151 46471 161 46527
rect 217 46471 303 46527
rect 359 46471 445 46527
rect 501 46471 587 46527
rect 643 46471 729 46527
rect 785 46471 871 46527
rect 927 46471 1013 46527
rect 1069 46471 1155 46527
rect 1211 46471 1297 46527
rect 1353 46471 1439 46527
rect 1495 46471 1581 46527
rect 1637 46471 1723 46527
rect 1779 46471 1865 46527
rect 1921 46471 2007 46527
rect 2063 46471 2149 46527
rect 2205 46471 2291 46527
rect 2347 46471 2433 46527
rect 2489 46471 2575 46527
rect 2631 46471 2717 46527
rect 2773 46471 2859 46527
rect 2915 46471 3001 46527
rect 3057 46471 3143 46527
rect 3199 46471 3285 46527
rect 3341 46471 3427 46527
rect 3483 46471 3569 46527
rect 3625 46471 3711 46527
rect 3767 46471 3853 46527
rect 3909 46471 3995 46527
rect 4051 46471 4137 46527
rect 4193 46471 4279 46527
rect 4335 46471 4421 46527
rect 4477 46471 4563 46527
rect 4619 46471 4705 46527
rect 4761 46471 4847 46527
rect 4903 46471 4989 46527
rect 5045 46471 5131 46527
rect 5187 46471 5273 46527
rect 5329 46471 5415 46527
rect 5471 46471 5557 46527
rect 5613 46471 5699 46527
rect 5755 46471 5841 46527
rect 5897 46471 5983 46527
rect 6039 46471 6125 46527
rect 6181 46471 6267 46527
rect 6323 46471 6409 46527
rect 6465 46471 6551 46527
rect 6607 46471 6693 46527
rect 6749 46471 6835 46527
rect 6891 46471 6977 46527
rect 7033 46471 7119 46527
rect 7175 46471 7261 46527
rect 7317 46471 7403 46527
rect 7459 46471 7545 46527
rect 7601 46471 7687 46527
rect 7743 46471 7829 46527
rect 7885 46471 7971 46527
rect 8027 46471 8113 46527
rect 8169 46471 8255 46527
rect 8311 46471 8397 46527
rect 8453 46471 8539 46527
rect 8595 46471 8681 46527
rect 8737 46471 8823 46527
rect 8879 46471 8965 46527
rect 9021 46471 9107 46527
rect 9163 46471 9249 46527
rect 9305 46471 9391 46527
rect 9447 46471 9533 46527
rect 9589 46471 9675 46527
rect 9731 46471 9817 46527
rect 9873 46471 9959 46527
rect 10015 46471 10101 46527
rect 10157 46471 10243 46527
rect 10299 46471 10385 46527
rect 10441 46471 10527 46527
rect 10583 46471 10669 46527
rect 10725 46471 10811 46527
rect 10867 46471 10953 46527
rect 11009 46471 11095 46527
rect 11151 46471 11237 46527
rect 11293 46471 11379 46527
rect 11435 46471 11521 46527
rect 11577 46471 11663 46527
rect 11719 46471 11805 46527
rect 11861 46471 11947 46527
rect 12003 46471 12089 46527
rect 12145 46471 12231 46527
rect 12287 46471 12373 46527
rect 12429 46471 12515 46527
rect 12571 46471 12657 46527
rect 12713 46471 12799 46527
rect 12855 46471 12941 46527
rect 12997 46471 13083 46527
rect 13139 46471 13225 46527
rect 13281 46471 13367 46527
rect 13423 46471 13509 46527
rect 13565 46471 13651 46527
rect 13707 46471 13793 46527
rect 13849 46471 13935 46527
rect 13991 46471 14077 46527
rect 14133 46471 14219 46527
rect 14275 46471 14361 46527
rect 14417 46471 14503 46527
rect 14559 46471 14645 46527
rect 14701 46471 14787 46527
rect 14843 46471 14853 46527
rect 151 46385 14853 46471
rect 151 46329 161 46385
rect 217 46329 303 46385
rect 359 46329 445 46385
rect 501 46329 587 46385
rect 643 46329 729 46385
rect 785 46329 871 46385
rect 927 46329 1013 46385
rect 1069 46329 1155 46385
rect 1211 46329 1297 46385
rect 1353 46329 1439 46385
rect 1495 46329 1581 46385
rect 1637 46329 1723 46385
rect 1779 46329 1865 46385
rect 1921 46329 2007 46385
rect 2063 46329 2149 46385
rect 2205 46329 2291 46385
rect 2347 46329 2433 46385
rect 2489 46329 2575 46385
rect 2631 46329 2717 46385
rect 2773 46329 2859 46385
rect 2915 46329 3001 46385
rect 3057 46329 3143 46385
rect 3199 46329 3285 46385
rect 3341 46329 3427 46385
rect 3483 46329 3569 46385
rect 3625 46329 3711 46385
rect 3767 46329 3853 46385
rect 3909 46329 3995 46385
rect 4051 46329 4137 46385
rect 4193 46329 4279 46385
rect 4335 46329 4421 46385
rect 4477 46329 4563 46385
rect 4619 46329 4705 46385
rect 4761 46329 4847 46385
rect 4903 46329 4989 46385
rect 5045 46329 5131 46385
rect 5187 46329 5273 46385
rect 5329 46329 5415 46385
rect 5471 46329 5557 46385
rect 5613 46329 5699 46385
rect 5755 46329 5841 46385
rect 5897 46329 5983 46385
rect 6039 46329 6125 46385
rect 6181 46329 6267 46385
rect 6323 46329 6409 46385
rect 6465 46329 6551 46385
rect 6607 46329 6693 46385
rect 6749 46329 6835 46385
rect 6891 46329 6977 46385
rect 7033 46329 7119 46385
rect 7175 46329 7261 46385
rect 7317 46329 7403 46385
rect 7459 46329 7545 46385
rect 7601 46329 7687 46385
rect 7743 46329 7829 46385
rect 7885 46329 7971 46385
rect 8027 46329 8113 46385
rect 8169 46329 8255 46385
rect 8311 46329 8397 46385
rect 8453 46329 8539 46385
rect 8595 46329 8681 46385
rect 8737 46329 8823 46385
rect 8879 46329 8965 46385
rect 9021 46329 9107 46385
rect 9163 46329 9249 46385
rect 9305 46329 9391 46385
rect 9447 46329 9533 46385
rect 9589 46329 9675 46385
rect 9731 46329 9817 46385
rect 9873 46329 9959 46385
rect 10015 46329 10101 46385
rect 10157 46329 10243 46385
rect 10299 46329 10385 46385
rect 10441 46329 10527 46385
rect 10583 46329 10669 46385
rect 10725 46329 10811 46385
rect 10867 46329 10953 46385
rect 11009 46329 11095 46385
rect 11151 46329 11237 46385
rect 11293 46329 11379 46385
rect 11435 46329 11521 46385
rect 11577 46329 11663 46385
rect 11719 46329 11805 46385
rect 11861 46329 11947 46385
rect 12003 46329 12089 46385
rect 12145 46329 12231 46385
rect 12287 46329 12373 46385
rect 12429 46329 12515 46385
rect 12571 46329 12657 46385
rect 12713 46329 12799 46385
rect 12855 46329 12941 46385
rect 12997 46329 13083 46385
rect 13139 46329 13225 46385
rect 13281 46329 13367 46385
rect 13423 46329 13509 46385
rect 13565 46329 13651 46385
rect 13707 46329 13793 46385
rect 13849 46329 13935 46385
rect 13991 46329 14077 46385
rect 14133 46329 14219 46385
rect 14275 46329 14361 46385
rect 14417 46329 14503 46385
rect 14559 46329 14645 46385
rect 14701 46329 14787 46385
rect 14843 46329 14853 46385
rect 151 46243 14853 46329
rect 151 46187 161 46243
rect 217 46187 303 46243
rect 359 46187 445 46243
rect 501 46187 587 46243
rect 643 46187 729 46243
rect 785 46187 871 46243
rect 927 46187 1013 46243
rect 1069 46187 1155 46243
rect 1211 46187 1297 46243
rect 1353 46187 1439 46243
rect 1495 46187 1581 46243
rect 1637 46187 1723 46243
rect 1779 46187 1865 46243
rect 1921 46187 2007 46243
rect 2063 46187 2149 46243
rect 2205 46187 2291 46243
rect 2347 46187 2433 46243
rect 2489 46187 2575 46243
rect 2631 46187 2717 46243
rect 2773 46187 2859 46243
rect 2915 46187 3001 46243
rect 3057 46187 3143 46243
rect 3199 46187 3285 46243
rect 3341 46187 3427 46243
rect 3483 46187 3569 46243
rect 3625 46187 3711 46243
rect 3767 46187 3853 46243
rect 3909 46187 3995 46243
rect 4051 46187 4137 46243
rect 4193 46187 4279 46243
rect 4335 46187 4421 46243
rect 4477 46187 4563 46243
rect 4619 46187 4705 46243
rect 4761 46187 4847 46243
rect 4903 46187 4989 46243
rect 5045 46187 5131 46243
rect 5187 46187 5273 46243
rect 5329 46187 5415 46243
rect 5471 46187 5557 46243
rect 5613 46187 5699 46243
rect 5755 46187 5841 46243
rect 5897 46187 5983 46243
rect 6039 46187 6125 46243
rect 6181 46187 6267 46243
rect 6323 46187 6409 46243
rect 6465 46187 6551 46243
rect 6607 46187 6693 46243
rect 6749 46187 6835 46243
rect 6891 46187 6977 46243
rect 7033 46187 7119 46243
rect 7175 46187 7261 46243
rect 7317 46187 7403 46243
rect 7459 46187 7545 46243
rect 7601 46187 7687 46243
rect 7743 46187 7829 46243
rect 7885 46187 7971 46243
rect 8027 46187 8113 46243
rect 8169 46187 8255 46243
rect 8311 46187 8397 46243
rect 8453 46187 8539 46243
rect 8595 46187 8681 46243
rect 8737 46187 8823 46243
rect 8879 46187 8965 46243
rect 9021 46187 9107 46243
rect 9163 46187 9249 46243
rect 9305 46187 9391 46243
rect 9447 46187 9533 46243
rect 9589 46187 9675 46243
rect 9731 46187 9817 46243
rect 9873 46187 9959 46243
rect 10015 46187 10101 46243
rect 10157 46187 10243 46243
rect 10299 46187 10385 46243
rect 10441 46187 10527 46243
rect 10583 46187 10669 46243
rect 10725 46187 10811 46243
rect 10867 46187 10953 46243
rect 11009 46187 11095 46243
rect 11151 46187 11237 46243
rect 11293 46187 11379 46243
rect 11435 46187 11521 46243
rect 11577 46187 11663 46243
rect 11719 46187 11805 46243
rect 11861 46187 11947 46243
rect 12003 46187 12089 46243
rect 12145 46187 12231 46243
rect 12287 46187 12373 46243
rect 12429 46187 12515 46243
rect 12571 46187 12657 46243
rect 12713 46187 12799 46243
rect 12855 46187 12941 46243
rect 12997 46187 13083 46243
rect 13139 46187 13225 46243
rect 13281 46187 13367 46243
rect 13423 46187 13509 46243
rect 13565 46187 13651 46243
rect 13707 46187 13793 46243
rect 13849 46187 13935 46243
rect 13991 46187 14077 46243
rect 14133 46187 14219 46243
rect 14275 46187 14361 46243
rect 14417 46187 14503 46243
rect 14559 46187 14645 46243
rect 14701 46187 14787 46243
rect 14843 46187 14853 46243
rect 151 46101 14853 46187
rect 151 46045 161 46101
rect 217 46045 303 46101
rect 359 46045 445 46101
rect 501 46045 587 46101
rect 643 46045 729 46101
rect 785 46045 871 46101
rect 927 46045 1013 46101
rect 1069 46045 1155 46101
rect 1211 46045 1297 46101
rect 1353 46045 1439 46101
rect 1495 46045 1581 46101
rect 1637 46045 1723 46101
rect 1779 46045 1865 46101
rect 1921 46045 2007 46101
rect 2063 46045 2149 46101
rect 2205 46045 2291 46101
rect 2347 46045 2433 46101
rect 2489 46045 2575 46101
rect 2631 46045 2717 46101
rect 2773 46045 2859 46101
rect 2915 46045 3001 46101
rect 3057 46045 3143 46101
rect 3199 46045 3285 46101
rect 3341 46045 3427 46101
rect 3483 46045 3569 46101
rect 3625 46045 3711 46101
rect 3767 46045 3853 46101
rect 3909 46045 3995 46101
rect 4051 46045 4137 46101
rect 4193 46045 4279 46101
rect 4335 46045 4421 46101
rect 4477 46045 4563 46101
rect 4619 46045 4705 46101
rect 4761 46045 4847 46101
rect 4903 46045 4989 46101
rect 5045 46045 5131 46101
rect 5187 46045 5273 46101
rect 5329 46045 5415 46101
rect 5471 46045 5557 46101
rect 5613 46045 5699 46101
rect 5755 46045 5841 46101
rect 5897 46045 5983 46101
rect 6039 46045 6125 46101
rect 6181 46045 6267 46101
rect 6323 46045 6409 46101
rect 6465 46045 6551 46101
rect 6607 46045 6693 46101
rect 6749 46045 6835 46101
rect 6891 46045 6977 46101
rect 7033 46045 7119 46101
rect 7175 46045 7261 46101
rect 7317 46045 7403 46101
rect 7459 46045 7545 46101
rect 7601 46045 7687 46101
rect 7743 46045 7829 46101
rect 7885 46045 7971 46101
rect 8027 46045 8113 46101
rect 8169 46045 8255 46101
rect 8311 46045 8397 46101
rect 8453 46045 8539 46101
rect 8595 46045 8681 46101
rect 8737 46045 8823 46101
rect 8879 46045 8965 46101
rect 9021 46045 9107 46101
rect 9163 46045 9249 46101
rect 9305 46045 9391 46101
rect 9447 46045 9533 46101
rect 9589 46045 9675 46101
rect 9731 46045 9817 46101
rect 9873 46045 9959 46101
rect 10015 46045 10101 46101
rect 10157 46045 10243 46101
rect 10299 46045 10385 46101
rect 10441 46045 10527 46101
rect 10583 46045 10669 46101
rect 10725 46045 10811 46101
rect 10867 46045 10953 46101
rect 11009 46045 11095 46101
rect 11151 46045 11237 46101
rect 11293 46045 11379 46101
rect 11435 46045 11521 46101
rect 11577 46045 11663 46101
rect 11719 46045 11805 46101
rect 11861 46045 11947 46101
rect 12003 46045 12089 46101
rect 12145 46045 12231 46101
rect 12287 46045 12373 46101
rect 12429 46045 12515 46101
rect 12571 46045 12657 46101
rect 12713 46045 12799 46101
rect 12855 46045 12941 46101
rect 12997 46045 13083 46101
rect 13139 46045 13225 46101
rect 13281 46045 13367 46101
rect 13423 46045 13509 46101
rect 13565 46045 13651 46101
rect 13707 46045 13793 46101
rect 13849 46045 13935 46101
rect 13991 46045 14077 46101
rect 14133 46045 14219 46101
rect 14275 46045 14361 46101
rect 14417 46045 14503 46101
rect 14559 46045 14645 46101
rect 14701 46045 14787 46101
rect 14843 46045 14853 46101
rect 151 46035 14853 46045
rect 151 45741 14853 45751
rect 151 45685 161 45741
rect 217 45685 303 45741
rect 359 45685 445 45741
rect 501 45685 587 45741
rect 643 45685 729 45741
rect 785 45685 871 45741
rect 927 45685 1013 45741
rect 1069 45685 1155 45741
rect 1211 45685 1297 45741
rect 1353 45685 1439 45741
rect 1495 45685 1581 45741
rect 1637 45685 1723 45741
rect 1779 45685 1865 45741
rect 1921 45685 2007 45741
rect 2063 45685 2149 45741
rect 2205 45685 2291 45741
rect 2347 45685 2433 45741
rect 2489 45685 2575 45741
rect 2631 45685 2717 45741
rect 2773 45685 2859 45741
rect 2915 45685 3001 45741
rect 3057 45685 3143 45741
rect 3199 45685 3285 45741
rect 3341 45685 3427 45741
rect 3483 45685 3569 45741
rect 3625 45685 3711 45741
rect 3767 45685 3853 45741
rect 3909 45685 3995 45741
rect 4051 45685 4137 45741
rect 4193 45685 4279 45741
rect 4335 45685 4421 45741
rect 4477 45685 4563 45741
rect 4619 45685 4705 45741
rect 4761 45685 4847 45741
rect 4903 45685 4989 45741
rect 5045 45685 5131 45741
rect 5187 45685 5273 45741
rect 5329 45685 5415 45741
rect 5471 45685 5557 45741
rect 5613 45685 5699 45741
rect 5755 45685 5841 45741
rect 5897 45685 5983 45741
rect 6039 45685 6125 45741
rect 6181 45685 6267 45741
rect 6323 45685 6409 45741
rect 6465 45685 6551 45741
rect 6607 45685 6693 45741
rect 6749 45685 6835 45741
rect 6891 45685 6977 45741
rect 7033 45685 7119 45741
rect 7175 45685 7261 45741
rect 7317 45685 7403 45741
rect 7459 45685 7545 45741
rect 7601 45685 7687 45741
rect 7743 45685 7829 45741
rect 7885 45685 7971 45741
rect 8027 45685 8113 45741
rect 8169 45685 8255 45741
rect 8311 45685 8397 45741
rect 8453 45685 8539 45741
rect 8595 45685 8681 45741
rect 8737 45685 8823 45741
rect 8879 45685 8965 45741
rect 9021 45685 9107 45741
rect 9163 45685 9249 45741
rect 9305 45685 9391 45741
rect 9447 45685 9533 45741
rect 9589 45685 9675 45741
rect 9731 45685 9817 45741
rect 9873 45685 9959 45741
rect 10015 45685 10101 45741
rect 10157 45685 10243 45741
rect 10299 45685 10385 45741
rect 10441 45685 10527 45741
rect 10583 45685 10669 45741
rect 10725 45685 10811 45741
rect 10867 45685 10953 45741
rect 11009 45685 11095 45741
rect 11151 45685 11237 45741
rect 11293 45685 11379 45741
rect 11435 45685 11521 45741
rect 11577 45685 11663 45741
rect 11719 45685 11805 45741
rect 11861 45685 11947 45741
rect 12003 45685 12089 45741
rect 12145 45685 12231 45741
rect 12287 45685 12373 45741
rect 12429 45685 12515 45741
rect 12571 45685 12657 45741
rect 12713 45685 12799 45741
rect 12855 45685 12941 45741
rect 12997 45685 13083 45741
rect 13139 45685 13225 45741
rect 13281 45685 13367 45741
rect 13423 45685 13509 45741
rect 13565 45685 13651 45741
rect 13707 45685 13793 45741
rect 13849 45685 13935 45741
rect 13991 45685 14077 45741
rect 14133 45685 14219 45741
rect 14275 45685 14361 45741
rect 14417 45685 14503 45741
rect 14559 45685 14645 45741
rect 14701 45685 14787 45741
rect 14843 45685 14853 45741
rect 151 45599 14853 45685
rect 151 45543 161 45599
rect 217 45543 303 45599
rect 359 45543 445 45599
rect 501 45543 587 45599
rect 643 45543 729 45599
rect 785 45543 871 45599
rect 927 45543 1013 45599
rect 1069 45543 1155 45599
rect 1211 45543 1297 45599
rect 1353 45543 1439 45599
rect 1495 45543 1581 45599
rect 1637 45543 1723 45599
rect 1779 45543 1865 45599
rect 1921 45543 2007 45599
rect 2063 45543 2149 45599
rect 2205 45543 2291 45599
rect 2347 45543 2433 45599
rect 2489 45543 2575 45599
rect 2631 45543 2717 45599
rect 2773 45543 2859 45599
rect 2915 45543 3001 45599
rect 3057 45543 3143 45599
rect 3199 45543 3285 45599
rect 3341 45543 3427 45599
rect 3483 45543 3569 45599
rect 3625 45543 3711 45599
rect 3767 45543 3853 45599
rect 3909 45543 3995 45599
rect 4051 45543 4137 45599
rect 4193 45543 4279 45599
rect 4335 45543 4421 45599
rect 4477 45543 4563 45599
rect 4619 45543 4705 45599
rect 4761 45543 4847 45599
rect 4903 45543 4989 45599
rect 5045 45543 5131 45599
rect 5187 45543 5273 45599
rect 5329 45543 5415 45599
rect 5471 45543 5557 45599
rect 5613 45543 5699 45599
rect 5755 45543 5841 45599
rect 5897 45543 5983 45599
rect 6039 45543 6125 45599
rect 6181 45543 6267 45599
rect 6323 45543 6409 45599
rect 6465 45543 6551 45599
rect 6607 45543 6693 45599
rect 6749 45543 6835 45599
rect 6891 45543 6977 45599
rect 7033 45543 7119 45599
rect 7175 45543 7261 45599
rect 7317 45543 7403 45599
rect 7459 45543 7545 45599
rect 7601 45543 7687 45599
rect 7743 45543 7829 45599
rect 7885 45543 7971 45599
rect 8027 45543 8113 45599
rect 8169 45543 8255 45599
rect 8311 45543 8397 45599
rect 8453 45543 8539 45599
rect 8595 45543 8681 45599
rect 8737 45543 8823 45599
rect 8879 45543 8965 45599
rect 9021 45543 9107 45599
rect 9163 45543 9249 45599
rect 9305 45543 9391 45599
rect 9447 45543 9533 45599
rect 9589 45543 9675 45599
rect 9731 45543 9817 45599
rect 9873 45543 9959 45599
rect 10015 45543 10101 45599
rect 10157 45543 10243 45599
rect 10299 45543 10385 45599
rect 10441 45543 10527 45599
rect 10583 45543 10669 45599
rect 10725 45543 10811 45599
rect 10867 45543 10953 45599
rect 11009 45543 11095 45599
rect 11151 45543 11237 45599
rect 11293 45543 11379 45599
rect 11435 45543 11521 45599
rect 11577 45543 11663 45599
rect 11719 45543 11805 45599
rect 11861 45543 11947 45599
rect 12003 45543 12089 45599
rect 12145 45543 12231 45599
rect 12287 45543 12373 45599
rect 12429 45543 12515 45599
rect 12571 45543 12657 45599
rect 12713 45543 12799 45599
rect 12855 45543 12941 45599
rect 12997 45543 13083 45599
rect 13139 45543 13225 45599
rect 13281 45543 13367 45599
rect 13423 45543 13509 45599
rect 13565 45543 13651 45599
rect 13707 45543 13793 45599
rect 13849 45543 13935 45599
rect 13991 45543 14077 45599
rect 14133 45543 14219 45599
rect 14275 45543 14361 45599
rect 14417 45543 14503 45599
rect 14559 45543 14645 45599
rect 14701 45543 14787 45599
rect 14843 45543 14853 45599
rect 151 45457 14853 45543
rect 151 45401 161 45457
rect 217 45401 303 45457
rect 359 45401 445 45457
rect 501 45401 587 45457
rect 643 45401 729 45457
rect 785 45401 871 45457
rect 927 45401 1013 45457
rect 1069 45401 1155 45457
rect 1211 45401 1297 45457
rect 1353 45401 1439 45457
rect 1495 45401 1581 45457
rect 1637 45401 1723 45457
rect 1779 45401 1865 45457
rect 1921 45401 2007 45457
rect 2063 45401 2149 45457
rect 2205 45401 2291 45457
rect 2347 45401 2433 45457
rect 2489 45401 2575 45457
rect 2631 45401 2717 45457
rect 2773 45401 2859 45457
rect 2915 45401 3001 45457
rect 3057 45401 3143 45457
rect 3199 45401 3285 45457
rect 3341 45401 3427 45457
rect 3483 45401 3569 45457
rect 3625 45401 3711 45457
rect 3767 45401 3853 45457
rect 3909 45401 3995 45457
rect 4051 45401 4137 45457
rect 4193 45401 4279 45457
rect 4335 45401 4421 45457
rect 4477 45401 4563 45457
rect 4619 45401 4705 45457
rect 4761 45401 4847 45457
rect 4903 45401 4989 45457
rect 5045 45401 5131 45457
rect 5187 45401 5273 45457
rect 5329 45401 5415 45457
rect 5471 45401 5557 45457
rect 5613 45401 5699 45457
rect 5755 45401 5841 45457
rect 5897 45401 5983 45457
rect 6039 45401 6125 45457
rect 6181 45401 6267 45457
rect 6323 45401 6409 45457
rect 6465 45401 6551 45457
rect 6607 45401 6693 45457
rect 6749 45401 6835 45457
rect 6891 45401 6977 45457
rect 7033 45401 7119 45457
rect 7175 45401 7261 45457
rect 7317 45401 7403 45457
rect 7459 45401 7545 45457
rect 7601 45401 7687 45457
rect 7743 45401 7829 45457
rect 7885 45401 7971 45457
rect 8027 45401 8113 45457
rect 8169 45401 8255 45457
rect 8311 45401 8397 45457
rect 8453 45401 8539 45457
rect 8595 45401 8681 45457
rect 8737 45401 8823 45457
rect 8879 45401 8965 45457
rect 9021 45401 9107 45457
rect 9163 45401 9249 45457
rect 9305 45401 9391 45457
rect 9447 45401 9533 45457
rect 9589 45401 9675 45457
rect 9731 45401 9817 45457
rect 9873 45401 9959 45457
rect 10015 45401 10101 45457
rect 10157 45401 10243 45457
rect 10299 45401 10385 45457
rect 10441 45401 10527 45457
rect 10583 45401 10669 45457
rect 10725 45401 10811 45457
rect 10867 45401 10953 45457
rect 11009 45401 11095 45457
rect 11151 45401 11237 45457
rect 11293 45401 11379 45457
rect 11435 45401 11521 45457
rect 11577 45401 11663 45457
rect 11719 45401 11805 45457
rect 11861 45401 11947 45457
rect 12003 45401 12089 45457
rect 12145 45401 12231 45457
rect 12287 45401 12373 45457
rect 12429 45401 12515 45457
rect 12571 45401 12657 45457
rect 12713 45401 12799 45457
rect 12855 45401 12941 45457
rect 12997 45401 13083 45457
rect 13139 45401 13225 45457
rect 13281 45401 13367 45457
rect 13423 45401 13509 45457
rect 13565 45401 13651 45457
rect 13707 45401 13793 45457
rect 13849 45401 13935 45457
rect 13991 45401 14077 45457
rect 14133 45401 14219 45457
rect 14275 45401 14361 45457
rect 14417 45401 14503 45457
rect 14559 45401 14645 45457
rect 14701 45401 14787 45457
rect 14843 45401 14853 45457
rect 151 45315 14853 45401
rect 151 45259 161 45315
rect 217 45259 303 45315
rect 359 45259 445 45315
rect 501 45259 587 45315
rect 643 45259 729 45315
rect 785 45259 871 45315
rect 927 45259 1013 45315
rect 1069 45259 1155 45315
rect 1211 45259 1297 45315
rect 1353 45259 1439 45315
rect 1495 45259 1581 45315
rect 1637 45259 1723 45315
rect 1779 45259 1865 45315
rect 1921 45259 2007 45315
rect 2063 45259 2149 45315
rect 2205 45259 2291 45315
rect 2347 45259 2433 45315
rect 2489 45259 2575 45315
rect 2631 45259 2717 45315
rect 2773 45259 2859 45315
rect 2915 45259 3001 45315
rect 3057 45259 3143 45315
rect 3199 45259 3285 45315
rect 3341 45259 3427 45315
rect 3483 45259 3569 45315
rect 3625 45259 3711 45315
rect 3767 45259 3853 45315
rect 3909 45259 3995 45315
rect 4051 45259 4137 45315
rect 4193 45259 4279 45315
rect 4335 45259 4421 45315
rect 4477 45259 4563 45315
rect 4619 45259 4705 45315
rect 4761 45259 4847 45315
rect 4903 45259 4989 45315
rect 5045 45259 5131 45315
rect 5187 45259 5273 45315
rect 5329 45259 5415 45315
rect 5471 45259 5557 45315
rect 5613 45259 5699 45315
rect 5755 45259 5841 45315
rect 5897 45259 5983 45315
rect 6039 45259 6125 45315
rect 6181 45259 6267 45315
rect 6323 45259 6409 45315
rect 6465 45259 6551 45315
rect 6607 45259 6693 45315
rect 6749 45259 6835 45315
rect 6891 45259 6977 45315
rect 7033 45259 7119 45315
rect 7175 45259 7261 45315
rect 7317 45259 7403 45315
rect 7459 45259 7545 45315
rect 7601 45259 7687 45315
rect 7743 45259 7829 45315
rect 7885 45259 7971 45315
rect 8027 45259 8113 45315
rect 8169 45259 8255 45315
rect 8311 45259 8397 45315
rect 8453 45259 8539 45315
rect 8595 45259 8681 45315
rect 8737 45259 8823 45315
rect 8879 45259 8965 45315
rect 9021 45259 9107 45315
rect 9163 45259 9249 45315
rect 9305 45259 9391 45315
rect 9447 45259 9533 45315
rect 9589 45259 9675 45315
rect 9731 45259 9817 45315
rect 9873 45259 9959 45315
rect 10015 45259 10101 45315
rect 10157 45259 10243 45315
rect 10299 45259 10385 45315
rect 10441 45259 10527 45315
rect 10583 45259 10669 45315
rect 10725 45259 10811 45315
rect 10867 45259 10953 45315
rect 11009 45259 11095 45315
rect 11151 45259 11237 45315
rect 11293 45259 11379 45315
rect 11435 45259 11521 45315
rect 11577 45259 11663 45315
rect 11719 45259 11805 45315
rect 11861 45259 11947 45315
rect 12003 45259 12089 45315
rect 12145 45259 12231 45315
rect 12287 45259 12373 45315
rect 12429 45259 12515 45315
rect 12571 45259 12657 45315
rect 12713 45259 12799 45315
rect 12855 45259 12941 45315
rect 12997 45259 13083 45315
rect 13139 45259 13225 45315
rect 13281 45259 13367 45315
rect 13423 45259 13509 45315
rect 13565 45259 13651 45315
rect 13707 45259 13793 45315
rect 13849 45259 13935 45315
rect 13991 45259 14077 45315
rect 14133 45259 14219 45315
rect 14275 45259 14361 45315
rect 14417 45259 14503 45315
rect 14559 45259 14645 45315
rect 14701 45259 14787 45315
rect 14843 45259 14853 45315
rect 151 45173 14853 45259
rect 151 45117 161 45173
rect 217 45117 303 45173
rect 359 45117 445 45173
rect 501 45117 587 45173
rect 643 45117 729 45173
rect 785 45117 871 45173
rect 927 45117 1013 45173
rect 1069 45117 1155 45173
rect 1211 45117 1297 45173
rect 1353 45117 1439 45173
rect 1495 45117 1581 45173
rect 1637 45117 1723 45173
rect 1779 45117 1865 45173
rect 1921 45117 2007 45173
rect 2063 45117 2149 45173
rect 2205 45117 2291 45173
rect 2347 45117 2433 45173
rect 2489 45117 2575 45173
rect 2631 45117 2717 45173
rect 2773 45117 2859 45173
rect 2915 45117 3001 45173
rect 3057 45117 3143 45173
rect 3199 45117 3285 45173
rect 3341 45117 3427 45173
rect 3483 45117 3569 45173
rect 3625 45117 3711 45173
rect 3767 45117 3853 45173
rect 3909 45117 3995 45173
rect 4051 45117 4137 45173
rect 4193 45117 4279 45173
rect 4335 45117 4421 45173
rect 4477 45117 4563 45173
rect 4619 45117 4705 45173
rect 4761 45117 4847 45173
rect 4903 45117 4989 45173
rect 5045 45117 5131 45173
rect 5187 45117 5273 45173
rect 5329 45117 5415 45173
rect 5471 45117 5557 45173
rect 5613 45117 5699 45173
rect 5755 45117 5841 45173
rect 5897 45117 5983 45173
rect 6039 45117 6125 45173
rect 6181 45117 6267 45173
rect 6323 45117 6409 45173
rect 6465 45117 6551 45173
rect 6607 45117 6693 45173
rect 6749 45117 6835 45173
rect 6891 45117 6977 45173
rect 7033 45117 7119 45173
rect 7175 45117 7261 45173
rect 7317 45117 7403 45173
rect 7459 45117 7545 45173
rect 7601 45117 7687 45173
rect 7743 45117 7829 45173
rect 7885 45117 7971 45173
rect 8027 45117 8113 45173
rect 8169 45117 8255 45173
rect 8311 45117 8397 45173
rect 8453 45117 8539 45173
rect 8595 45117 8681 45173
rect 8737 45117 8823 45173
rect 8879 45117 8965 45173
rect 9021 45117 9107 45173
rect 9163 45117 9249 45173
rect 9305 45117 9391 45173
rect 9447 45117 9533 45173
rect 9589 45117 9675 45173
rect 9731 45117 9817 45173
rect 9873 45117 9959 45173
rect 10015 45117 10101 45173
rect 10157 45117 10243 45173
rect 10299 45117 10385 45173
rect 10441 45117 10527 45173
rect 10583 45117 10669 45173
rect 10725 45117 10811 45173
rect 10867 45117 10953 45173
rect 11009 45117 11095 45173
rect 11151 45117 11237 45173
rect 11293 45117 11379 45173
rect 11435 45117 11521 45173
rect 11577 45117 11663 45173
rect 11719 45117 11805 45173
rect 11861 45117 11947 45173
rect 12003 45117 12089 45173
rect 12145 45117 12231 45173
rect 12287 45117 12373 45173
rect 12429 45117 12515 45173
rect 12571 45117 12657 45173
rect 12713 45117 12799 45173
rect 12855 45117 12941 45173
rect 12997 45117 13083 45173
rect 13139 45117 13225 45173
rect 13281 45117 13367 45173
rect 13423 45117 13509 45173
rect 13565 45117 13651 45173
rect 13707 45117 13793 45173
rect 13849 45117 13935 45173
rect 13991 45117 14077 45173
rect 14133 45117 14219 45173
rect 14275 45117 14361 45173
rect 14417 45117 14503 45173
rect 14559 45117 14645 45173
rect 14701 45117 14787 45173
rect 14843 45117 14853 45173
rect 151 45031 14853 45117
rect 151 44975 161 45031
rect 217 44975 303 45031
rect 359 44975 445 45031
rect 501 44975 587 45031
rect 643 44975 729 45031
rect 785 44975 871 45031
rect 927 44975 1013 45031
rect 1069 44975 1155 45031
rect 1211 44975 1297 45031
rect 1353 44975 1439 45031
rect 1495 44975 1581 45031
rect 1637 44975 1723 45031
rect 1779 44975 1865 45031
rect 1921 44975 2007 45031
rect 2063 44975 2149 45031
rect 2205 44975 2291 45031
rect 2347 44975 2433 45031
rect 2489 44975 2575 45031
rect 2631 44975 2717 45031
rect 2773 44975 2859 45031
rect 2915 44975 3001 45031
rect 3057 44975 3143 45031
rect 3199 44975 3285 45031
rect 3341 44975 3427 45031
rect 3483 44975 3569 45031
rect 3625 44975 3711 45031
rect 3767 44975 3853 45031
rect 3909 44975 3995 45031
rect 4051 44975 4137 45031
rect 4193 44975 4279 45031
rect 4335 44975 4421 45031
rect 4477 44975 4563 45031
rect 4619 44975 4705 45031
rect 4761 44975 4847 45031
rect 4903 44975 4989 45031
rect 5045 44975 5131 45031
rect 5187 44975 5273 45031
rect 5329 44975 5415 45031
rect 5471 44975 5557 45031
rect 5613 44975 5699 45031
rect 5755 44975 5841 45031
rect 5897 44975 5983 45031
rect 6039 44975 6125 45031
rect 6181 44975 6267 45031
rect 6323 44975 6409 45031
rect 6465 44975 6551 45031
rect 6607 44975 6693 45031
rect 6749 44975 6835 45031
rect 6891 44975 6977 45031
rect 7033 44975 7119 45031
rect 7175 44975 7261 45031
rect 7317 44975 7403 45031
rect 7459 44975 7545 45031
rect 7601 44975 7687 45031
rect 7743 44975 7829 45031
rect 7885 44975 7971 45031
rect 8027 44975 8113 45031
rect 8169 44975 8255 45031
rect 8311 44975 8397 45031
rect 8453 44975 8539 45031
rect 8595 44975 8681 45031
rect 8737 44975 8823 45031
rect 8879 44975 8965 45031
rect 9021 44975 9107 45031
rect 9163 44975 9249 45031
rect 9305 44975 9391 45031
rect 9447 44975 9533 45031
rect 9589 44975 9675 45031
rect 9731 44975 9817 45031
rect 9873 44975 9959 45031
rect 10015 44975 10101 45031
rect 10157 44975 10243 45031
rect 10299 44975 10385 45031
rect 10441 44975 10527 45031
rect 10583 44975 10669 45031
rect 10725 44975 10811 45031
rect 10867 44975 10953 45031
rect 11009 44975 11095 45031
rect 11151 44975 11237 45031
rect 11293 44975 11379 45031
rect 11435 44975 11521 45031
rect 11577 44975 11663 45031
rect 11719 44975 11805 45031
rect 11861 44975 11947 45031
rect 12003 44975 12089 45031
rect 12145 44975 12231 45031
rect 12287 44975 12373 45031
rect 12429 44975 12515 45031
rect 12571 44975 12657 45031
rect 12713 44975 12799 45031
rect 12855 44975 12941 45031
rect 12997 44975 13083 45031
rect 13139 44975 13225 45031
rect 13281 44975 13367 45031
rect 13423 44975 13509 45031
rect 13565 44975 13651 45031
rect 13707 44975 13793 45031
rect 13849 44975 13935 45031
rect 13991 44975 14077 45031
rect 14133 44975 14219 45031
rect 14275 44975 14361 45031
rect 14417 44975 14503 45031
rect 14559 44975 14645 45031
rect 14701 44975 14787 45031
rect 14843 44975 14853 45031
rect 151 44889 14853 44975
rect 151 44833 161 44889
rect 217 44833 303 44889
rect 359 44833 445 44889
rect 501 44833 587 44889
rect 643 44833 729 44889
rect 785 44833 871 44889
rect 927 44833 1013 44889
rect 1069 44833 1155 44889
rect 1211 44833 1297 44889
rect 1353 44833 1439 44889
rect 1495 44833 1581 44889
rect 1637 44833 1723 44889
rect 1779 44833 1865 44889
rect 1921 44833 2007 44889
rect 2063 44833 2149 44889
rect 2205 44833 2291 44889
rect 2347 44833 2433 44889
rect 2489 44833 2575 44889
rect 2631 44833 2717 44889
rect 2773 44833 2859 44889
rect 2915 44833 3001 44889
rect 3057 44833 3143 44889
rect 3199 44833 3285 44889
rect 3341 44833 3427 44889
rect 3483 44833 3569 44889
rect 3625 44833 3711 44889
rect 3767 44833 3853 44889
rect 3909 44833 3995 44889
rect 4051 44833 4137 44889
rect 4193 44833 4279 44889
rect 4335 44833 4421 44889
rect 4477 44833 4563 44889
rect 4619 44833 4705 44889
rect 4761 44833 4847 44889
rect 4903 44833 4989 44889
rect 5045 44833 5131 44889
rect 5187 44833 5273 44889
rect 5329 44833 5415 44889
rect 5471 44833 5557 44889
rect 5613 44833 5699 44889
rect 5755 44833 5841 44889
rect 5897 44833 5983 44889
rect 6039 44833 6125 44889
rect 6181 44833 6267 44889
rect 6323 44833 6409 44889
rect 6465 44833 6551 44889
rect 6607 44833 6693 44889
rect 6749 44833 6835 44889
rect 6891 44833 6977 44889
rect 7033 44833 7119 44889
rect 7175 44833 7261 44889
rect 7317 44833 7403 44889
rect 7459 44833 7545 44889
rect 7601 44833 7687 44889
rect 7743 44833 7829 44889
rect 7885 44833 7971 44889
rect 8027 44833 8113 44889
rect 8169 44833 8255 44889
rect 8311 44833 8397 44889
rect 8453 44833 8539 44889
rect 8595 44833 8681 44889
rect 8737 44833 8823 44889
rect 8879 44833 8965 44889
rect 9021 44833 9107 44889
rect 9163 44833 9249 44889
rect 9305 44833 9391 44889
rect 9447 44833 9533 44889
rect 9589 44833 9675 44889
rect 9731 44833 9817 44889
rect 9873 44833 9959 44889
rect 10015 44833 10101 44889
rect 10157 44833 10243 44889
rect 10299 44833 10385 44889
rect 10441 44833 10527 44889
rect 10583 44833 10669 44889
rect 10725 44833 10811 44889
rect 10867 44833 10953 44889
rect 11009 44833 11095 44889
rect 11151 44833 11237 44889
rect 11293 44833 11379 44889
rect 11435 44833 11521 44889
rect 11577 44833 11663 44889
rect 11719 44833 11805 44889
rect 11861 44833 11947 44889
rect 12003 44833 12089 44889
rect 12145 44833 12231 44889
rect 12287 44833 12373 44889
rect 12429 44833 12515 44889
rect 12571 44833 12657 44889
rect 12713 44833 12799 44889
rect 12855 44833 12941 44889
rect 12997 44833 13083 44889
rect 13139 44833 13225 44889
rect 13281 44833 13367 44889
rect 13423 44833 13509 44889
rect 13565 44833 13651 44889
rect 13707 44833 13793 44889
rect 13849 44833 13935 44889
rect 13991 44833 14077 44889
rect 14133 44833 14219 44889
rect 14275 44833 14361 44889
rect 14417 44833 14503 44889
rect 14559 44833 14645 44889
rect 14701 44833 14787 44889
rect 14843 44833 14853 44889
rect 151 44747 14853 44833
rect 151 44691 161 44747
rect 217 44691 303 44747
rect 359 44691 445 44747
rect 501 44691 587 44747
rect 643 44691 729 44747
rect 785 44691 871 44747
rect 927 44691 1013 44747
rect 1069 44691 1155 44747
rect 1211 44691 1297 44747
rect 1353 44691 1439 44747
rect 1495 44691 1581 44747
rect 1637 44691 1723 44747
rect 1779 44691 1865 44747
rect 1921 44691 2007 44747
rect 2063 44691 2149 44747
rect 2205 44691 2291 44747
rect 2347 44691 2433 44747
rect 2489 44691 2575 44747
rect 2631 44691 2717 44747
rect 2773 44691 2859 44747
rect 2915 44691 3001 44747
rect 3057 44691 3143 44747
rect 3199 44691 3285 44747
rect 3341 44691 3427 44747
rect 3483 44691 3569 44747
rect 3625 44691 3711 44747
rect 3767 44691 3853 44747
rect 3909 44691 3995 44747
rect 4051 44691 4137 44747
rect 4193 44691 4279 44747
rect 4335 44691 4421 44747
rect 4477 44691 4563 44747
rect 4619 44691 4705 44747
rect 4761 44691 4847 44747
rect 4903 44691 4989 44747
rect 5045 44691 5131 44747
rect 5187 44691 5273 44747
rect 5329 44691 5415 44747
rect 5471 44691 5557 44747
rect 5613 44691 5699 44747
rect 5755 44691 5841 44747
rect 5897 44691 5983 44747
rect 6039 44691 6125 44747
rect 6181 44691 6267 44747
rect 6323 44691 6409 44747
rect 6465 44691 6551 44747
rect 6607 44691 6693 44747
rect 6749 44691 6835 44747
rect 6891 44691 6977 44747
rect 7033 44691 7119 44747
rect 7175 44691 7261 44747
rect 7317 44691 7403 44747
rect 7459 44691 7545 44747
rect 7601 44691 7687 44747
rect 7743 44691 7829 44747
rect 7885 44691 7971 44747
rect 8027 44691 8113 44747
rect 8169 44691 8255 44747
rect 8311 44691 8397 44747
rect 8453 44691 8539 44747
rect 8595 44691 8681 44747
rect 8737 44691 8823 44747
rect 8879 44691 8965 44747
rect 9021 44691 9107 44747
rect 9163 44691 9249 44747
rect 9305 44691 9391 44747
rect 9447 44691 9533 44747
rect 9589 44691 9675 44747
rect 9731 44691 9817 44747
rect 9873 44691 9959 44747
rect 10015 44691 10101 44747
rect 10157 44691 10243 44747
rect 10299 44691 10385 44747
rect 10441 44691 10527 44747
rect 10583 44691 10669 44747
rect 10725 44691 10811 44747
rect 10867 44691 10953 44747
rect 11009 44691 11095 44747
rect 11151 44691 11237 44747
rect 11293 44691 11379 44747
rect 11435 44691 11521 44747
rect 11577 44691 11663 44747
rect 11719 44691 11805 44747
rect 11861 44691 11947 44747
rect 12003 44691 12089 44747
rect 12145 44691 12231 44747
rect 12287 44691 12373 44747
rect 12429 44691 12515 44747
rect 12571 44691 12657 44747
rect 12713 44691 12799 44747
rect 12855 44691 12941 44747
rect 12997 44691 13083 44747
rect 13139 44691 13225 44747
rect 13281 44691 13367 44747
rect 13423 44691 13509 44747
rect 13565 44691 13651 44747
rect 13707 44691 13793 44747
rect 13849 44691 13935 44747
rect 13991 44691 14077 44747
rect 14133 44691 14219 44747
rect 14275 44691 14361 44747
rect 14417 44691 14503 44747
rect 14559 44691 14645 44747
rect 14701 44691 14787 44747
rect 14843 44691 14853 44747
rect 151 44605 14853 44691
rect 151 44549 161 44605
rect 217 44549 303 44605
rect 359 44549 445 44605
rect 501 44549 587 44605
rect 643 44549 729 44605
rect 785 44549 871 44605
rect 927 44549 1013 44605
rect 1069 44549 1155 44605
rect 1211 44549 1297 44605
rect 1353 44549 1439 44605
rect 1495 44549 1581 44605
rect 1637 44549 1723 44605
rect 1779 44549 1865 44605
rect 1921 44549 2007 44605
rect 2063 44549 2149 44605
rect 2205 44549 2291 44605
rect 2347 44549 2433 44605
rect 2489 44549 2575 44605
rect 2631 44549 2717 44605
rect 2773 44549 2859 44605
rect 2915 44549 3001 44605
rect 3057 44549 3143 44605
rect 3199 44549 3285 44605
rect 3341 44549 3427 44605
rect 3483 44549 3569 44605
rect 3625 44549 3711 44605
rect 3767 44549 3853 44605
rect 3909 44549 3995 44605
rect 4051 44549 4137 44605
rect 4193 44549 4279 44605
rect 4335 44549 4421 44605
rect 4477 44549 4563 44605
rect 4619 44549 4705 44605
rect 4761 44549 4847 44605
rect 4903 44549 4989 44605
rect 5045 44549 5131 44605
rect 5187 44549 5273 44605
rect 5329 44549 5415 44605
rect 5471 44549 5557 44605
rect 5613 44549 5699 44605
rect 5755 44549 5841 44605
rect 5897 44549 5983 44605
rect 6039 44549 6125 44605
rect 6181 44549 6267 44605
rect 6323 44549 6409 44605
rect 6465 44549 6551 44605
rect 6607 44549 6693 44605
rect 6749 44549 6835 44605
rect 6891 44549 6977 44605
rect 7033 44549 7119 44605
rect 7175 44549 7261 44605
rect 7317 44549 7403 44605
rect 7459 44549 7545 44605
rect 7601 44549 7687 44605
rect 7743 44549 7829 44605
rect 7885 44549 7971 44605
rect 8027 44549 8113 44605
rect 8169 44549 8255 44605
rect 8311 44549 8397 44605
rect 8453 44549 8539 44605
rect 8595 44549 8681 44605
rect 8737 44549 8823 44605
rect 8879 44549 8965 44605
rect 9021 44549 9107 44605
rect 9163 44549 9249 44605
rect 9305 44549 9391 44605
rect 9447 44549 9533 44605
rect 9589 44549 9675 44605
rect 9731 44549 9817 44605
rect 9873 44549 9959 44605
rect 10015 44549 10101 44605
rect 10157 44549 10243 44605
rect 10299 44549 10385 44605
rect 10441 44549 10527 44605
rect 10583 44549 10669 44605
rect 10725 44549 10811 44605
rect 10867 44549 10953 44605
rect 11009 44549 11095 44605
rect 11151 44549 11237 44605
rect 11293 44549 11379 44605
rect 11435 44549 11521 44605
rect 11577 44549 11663 44605
rect 11719 44549 11805 44605
rect 11861 44549 11947 44605
rect 12003 44549 12089 44605
rect 12145 44549 12231 44605
rect 12287 44549 12373 44605
rect 12429 44549 12515 44605
rect 12571 44549 12657 44605
rect 12713 44549 12799 44605
rect 12855 44549 12941 44605
rect 12997 44549 13083 44605
rect 13139 44549 13225 44605
rect 13281 44549 13367 44605
rect 13423 44549 13509 44605
rect 13565 44549 13651 44605
rect 13707 44549 13793 44605
rect 13849 44549 13935 44605
rect 13991 44549 14077 44605
rect 14133 44549 14219 44605
rect 14275 44549 14361 44605
rect 14417 44549 14503 44605
rect 14559 44549 14645 44605
rect 14701 44549 14787 44605
rect 14843 44549 14853 44605
rect 151 44463 14853 44549
rect 151 44407 161 44463
rect 217 44407 303 44463
rect 359 44407 445 44463
rect 501 44407 587 44463
rect 643 44407 729 44463
rect 785 44407 871 44463
rect 927 44407 1013 44463
rect 1069 44407 1155 44463
rect 1211 44407 1297 44463
rect 1353 44407 1439 44463
rect 1495 44407 1581 44463
rect 1637 44407 1723 44463
rect 1779 44407 1865 44463
rect 1921 44407 2007 44463
rect 2063 44407 2149 44463
rect 2205 44407 2291 44463
rect 2347 44407 2433 44463
rect 2489 44407 2575 44463
rect 2631 44407 2717 44463
rect 2773 44407 2859 44463
rect 2915 44407 3001 44463
rect 3057 44407 3143 44463
rect 3199 44407 3285 44463
rect 3341 44407 3427 44463
rect 3483 44407 3569 44463
rect 3625 44407 3711 44463
rect 3767 44407 3853 44463
rect 3909 44407 3995 44463
rect 4051 44407 4137 44463
rect 4193 44407 4279 44463
rect 4335 44407 4421 44463
rect 4477 44407 4563 44463
rect 4619 44407 4705 44463
rect 4761 44407 4847 44463
rect 4903 44407 4989 44463
rect 5045 44407 5131 44463
rect 5187 44407 5273 44463
rect 5329 44407 5415 44463
rect 5471 44407 5557 44463
rect 5613 44407 5699 44463
rect 5755 44407 5841 44463
rect 5897 44407 5983 44463
rect 6039 44407 6125 44463
rect 6181 44407 6267 44463
rect 6323 44407 6409 44463
rect 6465 44407 6551 44463
rect 6607 44407 6693 44463
rect 6749 44407 6835 44463
rect 6891 44407 6977 44463
rect 7033 44407 7119 44463
rect 7175 44407 7261 44463
rect 7317 44407 7403 44463
rect 7459 44407 7545 44463
rect 7601 44407 7687 44463
rect 7743 44407 7829 44463
rect 7885 44407 7971 44463
rect 8027 44407 8113 44463
rect 8169 44407 8255 44463
rect 8311 44407 8397 44463
rect 8453 44407 8539 44463
rect 8595 44407 8681 44463
rect 8737 44407 8823 44463
rect 8879 44407 8965 44463
rect 9021 44407 9107 44463
rect 9163 44407 9249 44463
rect 9305 44407 9391 44463
rect 9447 44407 9533 44463
rect 9589 44407 9675 44463
rect 9731 44407 9817 44463
rect 9873 44407 9959 44463
rect 10015 44407 10101 44463
rect 10157 44407 10243 44463
rect 10299 44407 10385 44463
rect 10441 44407 10527 44463
rect 10583 44407 10669 44463
rect 10725 44407 10811 44463
rect 10867 44407 10953 44463
rect 11009 44407 11095 44463
rect 11151 44407 11237 44463
rect 11293 44407 11379 44463
rect 11435 44407 11521 44463
rect 11577 44407 11663 44463
rect 11719 44407 11805 44463
rect 11861 44407 11947 44463
rect 12003 44407 12089 44463
rect 12145 44407 12231 44463
rect 12287 44407 12373 44463
rect 12429 44407 12515 44463
rect 12571 44407 12657 44463
rect 12713 44407 12799 44463
rect 12855 44407 12941 44463
rect 12997 44407 13083 44463
rect 13139 44407 13225 44463
rect 13281 44407 13367 44463
rect 13423 44407 13509 44463
rect 13565 44407 13651 44463
rect 13707 44407 13793 44463
rect 13849 44407 13935 44463
rect 13991 44407 14077 44463
rect 14133 44407 14219 44463
rect 14275 44407 14361 44463
rect 14417 44407 14503 44463
rect 14559 44407 14645 44463
rect 14701 44407 14787 44463
rect 14843 44407 14853 44463
rect 151 44321 14853 44407
rect 151 44265 161 44321
rect 217 44265 303 44321
rect 359 44265 445 44321
rect 501 44265 587 44321
rect 643 44265 729 44321
rect 785 44265 871 44321
rect 927 44265 1013 44321
rect 1069 44265 1155 44321
rect 1211 44265 1297 44321
rect 1353 44265 1439 44321
rect 1495 44265 1581 44321
rect 1637 44265 1723 44321
rect 1779 44265 1865 44321
rect 1921 44265 2007 44321
rect 2063 44265 2149 44321
rect 2205 44265 2291 44321
rect 2347 44265 2433 44321
rect 2489 44265 2575 44321
rect 2631 44265 2717 44321
rect 2773 44265 2859 44321
rect 2915 44265 3001 44321
rect 3057 44265 3143 44321
rect 3199 44265 3285 44321
rect 3341 44265 3427 44321
rect 3483 44265 3569 44321
rect 3625 44265 3711 44321
rect 3767 44265 3853 44321
rect 3909 44265 3995 44321
rect 4051 44265 4137 44321
rect 4193 44265 4279 44321
rect 4335 44265 4421 44321
rect 4477 44265 4563 44321
rect 4619 44265 4705 44321
rect 4761 44265 4847 44321
rect 4903 44265 4989 44321
rect 5045 44265 5131 44321
rect 5187 44265 5273 44321
rect 5329 44265 5415 44321
rect 5471 44265 5557 44321
rect 5613 44265 5699 44321
rect 5755 44265 5841 44321
rect 5897 44265 5983 44321
rect 6039 44265 6125 44321
rect 6181 44265 6267 44321
rect 6323 44265 6409 44321
rect 6465 44265 6551 44321
rect 6607 44265 6693 44321
rect 6749 44265 6835 44321
rect 6891 44265 6977 44321
rect 7033 44265 7119 44321
rect 7175 44265 7261 44321
rect 7317 44265 7403 44321
rect 7459 44265 7545 44321
rect 7601 44265 7687 44321
rect 7743 44265 7829 44321
rect 7885 44265 7971 44321
rect 8027 44265 8113 44321
rect 8169 44265 8255 44321
rect 8311 44265 8397 44321
rect 8453 44265 8539 44321
rect 8595 44265 8681 44321
rect 8737 44265 8823 44321
rect 8879 44265 8965 44321
rect 9021 44265 9107 44321
rect 9163 44265 9249 44321
rect 9305 44265 9391 44321
rect 9447 44265 9533 44321
rect 9589 44265 9675 44321
rect 9731 44265 9817 44321
rect 9873 44265 9959 44321
rect 10015 44265 10101 44321
rect 10157 44265 10243 44321
rect 10299 44265 10385 44321
rect 10441 44265 10527 44321
rect 10583 44265 10669 44321
rect 10725 44265 10811 44321
rect 10867 44265 10953 44321
rect 11009 44265 11095 44321
rect 11151 44265 11237 44321
rect 11293 44265 11379 44321
rect 11435 44265 11521 44321
rect 11577 44265 11663 44321
rect 11719 44265 11805 44321
rect 11861 44265 11947 44321
rect 12003 44265 12089 44321
rect 12145 44265 12231 44321
rect 12287 44265 12373 44321
rect 12429 44265 12515 44321
rect 12571 44265 12657 44321
rect 12713 44265 12799 44321
rect 12855 44265 12941 44321
rect 12997 44265 13083 44321
rect 13139 44265 13225 44321
rect 13281 44265 13367 44321
rect 13423 44265 13509 44321
rect 13565 44265 13651 44321
rect 13707 44265 13793 44321
rect 13849 44265 13935 44321
rect 13991 44265 14077 44321
rect 14133 44265 14219 44321
rect 14275 44265 14361 44321
rect 14417 44265 14503 44321
rect 14559 44265 14645 44321
rect 14701 44265 14787 44321
rect 14843 44265 14853 44321
rect 151 44179 14853 44265
rect 151 44123 161 44179
rect 217 44123 303 44179
rect 359 44123 445 44179
rect 501 44123 587 44179
rect 643 44123 729 44179
rect 785 44123 871 44179
rect 927 44123 1013 44179
rect 1069 44123 1155 44179
rect 1211 44123 1297 44179
rect 1353 44123 1439 44179
rect 1495 44123 1581 44179
rect 1637 44123 1723 44179
rect 1779 44123 1865 44179
rect 1921 44123 2007 44179
rect 2063 44123 2149 44179
rect 2205 44123 2291 44179
rect 2347 44123 2433 44179
rect 2489 44123 2575 44179
rect 2631 44123 2717 44179
rect 2773 44123 2859 44179
rect 2915 44123 3001 44179
rect 3057 44123 3143 44179
rect 3199 44123 3285 44179
rect 3341 44123 3427 44179
rect 3483 44123 3569 44179
rect 3625 44123 3711 44179
rect 3767 44123 3853 44179
rect 3909 44123 3995 44179
rect 4051 44123 4137 44179
rect 4193 44123 4279 44179
rect 4335 44123 4421 44179
rect 4477 44123 4563 44179
rect 4619 44123 4705 44179
rect 4761 44123 4847 44179
rect 4903 44123 4989 44179
rect 5045 44123 5131 44179
rect 5187 44123 5273 44179
rect 5329 44123 5415 44179
rect 5471 44123 5557 44179
rect 5613 44123 5699 44179
rect 5755 44123 5841 44179
rect 5897 44123 5983 44179
rect 6039 44123 6125 44179
rect 6181 44123 6267 44179
rect 6323 44123 6409 44179
rect 6465 44123 6551 44179
rect 6607 44123 6693 44179
rect 6749 44123 6835 44179
rect 6891 44123 6977 44179
rect 7033 44123 7119 44179
rect 7175 44123 7261 44179
rect 7317 44123 7403 44179
rect 7459 44123 7545 44179
rect 7601 44123 7687 44179
rect 7743 44123 7829 44179
rect 7885 44123 7971 44179
rect 8027 44123 8113 44179
rect 8169 44123 8255 44179
rect 8311 44123 8397 44179
rect 8453 44123 8539 44179
rect 8595 44123 8681 44179
rect 8737 44123 8823 44179
rect 8879 44123 8965 44179
rect 9021 44123 9107 44179
rect 9163 44123 9249 44179
rect 9305 44123 9391 44179
rect 9447 44123 9533 44179
rect 9589 44123 9675 44179
rect 9731 44123 9817 44179
rect 9873 44123 9959 44179
rect 10015 44123 10101 44179
rect 10157 44123 10243 44179
rect 10299 44123 10385 44179
rect 10441 44123 10527 44179
rect 10583 44123 10669 44179
rect 10725 44123 10811 44179
rect 10867 44123 10953 44179
rect 11009 44123 11095 44179
rect 11151 44123 11237 44179
rect 11293 44123 11379 44179
rect 11435 44123 11521 44179
rect 11577 44123 11663 44179
rect 11719 44123 11805 44179
rect 11861 44123 11947 44179
rect 12003 44123 12089 44179
rect 12145 44123 12231 44179
rect 12287 44123 12373 44179
rect 12429 44123 12515 44179
rect 12571 44123 12657 44179
rect 12713 44123 12799 44179
rect 12855 44123 12941 44179
rect 12997 44123 13083 44179
rect 13139 44123 13225 44179
rect 13281 44123 13367 44179
rect 13423 44123 13509 44179
rect 13565 44123 13651 44179
rect 13707 44123 13793 44179
rect 13849 44123 13935 44179
rect 13991 44123 14077 44179
rect 14133 44123 14219 44179
rect 14275 44123 14361 44179
rect 14417 44123 14503 44179
rect 14559 44123 14645 44179
rect 14701 44123 14787 44179
rect 14843 44123 14853 44179
rect 151 44037 14853 44123
rect 151 43981 161 44037
rect 217 43981 303 44037
rect 359 43981 445 44037
rect 501 43981 587 44037
rect 643 43981 729 44037
rect 785 43981 871 44037
rect 927 43981 1013 44037
rect 1069 43981 1155 44037
rect 1211 43981 1297 44037
rect 1353 43981 1439 44037
rect 1495 43981 1581 44037
rect 1637 43981 1723 44037
rect 1779 43981 1865 44037
rect 1921 43981 2007 44037
rect 2063 43981 2149 44037
rect 2205 43981 2291 44037
rect 2347 43981 2433 44037
rect 2489 43981 2575 44037
rect 2631 43981 2717 44037
rect 2773 43981 2859 44037
rect 2915 43981 3001 44037
rect 3057 43981 3143 44037
rect 3199 43981 3285 44037
rect 3341 43981 3427 44037
rect 3483 43981 3569 44037
rect 3625 43981 3711 44037
rect 3767 43981 3853 44037
rect 3909 43981 3995 44037
rect 4051 43981 4137 44037
rect 4193 43981 4279 44037
rect 4335 43981 4421 44037
rect 4477 43981 4563 44037
rect 4619 43981 4705 44037
rect 4761 43981 4847 44037
rect 4903 43981 4989 44037
rect 5045 43981 5131 44037
rect 5187 43981 5273 44037
rect 5329 43981 5415 44037
rect 5471 43981 5557 44037
rect 5613 43981 5699 44037
rect 5755 43981 5841 44037
rect 5897 43981 5983 44037
rect 6039 43981 6125 44037
rect 6181 43981 6267 44037
rect 6323 43981 6409 44037
rect 6465 43981 6551 44037
rect 6607 43981 6693 44037
rect 6749 43981 6835 44037
rect 6891 43981 6977 44037
rect 7033 43981 7119 44037
rect 7175 43981 7261 44037
rect 7317 43981 7403 44037
rect 7459 43981 7545 44037
rect 7601 43981 7687 44037
rect 7743 43981 7829 44037
rect 7885 43981 7971 44037
rect 8027 43981 8113 44037
rect 8169 43981 8255 44037
rect 8311 43981 8397 44037
rect 8453 43981 8539 44037
rect 8595 43981 8681 44037
rect 8737 43981 8823 44037
rect 8879 43981 8965 44037
rect 9021 43981 9107 44037
rect 9163 43981 9249 44037
rect 9305 43981 9391 44037
rect 9447 43981 9533 44037
rect 9589 43981 9675 44037
rect 9731 43981 9817 44037
rect 9873 43981 9959 44037
rect 10015 43981 10101 44037
rect 10157 43981 10243 44037
rect 10299 43981 10385 44037
rect 10441 43981 10527 44037
rect 10583 43981 10669 44037
rect 10725 43981 10811 44037
rect 10867 43981 10953 44037
rect 11009 43981 11095 44037
rect 11151 43981 11237 44037
rect 11293 43981 11379 44037
rect 11435 43981 11521 44037
rect 11577 43981 11663 44037
rect 11719 43981 11805 44037
rect 11861 43981 11947 44037
rect 12003 43981 12089 44037
rect 12145 43981 12231 44037
rect 12287 43981 12373 44037
rect 12429 43981 12515 44037
rect 12571 43981 12657 44037
rect 12713 43981 12799 44037
rect 12855 43981 12941 44037
rect 12997 43981 13083 44037
rect 13139 43981 13225 44037
rect 13281 43981 13367 44037
rect 13423 43981 13509 44037
rect 13565 43981 13651 44037
rect 13707 43981 13793 44037
rect 13849 43981 13935 44037
rect 13991 43981 14077 44037
rect 14133 43981 14219 44037
rect 14275 43981 14361 44037
rect 14417 43981 14503 44037
rect 14559 43981 14645 44037
rect 14701 43981 14787 44037
rect 14843 43981 14853 44037
rect 151 43895 14853 43981
rect 151 43839 161 43895
rect 217 43839 303 43895
rect 359 43839 445 43895
rect 501 43839 587 43895
rect 643 43839 729 43895
rect 785 43839 871 43895
rect 927 43839 1013 43895
rect 1069 43839 1155 43895
rect 1211 43839 1297 43895
rect 1353 43839 1439 43895
rect 1495 43839 1581 43895
rect 1637 43839 1723 43895
rect 1779 43839 1865 43895
rect 1921 43839 2007 43895
rect 2063 43839 2149 43895
rect 2205 43839 2291 43895
rect 2347 43839 2433 43895
rect 2489 43839 2575 43895
rect 2631 43839 2717 43895
rect 2773 43839 2859 43895
rect 2915 43839 3001 43895
rect 3057 43839 3143 43895
rect 3199 43839 3285 43895
rect 3341 43839 3427 43895
rect 3483 43839 3569 43895
rect 3625 43839 3711 43895
rect 3767 43839 3853 43895
rect 3909 43839 3995 43895
rect 4051 43839 4137 43895
rect 4193 43839 4279 43895
rect 4335 43839 4421 43895
rect 4477 43839 4563 43895
rect 4619 43839 4705 43895
rect 4761 43839 4847 43895
rect 4903 43839 4989 43895
rect 5045 43839 5131 43895
rect 5187 43839 5273 43895
rect 5329 43839 5415 43895
rect 5471 43839 5557 43895
rect 5613 43839 5699 43895
rect 5755 43839 5841 43895
rect 5897 43839 5983 43895
rect 6039 43839 6125 43895
rect 6181 43839 6267 43895
rect 6323 43839 6409 43895
rect 6465 43839 6551 43895
rect 6607 43839 6693 43895
rect 6749 43839 6835 43895
rect 6891 43839 6977 43895
rect 7033 43839 7119 43895
rect 7175 43839 7261 43895
rect 7317 43839 7403 43895
rect 7459 43839 7545 43895
rect 7601 43839 7687 43895
rect 7743 43839 7829 43895
rect 7885 43839 7971 43895
rect 8027 43839 8113 43895
rect 8169 43839 8255 43895
rect 8311 43839 8397 43895
rect 8453 43839 8539 43895
rect 8595 43839 8681 43895
rect 8737 43839 8823 43895
rect 8879 43839 8965 43895
rect 9021 43839 9107 43895
rect 9163 43839 9249 43895
rect 9305 43839 9391 43895
rect 9447 43839 9533 43895
rect 9589 43839 9675 43895
rect 9731 43839 9817 43895
rect 9873 43839 9959 43895
rect 10015 43839 10101 43895
rect 10157 43839 10243 43895
rect 10299 43839 10385 43895
rect 10441 43839 10527 43895
rect 10583 43839 10669 43895
rect 10725 43839 10811 43895
rect 10867 43839 10953 43895
rect 11009 43839 11095 43895
rect 11151 43839 11237 43895
rect 11293 43839 11379 43895
rect 11435 43839 11521 43895
rect 11577 43839 11663 43895
rect 11719 43839 11805 43895
rect 11861 43839 11947 43895
rect 12003 43839 12089 43895
rect 12145 43839 12231 43895
rect 12287 43839 12373 43895
rect 12429 43839 12515 43895
rect 12571 43839 12657 43895
rect 12713 43839 12799 43895
rect 12855 43839 12941 43895
rect 12997 43839 13083 43895
rect 13139 43839 13225 43895
rect 13281 43839 13367 43895
rect 13423 43839 13509 43895
rect 13565 43839 13651 43895
rect 13707 43839 13793 43895
rect 13849 43839 13935 43895
rect 13991 43839 14077 43895
rect 14133 43839 14219 43895
rect 14275 43839 14361 43895
rect 14417 43839 14503 43895
rect 14559 43839 14645 43895
rect 14701 43839 14787 43895
rect 14843 43839 14853 43895
rect 151 43753 14853 43839
rect 151 43697 161 43753
rect 217 43697 303 43753
rect 359 43697 445 43753
rect 501 43697 587 43753
rect 643 43697 729 43753
rect 785 43697 871 43753
rect 927 43697 1013 43753
rect 1069 43697 1155 43753
rect 1211 43697 1297 43753
rect 1353 43697 1439 43753
rect 1495 43697 1581 43753
rect 1637 43697 1723 43753
rect 1779 43697 1865 43753
rect 1921 43697 2007 43753
rect 2063 43697 2149 43753
rect 2205 43697 2291 43753
rect 2347 43697 2433 43753
rect 2489 43697 2575 43753
rect 2631 43697 2717 43753
rect 2773 43697 2859 43753
rect 2915 43697 3001 43753
rect 3057 43697 3143 43753
rect 3199 43697 3285 43753
rect 3341 43697 3427 43753
rect 3483 43697 3569 43753
rect 3625 43697 3711 43753
rect 3767 43697 3853 43753
rect 3909 43697 3995 43753
rect 4051 43697 4137 43753
rect 4193 43697 4279 43753
rect 4335 43697 4421 43753
rect 4477 43697 4563 43753
rect 4619 43697 4705 43753
rect 4761 43697 4847 43753
rect 4903 43697 4989 43753
rect 5045 43697 5131 43753
rect 5187 43697 5273 43753
rect 5329 43697 5415 43753
rect 5471 43697 5557 43753
rect 5613 43697 5699 43753
rect 5755 43697 5841 43753
rect 5897 43697 5983 43753
rect 6039 43697 6125 43753
rect 6181 43697 6267 43753
rect 6323 43697 6409 43753
rect 6465 43697 6551 43753
rect 6607 43697 6693 43753
rect 6749 43697 6835 43753
rect 6891 43697 6977 43753
rect 7033 43697 7119 43753
rect 7175 43697 7261 43753
rect 7317 43697 7403 43753
rect 7459 43697 7545 43753
rect 7601 43697 7687 43753
rect 7743 43697 7829 43753
rect 7885 43697 7971 43753
rect 8027 43697 8113 43753
rect 8169 43697 8255 43753
rect 8311 43697 8397 43753
rect 8453 43697 8539 43753
rect 8595 43697 8681 43753
rect 8737 43697 8823 43753
rect 8879 43697 8965 43753
rect 9021 43697 9107 43753
rect 9163 43697 9249 43753
rect 9305 43697 9391 43753
rect 9447 43697 9533 43753
rect 9589 43697 9675 43753
rect 9731 43697 9817 43753
rect 9873 43697 9959 43753
rect 10015 43697 10101 43753
rect 10157 43697 10243 43753
rect 10299 43697 10385 43753
rect 10441 43697 10527 43753
rect 10583 43697 10669 43753
rect 10725 43697 10811 43753
rect 10867 43697 10953 43753
rect 11009 43697 11095 43753
rect 11151 43697 11237 43753
rect 11293 43697 11379 43753
rect 11435 43697 11521 43753
rect 11577 43697 11663 43753
rect 11719 43697 11805 43753
rect 11861 43697 11947 43753
rect 12003 43697 12089 43753
rect 12145 43697 12231 43753
rect 12287 43697 12373 43753
rect 12429 43697 12515 43753
rect 12571 43697 12657 43753
rect 12713 43697 12799 43753
rect 12855 43697 12941 43753
rect 12997 43697 13083 43753
rect 13139 43697 13225 43753
rect 13281 43697 13367 43753
rect 13423 43697 13509 43753
rect 13565 43697 13651 43753
rect 13707 43697 13793 43753
rect 13849 43697 13935 43753
rect 13991 43697 14077 43753
rect 14133 43697 14219 43753
rect 14275 43697 14361 43753
rect 14417 43697 14503 43753
rect 14559 43697 14645 43753
rect 14701 43697 14787 43753
rect 14843 43697 14853 43753
rect 151 43611 14853 43697
rect 151 43555 161 43611
rect 217 43555 303 43611
rect 359 43555 445 43611
rect 501 43555 587 43611
rect 643 43555 729 43611
rect 785 43555 871 43611
rect 927 43555 1013 43611
rect 1069 43555 1155 43611
rect 1211 43555 1297 43611
rect 1353 43555 1439 43611
rect 1495 43555 1581 43611
rect 1637 43555 1723 43611
rect 1779 43555 1865 43611
rect 1921 43555 2007 43611
rect 2063 43555 2149 43611
rect 2205 43555 2291 43611
rect 2347 43555 2433 43611
rect 2489 43555 2575 43611
rect 2631 43555 2717 43611
rect 2773 43555 2859 43611
rect 2915 43555 3001 43611
rect 3057 43555 3143 43611
rect 3199 43555 3285 43611
rect 3341 43555 3427 43611
rect 3483 43555 3569 43611
rect 3625 43555 3711 43611
rect 3767 43555 3853 43611
rect 3909 43555 3995 43611
rect 4051 43555 4137 43611
rect 4193 43555 4279 43611
rect 4335 43555 4421 43611
rect 4477 43555 4563 43611
rect 4619 43555 4705 43611
rect 4761 43555 4847 43611
rect 4903 43555 4989 43611
rect 5045 43555 5131 43611
rect 5187 43555 5273 43611
rect 5329 43555 5415 43611
rect 5471 43555 5557 43611
rect 5613 43555 5699 43611
rect 5755 43555 5841 43611
rect 5897 43555 5983 43611
rect 6039 43555 6125 43611
rect 6181 43555 6267 43611
rect 6323 43555 6409 43611
rect 6465 43555 6551 43611
rect 6607 43555 6693 43611
rect 6749 43555 6835 43611
rect 6891 43555 6977 43611
rect 7033 43555 7119 43611
rect 7175 43555 7261 43611
rect 7317 43555 7403 43611
rect 7459 43555 7545 43611
rect 7601 43555 7687 43611
rect 7743 43555 7829 43611
rect 7885 43555 7971 43611
rect 8027 43555 8113 43611
rect 8169 43555 8255 43611
rect 8311 43555 8397 43611
rect 8453 43555 8539 43611
rect 8595 43555 8681 43611
rect 8737 43555 8823 43611
rect 8879 43555 8965 43611
rect 9021 43555 9107 43611
rect 9163 43555 9249 43611
rect 9305 43555 9391 43611
rect 9447 43555 9533 43611
rect 9589 43555 9675 43611
rect 9731 43555 9817 43611
rect 9873 43555 9959 43611
rect 10015 43555 10101 43611
rect 10157 43555 10243 43611
rect 10299 43555 10385 43611
rect 10441 43555 10527 43611
rect 10583 43555 10669 43611
rect 10725 43555 10811 43611
rect 10867 43555 10953 43611
rect 11009 43555 11095 43611
rect 11151 43555 11237 43611
rect 11293 43555 11379 43611
rect 11435 43555 11521 43611
rect 11577 43555 11663 43611
rect 11719 43555 11805 43611
rect 11861 43555 11947 43611
rect 12003 43555 12089 43611
rect 12145 43555 12231 43611
rect 12287 43555 12373 43611
rect 12429 43555 12515 43611
rect 12571 43555 12657 43611
rect 12713 43555 12799 43611
rect 12855 43555 12941 43611
rect 12997 43555 13083 43611
rect 13139 43555 13225 43611
rect 13281 43555 13367 43611
rect 13423 43555 13509 43611
rect 13565 43555 13651 43611
rect 13707 43555 13793 43611
rect 13849 43555 13935 43611
rect 13991 43555 14077 43611
rect 14133 43555 14219 43611
rect 14275 43555 14361 43611
rect 14417 43555 14503 43611
rect 14559 43555 14645 43611
rect 14701 43555 14787 43611
rect 14843 43555 14853 43611
rect 151 43469 14853 43555
rect 151 43413 161 43469
rect 217 43413 303 43469
rect 359 43413 445 43469
rect 501 43413 587 43469
rect 643 43413 729 43469
rect 785 43413 871 43469
rect 927 43413 1013 43469
rect 1069 43413 1155 43469
rect 1211 43413 1297 43469
rect 1353 43413 1439 43469
rect 1495 43413 1581 43469
rect 1637 43413 1723 43469
rect 1779 43413 1865 43469
rect 1921 43413 2007 43469
rect 2063 43413 2149 43469
rect 2205 43413 2291 43469
rect 2347 43413 2433 43469
rect 2489 43413 2575 43469
rect 2631 43413 2717 43469
rect 2773 43413 2859 43469
rect 2915 43413 3001 43469
rect 3057 43413 3143 43469
rect 3199 43413 3285 43469
rect 3341 43413 3427 43469
rect 3483 43413 3569 43469
rect 3625 43413 3711 43469
rect 3767 43413 3853 43469
rect 3909 43413 3995 43469
rect 4051 43413 4137 43469
rect 4193 43413 4279 43469
rect 4335 43413 4421 43469
rect 4477 43413 4563 43469
rect 4619 43413 4705 43469
rect 4761 43413 4847 43469
rect 4903 43413 4989 43469
rect 5045 43413 5131 43469
rect 5187 43413 5273 43469
rect 5329 43413 5415 43469
rect 5471 43413 5557 43469
rect 5613 43413 5699 43469
rect 5755 43413 5841 43469
rect 5897 43413 5983 43469
rect 6039 43413 6125 43469
rect 6181 43413 6267 43469
rect 6323 43413 6409 43469
rect 6465 43413 6551 43469
rect 6607 43413 6693 43469
rect 6749 43413 6835 43469
rect 6891 43413 6977 43469
rect 7033 43413 7119 43469
rect 7175 43413 7261 43469
rect 7317 43413 7403 43469
rect 7459 43413 7545 43469
rect 7601 43413 7687 43469
rect 7743 43413 7829 43469
rect 7885 43413 7971 43469
rect 8027 43413 8113 43469
rect 8169 43413 8255 43469
rect 8311 43413 8397 43469
rect 8453 43413 8539 43469
rect 8595 43413 8681 43469
rect 8737 43413 8823 43469
rect 8879 43413 8965 43469
rect 9021 43413 9107 43469
rect 9163 43413 9249 43469
rect 9305 43413 9391 43469
rect 9447 43413 9533 43469
rect 9589 43413 9675 43469
rect 9731 43413 9817 43469
rect 9873 43413 9959 43469
rect 10015 43413 10101 43469
rect 10157 43413 10243 43469
rect 10299 43413 10385 43469
rect 10441 43413 10527 43469
rect 10583 43413 10669 43469
rect 10725 43413 10811 43469
rect 10867 43413 10953 43469
rect 11009 43413 11095 43469
rect 11151 43413 11237 43469
rect 11293 43413 11379 43469
rect 11435 43413 11521 43469
rect 11577 43413 11663 43469
rect 11719 43413 11805 43469
rect 11861 43413 11947 43469
rect 12003 43413 12089 43469
rect 12145 43413 12231 43469
rect 12287 43413 12373 43469
rect 12429 43413 12515 43469
rect 12571 43413 12657 43469
rect 12713 43413 12799 43469
rect 12855 43413 12941 43469
rect 12997 43413 13083 43469
rect 13139 43413 13225 43469
rect 13281 43413 13367 43469
rect 13423 43413 13509 43469
rect 13565 43413 13651 43469
rect 13707 43413 13793 43469
rect 13849 43413 13935 43469
rect 13991 43413 14077 43469
rect 14133 43413 14219 43469
rect 14275 43413 14361 43469
rect 14417 43413 14503 43469
rect 14559 43413 14645 43469
rect 14701 43413 14787 43469
rect 14843 43413 14853 43469
rect 151 43327 14853 43413
rect 151 43271 161 43327
rect 217 43271 303 43327
rect 359 43271 445 43327
rect 501 43271 587 43327
rect 643 43271 729 43327
rect 785 43271 871 43327
rect 927 43271 1013 43327
rect 1069 43271 1155 43327
rect 1211 43271 1297 43327
rect 1353 43271 1439 43327
rect 1495 43271 1581 43327
rect 1637 43271 1723 43327
rect 1779 43271 1865 43327
rect 1921 43271 2007 43327
rect 2063 43271 2149 43327
rect 2205 43271 2291 43327
rect 2347 43271 2433 43327
rect 2489 43271 2575 43327
rect 2631 43271 2717 43327
rect 2773 43271 2859 43327
rect 2915 43271 3001 43327
rect 3057 43271 3143 43327
rect 3199 43271 3285 43327
rect 3341 43271 3427 43327
rect 3483 43271 3569 43327
rect 3625 43271 3711 43327
rect 3767 43271 3853 43327
rect 3909 43271 3995 43327
rect 4051 43271 4137 43327
rect 4193 43271 4279 43327
rect 4335 43271 4421 43327
rect 4477 43271 4563 43327
rect 4619 43271 4705 43327
rect 4761 43271 4847 43327
rect 4903 43271 4989 43327
rect 5045 43271 5131 43327
rect 5187 43271 5273 43327
rect 5329 43271 5415 43327
rect 5471 43271 5557 43327
rect 5613 43271 5699 43327
rect 5755 43271 5841 43327
rect 5897 43271 5983 43327
rect 6039 43271 6125 43327
rect 6181 43271 6267 43327
rect 6323 43271 6409 43327
rect 6465 43271 6551 43327
rect 6607 43271 6693 43327
rect 6749 43271 6835 43327
rect 6891 43271 6977 43327
rect 7033 43271 7119 43327
rect 7175 43271 7261 43327
rect 7317 43271 7403 43327
rect 7459 43271 7545 43327
rect 7601 43271 7687 43327
rect 7743 43271 7829 43327
rect 7885 43271 7971 43327
rect 8027 43271 8113 43327
rect 8169 43271 8255 43327
rect 8311 43271 8397 43327
rect 8453 43271 8539 43327
rect 8595 43271 8681 43327
rect 8737 43271 8823 43327
rect 8879 43271 8965 43327
rect 9021 43271 9107 43327
rect 9163 43271 9249 43327
rect 9305 43271 9391 43327
rect 9447 43271 9533 43327
rect 9589 43271 9675 43327
rect 9731 43271 9817 43327
rect 9873 43271 9959 43327
rect 10015 43271 10101 43327
rect 10157 43271 10243 43327
rect 10299 43271 10385 43327
rect 10441 43271 10527 43327
rect 10583 43271 10669 43327
rect 10725 43271 10811 43327
rect 10867 43271 10953 43327
rect 11009 43271 11095 43327
rect 11151 43271 11237 43327
rect 11293 43271 11379 43327
rect 11435 43271 11521 43327
rect 11577 43271 11663 43327
rect 11719 43271 11805 43327
rect 11861 43271 11947 43327
rect 12003 43271 12089 43327
rect 12145 43271 12231 43327
rect 12287 43271 12373 43327
rect 12429 43271 12515 43327
rect 12571 43271 12657 43327
rect 12713 43271 12799 43327
rect 12855 43271 12941 43327
rect 12997 43271 13083 43327
rect 13139 43271 13225 43327
rect 13281 43271 13367 43327
rect 13423 43271 13509 43327
rect 13565 43271 13651 43327
rect 13707 43271 13793 43327
rect 13849 43271 13935 43327
rect 13991 43271 14077 43327
rect 14133 43271 14219 43327
rect 14275 43271 14361 43327
rect 14417 43271 14503 43327
rect 14559 43271 14645 43327
rect 14701 43271 14787 43327
rect 14843 43271 14853 43327
rect 151 43185 14853 43271
rect 151 43129 161 43185
rect 217 43129 303 43185
rect 359 43129 445 43185
rect 501 43129 587 43185
rect 643 43129 729 43185
rect 785 43129 871 43185
rect 927 43129 1013 43185
rect 1069 43129 1155 43185
rect 1211 43129 1297 43185
rect 1353 43129 1439 43185
rect 1495 43129 1581 43185
rect 1637 43129 1723 43185
rect 1779 43129 1865 43185
rect 1921 43129 2007 43185
rect 2063 43129 2149 43185
rect 2205 43129 2291 43185
rect 2347 43129 2433 43185
rect 2489 43129 2575 43185
rect 2631 43129 2717 43185
rect 2773 43129 2859 43185
rect 2915 43129 3001 43185
rect 3057 43129 3143 43185
rect 3199 43129 3285 43185
rect 3341 43129 3427 43185
rect 3483 43129 3569 43185
rect 3625 43129 3711 43185
rect 3767 43129 3853 43185
rect 3909 43129 3995 43185
rect 4051 43129 4137 43185
rect 4193 43129 4279 43185
rect 4335 43129 4421 43185
rect 4477 43129 4563 43185
rect 4619 43129 4705 43185
rect 4761 43129 4847 43185
rect 4903 43129 4989 43185
rect 5045 43129 5131 43185
rect 5187 43129 5273 43185
rect 5329 43129 5415 43185
rect 5471 43129 5557 43185
rect 5613 43129 5699 43185
rect 5755 43129 5841 43185
rect 5897 43129 5983 43185
rect 6039 43129 6125 43185
rect 6181 43129 6267 43185
rect 6323 43129 6409 43185
rect 6465 43129 6551 43185
rect 6607 43129 6693 43185
rect 6749 43129 6835 43185
rect 6891 43129 6977 43185
rect 7033 43129 7119 43185
rect 7175 43129 7261 43185
rect 7317 43129 7403 43185
rect 7459 43129 7545 43185
rect 7601 43129 7687 43185
rect 7743 43129 7829 43185
rect 7885 43129 7971 43185
rect 8027 43129 8113 43185
rect 8169 43129 8255 43185
rect 8311 43129 8397 43185
rect 8453 43129 8539 43185
rect 8595 43129 8681 43185
rect 8737 43129 8823 43185
rect 8879 43129 8965 43185
rect 9021 43129 9107 43185
rect 9163 43129 9249 43185
rect 9305 43129 9391 43185
rect 9447 43129 9533 43185
rect 9589 43129 9675 43185
rect 9731 43129 9817 43185
rect 9873 43129 9959 43185
rect 10015 43129 10101 43185
rect 10157 43129 10243 43185
rect 10299 43129 10385 43185
rect 10441 43129 10527 43185
rect 10583 43129 10669 43185
rect 10725 43129 10811 43185
rect 10867 43129 10953 43185
rect 11009 43129 11095 43185
rect 11151 43129 11237 43185
rect 11293 43129 11379 43185
rect 11435 43129 11521 43185
rect 11577 43129 11663 43185
rect 11719 43129 11805 43185
rect 11861 43129 11947 43185
rect 12003 43129 12089 43185
rect 12145 43129 12231 43185
rect 12287 43129 12373 43185
rect 12429 43129 12515 43185
rect 12571 43129 12657 43185
rect 12713 43129 12799 43185
rect 12855 43129 12941 43185
rect 12997 43129 13083 43185
rect 13139 43129 13225 43185
rect 13281 43129 13367 43185
rect 13423 43129 13509 43185
rect 13565 43129 13651 43185
rect 13707 43129 13793 43185
rect 13849 43129 13935 43185
rect 13991 43129 14077 43185
rect 14133 43129 14219 43185
rect 14275 43129 14361 43185
rect 14417 43129 14503 43185
rect 14559 43129 14645 43185
rect 14701 43129 14787 43185
rect 14843 43129 14853 43185
rect 151 43043 14853 43129
rect 151 42987 161 43043
rect 217 42987 303 43043
rect 359 42987 445 43043
rect 501 42987 587 43043
rect 643 42987 729 43043
rect 785 42987 871 43043
rect 927 42987 1013 43043
rect 1069 42987 1155 43043
rect 1211 42987 1297 43043
rect 1353 42987 1439 43043
rect 1495 42987 1581 43043
rect 1637 42987 1723 43043
rect 1779 42987 1865 43043
rect 1921 42987 2007 43043
rect 2063 42987 2149 43043
rect 2205 42987 2291 43043
rect 2347 42987 2433 43043
rect 2489 42987 2575 43043
rect 2631 42987 2717 43043
rect 2773 42987 2859 43043
rect 2915 42987 3001 43043
rect 3057 42987 3143 43043
rect 3199 42987 3285 43043
rect 3341 42987 3427 43043
rect 3483 42987 3569 43043
rect 3625 42987 3711 43043
rect 3767 42987 3853 43043
rect 3909 42987 3995 43043
rect 4051 42987 4137 43043
rect 4193 42987 4279 43043
rect 4335 42987 4421 43043
rect 4477 42987 4563 43043
rect 4619 42987 4705 43043
rect 4761 42987 4847 43043
rect 4903 42987 4989 43043
rect 5045 42987 5131 43043
rect 5187 42987 5273 43043
rect 5329 42987 5415 43043
rect 5471 42987 5557 43043
rect 5613 42987 5699 43043
rect 5755 42987 5841 43043
rect 5897 42987 5983 43043
rect 6039 42987 6125 43043
rect 6181 42987 6267 43043
rect 6323 42987 6409 43043
rect 6465 42987 6551 43043
rect 6607 42987 6693 43043
rect 6749 42987 6835 43043
rect 6891 42987 6977 43043
rect 7033 42987 7119 43043
rect 7175 42987 7261 43043
rect 7317 42987 7403 43043
rect 7459 42987 7545 43043
rect 7601 42987 7687 43043
rect 7743 42987 7829 43043
rect 7885 42987 7971 43043
rect 8027 42987 8113 43043
rect 8169 42987 8255 43043
rect 8311 42987 8397 43043
rect 8453 42987 8539 43043
rect 8595 42987 8681 43043
rect 8737 42987 8823 43043
rect 8879 42987 8965 43043
rect 9021 42987 9107 43043
rect 9163 42987 9249 43043
rect 9305 42987 9391 43043
rect 9447 42987 9533 43043
rect 9589 42987 9675 43043
rect 9731 42987 9817 43043
rect 9873 42987 9959 43043
rect 10015 42987 10101 43043
rect 10157 42987 10243 43043
rect 10299 42987 10385 43043
rect 10441 42987 10527 43043
rect 10583 42987 10669 43043
rect 10725 42987 10811 43043
rect 10867 42987 10953 43043
rect 11009 42987 11095 43043
rect 11151 42987 11237 43043
rect 11293 42987 11379 43043
rect 11435 42987 11521 43043
rect 11577 42987 11663 43043
rect 11719 42987 11805 43043
rect 11861 42987 11947 43043
rect 12003 42987 12089 43043
rect 12145 42987 12231 43043
rect 12287 42987 12373 43043
rect 12429 42987 12515 43043
rect 12571 42987 12657 43043
rect 12713 42987 12799 43043
rect 12855 42987 12941 43043
rect 12997 42987 13083 43043
rect 13139 42987 13225 43043
rect 13281 42987 13367 43043
rect 13423 42987 13509 43043
rect 13565 42987 13651 43043
rect 13707 42987 13793 43043
rect 13849 42987 13935 43043
rect 13991 42987 14077 43043
rect 14133 42987 14219 43043
rect 14275 42987 14361 43043
rect 14417 42987 14503 43043
rect 14559 42987 14645 43043
rect 14701 42987 14787 43043
rect 14843 42987 14853 43043
rect 151 42901 14853 42987
rect 151 42845 161 42901
rect 217 42845 303 42901
rect 359 42845 445 42901
rect 501 42845 587 42901
rect 643 42845 729 42901
rect 785 42845 871 42901
rect 927 42845 1013 42901
rect 1069 42845 1155 42901
rect 1211 42845 1297 42901
rect 1353 42845 1439 42901
rect 1495 42845 1581 42901
rect 1637 42845 1723 42901
rect 1779 42845 1865 42901
rect 1921 42845 2007 42901
rect 2063 42845 2149 42901
rect 2205 42845 2291 42901
rect 2347 42845 2433 42901
rect 2489 42845 2575 42901
rect 2631 42845 2717 42901
rect 2773 42845 2859 42901
rect 2915 42845 3001 42901
rect 3057 42845 3143 42901
rect 3199 42845 3285 42901
rect 3341 42845 3427 42901
rect 3483 42845 3569 42901
rect 3625 42845 3711 42901
rect 3767 42845 3853 42901
rect 3909 42845 3995 42901
rect 4051 42845 4137 42901
rect 4193 42845 4279 42901
rect 4335 42845 4421 42901
rect 4477 42845 4563 42901
rect 4619 42845 4705 42901
rect 4761 42845 4847 42901
rect 4903 42845 4989 42901
rect 5045 42845 5131 42901
rect 5187 42845 5273 42901
rect 5329 42845 5415 42901
rect 5471 42845 5557 42901
rect 5613 42845 5699 42901
rect 5755 42845 5841 42901
rect 5897 42845 5983 42901
rect 6039 42845 6125 42901
rect 6181 42845 6267 42901
rect 6323 42845 6409 42901
rect 6465 42845 6551 42901
rect 6607 42845 6693 42901
rect 6749 42845 6835 42901
rect 6891 42845 6977 42901
rect 7033 42845 7119 42901
rect 7175 42845 7261 42901
rect 7317 42845 7403 42901
rect 7459 42845 7545 42901
rect 7601 42845 7687 42901
rect 7743 42845 7829 42901
rect 7885 42845 7971 42901
rect 8027 42845 8113 42901
rect 8169 42845 8255 42901
rect 8311 42845 8397 42901
rect 8453 42845 8539 42901
rect 8595 42845 8681 42901
rect 8737 42845 8823 42901
rect 8879 42845 8965 42901
rect 9021 42845 9107 42901
rect 9163 42845 9249 42901
rect 9305 42845 9391 42901
rect 9447 42845 9533 42901
rect 9589 42845 9675 42901
rect 9731 42845 9817 42901
rect 9873 42845 9959 42901
rect 10015 42845 10101 42901
rect 10157 42845 10243 42901
rect 10299 42845 10385 42901
rect 10441 42845 10527 42901
rect 10583 42845 10669 42901
rect 10725 42845 10811 42901
rect 10867 42845 10953 42901
rect 11009 42845 11095 42901
rect 11151 42845 11237 42901
rect 11293 42845 11379 42901
rect 11435 42845 11521 42901
rect 11577 42845 11663 42901
rect 11719 42845 11805 42901
rect 11861 42845 11947 42901
rect 12003 42845 12089 42901
rect 12145 42845 12231 42901
rect 12287 42845 12373 42901
rect 12429 42845 12515 42901
rect 12571 42845 12657 42901
rect 12713 42845 12799 42901
rect 12855 42845 12941 42901
rect 12997 42845 13083 42901
rect 13139 42845 13225 42901
rect 13281 42845 13367 42901
rect 13423 42845 13509 42901
rect 13565 42845 13651 42901
rect 13707 42845 13793 42901
rect 13849 42845 13935 42901
rect 13991 42845 14077 42901
rect 14133 42845 14219 42901
rect 14275 42845 14361 42901
rect 14417 42845 14503 42901
rect 14559 42845 14645 42901
rect 14701 42845 14787 42901
rect 14843 42845 14853 42901
rect 151 42835 14853 42845
rect 151 42563 14853 42573
rect 151 42507 161 42563
rect 217 42507 303 42563
rect 359 42507 445 42563
rect 501 42507 587 42563
rect 643 42507 729 42563
rect 785 42507 871 42563
rect 927 42507 1013 42563
rect 1069 42507 1155 42563
rect 1211 42507 1297 42563
rect 1353 42507 1439 42563
rect 1495 42507 1581 42563
rect 1637 42507 1723 42563
rect 1779 42507 1865 42563
rect 1921 42507 2007 42563
rect 2063 42507 2149 42563
rect 2205 42507 2291 42563
rect 2347 42507 2433 42563
rect 2489 42507 2575 42563
rect 2631 42507 2717 42563
rect 2773 42507 2859 42563
rect 2915 42507 3001 42563
rect 3057 42507 3143 42563
rect 3199 42507 3285 42563
rect 3341 42507 3427 42563
rect 3483 42507 3569 42563
rect 3625 42507 3711 42563
rect 3767 42507 3853 42563
rect 3909 42507 3995 42563
rect 4051 42507 4137 42563
rect 4193 42507 4279 42563
rect 4335 42507 4421 42563
rect 4477 42507 4563 42563
rect 4619 42507 4705 42563
rect 4761 42507 4847 42563
rect 4903 42507 4989 42563
rect 5045 42507 5131 42563
rect 5187 42507 5273 42563
rect 5329 42507 5415 42563
rect 5471 42507 5557 42563
rect 5613 42507 5699 42563
rect 5755 42507 5841 42563
rect 5897 42507 5983 42563
rect 6039 42507 6125 42563
rect 6181 42507 6267 42563
rect 6323 42507 6409 42563
rect 6465 42507 6551 42563
rect 6607 42507 6693 42563
rect 6749 42507 6835 42563
rect 6891 42507 6977 42563
rect 7033 42507 7119 42563
rect 7175 42507 7261 42563
rect 7317 42507 7403 42563
rect 7459 42507 7545 42563
rect 7601 42507 7687 42563
rect 7743 42507 7829 42563
rect 7885 42507 7971 42563
rect 8027 42507 8113 42563
rect 8169 42507 8255 42563
rect 8311 42507 8397 42563
rect 8453 42507 8539 42563
rect 8595 42507 8681 42563
rect 8737 42507 8823 42563
rect 8879 42507 8965 42563
rect 9021 42507 9107 42563
rect 9163 42507 9249 42563
rect 9305 42507 9391 42563
rect 9447 42507 9533 42563
rect 9589 42507 9675 42563
rect 9731 42507 9817 42563
rect 9873 42507 9959 42563
rect 10015 42507 10101 42563
rect 10157 42507 10243 42563
rect 10299 42507 10385 42563
rect 10441 42507 10527 42563
rect 10583 42507 10669 42563
rect 10725 42507 10811 42563
rect 10867 42507 10953 42563
rect 11009 42507 11095 42563
rect 11151 42507 11237 42563
rect 11293 42507 11379 42563
rect 11435 42507 11521 42563
rect 11577 42507 11663 42563
rect 11719 42507 11805 42563
rect 11861 42507 11947 42563
rect 12003 42507 12089 42563
rect 12145 42507 12231 42563
rect 12287 42507 12373 42563
rect 12429 42507 12515 42563
rect 12571 42507 12657 42563
rect 12713 42507 12799 42563
rect 12855 42507 12941 42563
rect 12997 42507 13083 42563
rect 13139 42507 13225 42563
rect 13281 42507 13367 42563
rect 13423 42507 13509 42563
rect 13565 42507 13651 42563
rect 13707 42507 13793 42563
rect 13849 42507 13935 42563
rect 13991 42507 14077 42563
rect 14133 42507 14219 42563
rect 14275 42507 14361 42563
rect 14417 42507 14503 42563
rect 14559 42507 14645 42563
rect 14701 42507 14787 42563
rect 14843 42507 14853 42563
rect 151 42421 14853 42507
rect 151 42365 161 42421
rect 217 42365 303 42421
rect 359 42365 445 42421
rect 501 42365 587 42421
rect 643 42365 729 42421
rect 785 42365 871 42421
rect 927 42365 1013 42421
rect 1069 42365 1155 42421
rect 1211 42365 1297 42421
rect 1353 42365 1439 42421
rect 1495 42365 1581 42421
rect 1637 42365 1723 42421
rect 1779 42365 1865 42421
rect 1921 42365 2007 42421
rect 2063 42365 2149 42421
rect 2205 42365 2291 42421
rect 2347 42365 2433 42421
rect 2489 42365 2575 42421
rect 2631 42365 2717 42421
rect 2773 42365 2859 42421
rect 2915 42365 3001 42421
rect 3057 42365 3143 42421
rect 3199 42365 3285 42421
rect 3341 42365 3427 42421
rect 3483 42365 3569 42421
rect 3625 42365 3711 42421
rect 3767 42365 3853 42421
rect 3909 42365 3995 42421
rect 4051 42365 4137 42421
rect 4193 42365 4279 42421
rect 4335 42365 4421 42421
rect 4477 42365 4563 42421
rect 4619 42365 4705 42421
rect 4761 42365 4847 42421
rect 4903 42365 4989 42421
rect 5045 42365 5131 42421
rect 5187 42365 5273 42421
rect 5329 42365 5415 42421
rect 5471 42365 5557 42421
rect 5613 42365 5699 42421
rect 5755 42365 5841 42421
rect 5897 42365 5983 42421
rect 6039 42365 6125 42421
rect 6181 42365 6267 42421
rect 6323 42365 6409 42421
rect 6465 42365 6551 42421
rect 6607 42365 6693 42421
rect 6749 42365 6835 42421
rect 6891 42365 6977 42421
rect 7033 42365 7119 42421
rect 7175 42365 7261 42421
rect 7317 42365 7403 42421
rect 7459 42365 7545 42421
rect 7601 42365 7687 42421
rect 7743 42365 7829 42421
rect 7885 42365 7971 42421
rect 8027 42365 8113 42421
rect 8169 42365 8255 42421
rect 8311 42365 8397 42421
rect 8453 42365 8539 42421
rect 8595 42365 8681 42421
rect 8737 42365 8823 42421
rect 8879 42365 8965 42421
rect 9021 42365 9107 42421
rect 9163 42365 9249 42421
rect 9305 42365 9391 42421
rect 9447 42365 9533 42421
rect 9589 42365 9675 42421
rect 9731 42365 9817 42421
rect 9873 42365 9959 42421
rect 10015 42365 10101 42421
rect 10157 42365 10243 42421
rect 10299 42365 10385 42421
rect 10441 42365 10527 42421
rect 10583 42365 10669 42421
rect 10725 42365 10811 42421
rect 10867 42365 10953 42421
rect 11009 42365 11095 42421
rect 11151 42365 11237 42421
rect 11293 42365 11379 42421
rect 11435 42365 11521 42421
rect 11577 42365 11663 42421
rect 11719 42365 11805 42421
rect 11861 42365 11947 42421
rect 12003 42365 12089 42421
rect 12145 42365 12231 42421
rect 12287 42365 12373 42421
rect 12429 42365 12515 42421
rect 12571 42365 12657 42421
rect 12713 42365 12799 42421
rect 12855 42365 12941 42421
rect 12997 42365 13083 42421
rect 13139 42365 13225 42421
rect 13281 42365 13367 42421
rect 13423 42365 13509 42421
rect 13565 42365 13651 42421
rect 13707 42365 13793 42421
rect 13849 42365 13935 42421
rect 13991 42365 14077 42421
rect 14133 42365 14219 42421
rect 14275 42365 14361 42421
rect 14417 42365 14503 42421
rect 14559 42365 14645 42421
rect 14701 42365 14787 42421
rect 14843 42365 14853 42421
rect 151 42279 14853 42365
rect 151 42223 161 42279
rect 217 42223 303 42279
rect 359 42223 445 42279
rect 501 42223 587 42279
rect 643 42223 729 42279
rect 785 42223 871 42279
rect 927 42223 1013 42279
rect 1069 42223 1155 42279
rect 1211 42223 1297 42279
rect 1353 42223 1439 42279
rect 1495 42223 1581 42279
rect 1637 42223 1723 42279
rect 1779 42223 1865 42279
rect 1921 42223 2007 42279
rect 2063 42223 2149 42279
rect 2205 42223 2291 42279
rect 2347 42223 2433 42279
rect 2489 42223 2575 42279
rect 2631 42223 2717 42279
rect 2773 42223 2859 42279
rect 2915 42223 3001 42279
rect 3057 42223 3143 42279
rect 3199 42223 3285 42279
rect 3341 42223 3427 42279
rect 3483 42223 3569 42279
rect 3625 42223 3711 42279
rect 3767 42223 3853 42279
rect 3909 42223 3995 42279
rect 4051 42223 4137 42279
rect 4193 42223 4279 42279
rect 4335 42223 4421 42279
rect 4477 42223 4563 42279
rect 4619 42223 4705 42279
rect 4761 42223 4847 42279
rect 4903 42223 4989 42279
rect 5045 42223 5131 42279
rect 5187 42223 5273 42279
rect 5329 42223 5415 42279
rect 5471 42223 5557 42279
rect 5613 42223 5699 42279
rect 5755 42223 5841 42279
rect 5897 42223 5983 42279
rect 6039 42223 6125 42279
rect 6181 42223 6267 42279
rect 6323 42223 6409 42279
rect 6465 42223 6551 42279
rect 6607 42223 6693 42279
rect 6749 42223 6835 42279
rect 6891 42223 6977 42279
rect 7033 42223 7119 42279
rect 7175 42223 7261 42279
rect 7317 42223 7403 42279
rect 7459 42223 7545 42279
rect 7601 42223 7687 42279
rect 7743 42223 7829 42279
rect 7885 42223 7971 42279
rect 8027 42223 8113 42279
rect 8169 42223 8255 42279
rect 8311 42223 8397 42279
rect 8453 42223 8539 42279
rect 8595 42223 8681 42279
rect 8737 42223 8823 42279
rect 8879 42223 8965 42279
rect 9021 42223 9107 42279
rect 9163 42223 9249 42279
rect 9305 42223 9391 42279
rect 9447 42223 9533 42279
rect 9589 42223 9675 42279
rect 9731 42223 9817 42279
rect 9873 42223 9959 42279
rect 10015 42223 10101 42279
rect 10157 42223 10243 42279
rect 10299 42223 10385 42279
rect 10441 42223 10527 42279
rect 10583 42223 10669 42279
rect 10725 42223 10811 42279
rect 10867 42223 10953 42279
rect 11009 42223 11095 42279
rect 11151 42223 11237 42279
rect 11293 42223 11379 42279
rect 11435 42223 11521 42279
rect 11577 42223 11663 42279
rect 11719 42223 11805 42279
rect 11861 42223 11947 42279
rect 12003 42223 12089 42279
rect 12145 42223 12231 42279
rect 12287 42223 12373 42279
rect 12429 42223 12515 42279
rect 12571 42223 12657 42279
rect 12713 42223 12799 42279
rect 12855 42223 12941 42279
rect 12997 42223 13083 42279
rect 13139 42223 13225 42279
rect 13281 42223 13367 42279
rect 13423 42223 13509 42279
rect 13565 42223 13651 42279
rect 13707 42223 13793 42279
rect 13849 42223 13935 42279
rect 13991 42223 14077 42279
rect 14133 42223 14219 42279
rect 14275 42223 14361 42279
rect 14417 42223 14503 42279
rect 14559 42223 14645 42279
rect 14701 42223 14787 42279
rect 14843 42223 14853 42279
rect 151 42137 14853 42223
rect 151 42081 161 42137
rect 217 42081 303 42137
rect 359 42081 445 42137
rect 501 42081 587 42137
rect 643 42081 729 42137
rect 785 42081 871 42137
rect 927 42081 1013 42137
rect 1069 42081 1155 42137
rect 1211 42081 1297 42137
rect 1353 42081 1439 42137
rect 1495 42081 1581 42137
rect 1637 42081 1723 42137
rect 1779 42081 1865 42137
rect 1921 42081 2007 42137
rect 2063 42081 2149 42137
rect 2205 42081 2291 42137
rect 2347 42081 2433 42137
rect 2489 42081 2575 42137
rect 2631 42081 2717 42137
rect 2773 42081 2859 42137
rect 2915 42081 3001 42137
rect 3057 42081 3143 42137
rect 3199 42081 3285 42137
rect 3341 42081 3427 42137
rect 3483 42081 3569 42137
rect 3625 42081 3711 42137
rect 3767 42081 3853 42137
rect 3909 42081 3995 42137
rect 4051 42081 4137 42137
rect 4193 42081 4279 42137
rect 4335 42081 4421 42137
rect 4477 42081 4563 42137
rect 4619 42081 4705 42137
rect 4761 42081 4847 42137
rect 4903 42081 4989 42137
rect 5045 42081 5131 42137
rect 5187 42081 5273 42137
rect 5329 42081 5415 42137
rect 5471 42081 5557 42137
rect 5613 42081 5699 42137
rect 5755 42081 5841 42137
rect 5897 42081 5983 42137
rect 6039 42081 6125 42137
rect 6181 42081 6267 42137
rect 6323 42081 6409 42137
rect 6465 42081 6551 42137
rect 6607 42081 6693 42137
rect 6749 42081 6835 42137
rect 6891 42081 6977 42137
rect 7033 42081 7119 42137
rect 7175 42081 7261 42137
rect 7317 42081 7403 42137
rect 7459 42081 7545 42137
rect 7601 42081 7687 42137
rect 7743 42081 7829 42137
rect 7885 42081 7971 42137
rect 8027 42081 8113 42137
rect 8169 42081 8255 42137
rect 8311 42081 8397 42137
rect 8453 42081 8539 42137
rect 8595 42081 8681 42137
rect 8737 42081 8823 42137
rect 8879 42081 8965 42137
rect 9021 42081 9107 42137
rect 9163 42081 9249 42137
rect 9305 42081 9391 42137
rect 9447 42081 9533 42137
rect 9589 42081 9675 42137
rect 9731 42081 9817 42137
rect 9873 42081 9959 42137
rect 10015 42081 10101 42137
rect 10157 42081 10243 42137
rect 10299 42081 10385 42137
rect 10441 42081 10527 42137
rect 10583 42081 10669 42137
rect 10725 42081 10811 42137
rect 10867 42081 10953 42137
rect 11009 42081 11095 42137
rect 11151 42081 11237 42137
rect 11293 42081 11379 42137
rect 11435 42081 11521 42137
rect 11577 42081 11663 42137
rect 11719 42081 11805 42137
rect 11861 42081 11947 42137
rect 12003 42081 12089 42137
rect 12145 42081 12231 42137
rect 12287 42081 12373 42137
rect 12429 42081 12515 42137
rect 12571 42081 12657 42137
rect 12713 42081 12799 42137
rect 12855 42081 12941 42137
rect 12997 42081 13083 42137
rect 13139 42081 13225 42137
rect 13281 42081 13367 42137
rect 13423 42081 13509 42137
rect 13565 42081 13651 42137
rect 13707 42081 13793 42137
rect 13849 42081 13935 42137
rect 13991 42081 14077 42137
rect 14133 42081 14219 42137
rect 14275 42081 14361 42137
rect 14417 42081 14503 42137
rect 14559 42081 14645 42137
rect 14701 42081 14787 42137
rect 14843 42081 14853 42137
rect 151 41995 14853 42081
rect 151 41939 161 41995
rect 217 41939 303 41995
rect 359 41939 445 41995
rect 501 41939 587 41995
rect 643 41939 729 41995
rect 785 41939 871 41995
rect 927 41939 1013 41995
rect 1069 41939 1155 41995
rect 1211 41939 1297 41995
rect 1353 41939 1439 41995
rect 1495 41939 1581 41995
rect 1637 41939 1723 41995
rect 1779 41939 1865 41995
rect 1921 41939 2007 41995
rect 2063 41939 2149 41995
rect 2205 41939 2291 41995
rect 2347 41939 2433 41995
rect 2489 41939 2575 41995
rect 2631 41939 2717 41995
rect 2773 41939 2859 41995
rect 2915 41939 3001 41995
rect 3057 41939 3143 41995
rect 3199 41939 3285 41995
rect 3341 41939 3427 41995
rect 3483 41939 3569 41995
rect 3625 41939 3711 41995
rect 3767 41939 3853 41995
rect 3909 41939 3995 41995
rect 4051 41939 4137 41995
rect 4193 41939 4279 41995
rect 4335 41939 4421 41995
rect 4477 41939 4563 41995
rect 4619 41939 4705 41995
rect 4761 41939 4847 41995
rect 4903 41939 4989 41995
rect 5045 41939 5131 41995
rect 5187 41939 5273 41995
rect 5329 41939 5415 41995
rect 5471 41939 5557 41995
rect 5613 41939 5699 41995
rect 5755 41939 5841 41995
rect 5897 41939 5983 41995
rect 6039 41939 6125 41995
rect 6181 41939 6267 41995
rect 6323 41939 6409 41995
rect 6465 41939 6551 41995
rect 6607 41939 6693 41995
rect 6749 41939 6835 41995
rect 6891 41939 6977 41995
rect 7033 41939 7119 41995
rect 7175 41939 7261 41995
rect 7317 41939 7403 41995
rect 7459 41939 7545 41995
rect 7601 41939 7687 41995
rect 7743 41939 7829 41995
rect 7885 41939 7971 41995
rect 8027 41939 8113 41995
rect 8169 41939 8255 41995
rect 8311 41939 8397 41995
rect 8453 41939 8539 41995
rect 8595 41939 8681 41995
rect 8737 41939 8823 41995
rect 8879 41939 8965 41995
rect 9021 41939 9107 41995
rect 9163 41939 9249 41995
rect 9305 41939 9391 41995
rect 9447 41939 9533 41995
rect 9589 41939 9675 41995
rect 9731 41939 9817 41995
rect 9873 41939 9959 41995
rect 10015 41939 10101 41995
rect 10157 41939 10243 41995
rect 10299 41939 10385 41995
rect 10441 41939 10527 41995
rect 10583 41939 10669 41995
rect 10725 41939 10811 41995
rect 10867 41939 10953 41995
rect 11009 41939 11095 41995
rect 11151 41939 11237 41995
rect 11293 41939 11379 41995
rect 11435 41939 11521 41995
rect 11577 41939 11663 41995
rect 11719 41939 11805 41995
rect 11861 41939 11947 41995
rect 12003 41939 12089 41995
rect 12145 41939 12231 41995
rect 12287 41939 12373 41995
rect 12429 41939 12515 41995
rect 12571 41939 12657 41995
rect 12713 41939 12799 41995
rect 12855 41939 12941 41995
rect 12997 41939 13083 41995
rect 13139 41939 13225 41995
rect 13281 41939 13367 41995
rect 13423 41939 13509 41995
rect 13565 41939 13651 41995
rect 13707 41939 13793 41995
rect 13849 41939 13935 41995
rect 13991 41939 14077 41995
rect 14133 41939 14219 41995
rect 14275 41939 14361 41995
rect 14417 41939 14503 41995
rect 14559 41939 14645 41995
rect 14701 41939 14787 41995
rect 14843 41939 14853 41995
rect 151 41853 14853 41939
rect 151 41797 161 41853
rect 217 41797 303 41853
rect 359 41797 445 41853
rect 501 41797 587 41853
rect 643 41797 729 41853
rect 785 41797 871 41853
rect 927 41797 1013 41853
rect 1069 41797 1155 41853
rect 1211 41797 1297 41853
rect 1353 41797 1439 41853
rect 1495 41797 1581 41853
rect 1637 41797 1723 41853
rect 1779 41797 1865 41853
rect 1921 41797 2007 41853
rect 2063 41797 2149 41853
rect 2205 41797 2291 41853
rect 2347 41797 2433 41853
rect 2489 41797 2575 41853
rect 2631 41797 2717 41853
rect 2773 41797 2859 41853
rect 2915 41797 3001 41853
rect 3057 41797 3143 41853
rect 3199 41797 3285 41853
rect 3341 41797 3427 41853
rect 3483 41797 3569 41853
rect 3625 41797 3711 41853
rect 3767 41797 3853 41853
rect 3909 41797 3995 41853
rect 4051 41797 4137 41853
rect 4193 41797 4279 41853
rect 4335 41797 4421 41853
rect 4477 41797 4563 41853
rect 4619 41797 4705 41853
rect 4761 41797 4847 41853
rect 4903 41797 4989 41853
rect 5045 41797 5131 41853
rect 5187 41797 5273 41853
rect 5329 41797 5415 41853
rect 5471 41797 5557 41853
rect 5613 41797 5699 41853
rect 5755 41797 5841 41853
rect 5897 41797 5983 41853
rect 6039 41797 6125 41853
rect 6181 41797 6267 41853
rect 6323 41797 6409 41853
rect 6465 41797 6551 41853
rect 6607 41797 6693 41853
rect 6749 41797 6835 41853
rect 6891 41797 6977 41853
rect 7033 41797 7119 41853
rect 7175 41797 7261 41853
rect 7317 41797 7403 41853
rect 7459 41797 7545 41853
rect 7601 41797 7687 41853
rect 7743 41797 7829 41853
rect 7885 41797 7971 41853
rect 8027 41797 8113 41853
rect 8169 41797 8255 41853
rect 8311 41797 8397 41853
rect 8453 41797 8539 41853
rect 8595 41797 8681 41853
rect 8737 41797 8823 41853
rect 8879 41797 8965 41853
rect 9021 41797 9107 41853
rect 9163 41797 9249 41853
rect 9305 41797 9391 41853
rect 9447 41797 9533 41853
rect 9589 41797 9675 41853
rect 9731 41797 9817 41853
rect 9873 41797 9959 41853
rect 10015 41797 10101 41853
rect 10157 41797 10243 41853
rect 10299 41797 10385 41853
rect 10441 41797 10527 41853
rect 10583 41797 10669 41853
rect 10725 41797 10811 41853
rect 10867 41797 10953 41853
rect 11009 41797 11095 41853
rect 11151 41797 11237 41853
rect 11293 41797 11379 41853
rect 11435 41797 11521 41853
rect 11577 41797 11663 41853
rect 11719 41797 11805 41853
rect 11861 41797 11947 41853
rect 12003 41797 12089 41853
rect 12145 41797 12231 41853
rect 12287 41797 12373 41853
rect 12429 41797 12515 41853
rect 12571 41797 12657 41853
rect 12713 41797 12799 41853
rect 12855 41797 12941 41853
rect 12997 41797 13083 41853
rect 13139 41797 13225 41853
rect 13281 41797 13367 41853
rect 13423 41797 13509 41853
rect 13565 41797 13651 41853
rect 13707 41797 13793 41853
rect 13849 41797 13935 41853
rect 13991 41797 14077 41853
rect 14133 41797 14219 41853
rect 14275 41797 14361 41853
rect 14417 41797 14503 41853
rect 14559 41797 14645 41853
rect 14701 41797 14787 41853
rect 14843 41797 14853 41853
rect 151 41711 14853 41797
rect 151 41655 161 41711
rect 217 41655 303 41711
rect 359 41655 445 41711
rect 501 41655 587 41711
rect 643 41655 729 41711
rect 785 41655 871 41711
rect 927 41655 1013 41711
rect 1069 41655 1155 41711
rect 1211 41655 1297 41711
rect 1353 41655 1439 41711
rect 1495 41655 1581 41711
rect 1637 41655 1723 41711
rect 1779 41655 1865 41711
rect 1921 41655 2007 41711
rect 2063 41655 2149 41711
rect 2205 41655 2291 41711
rect 2347 41655 2433 41711
rect 2489 41655 2575 41711
rect 2631 41655 2717 41711
rect 2773 41655 2859 41711
rect 2915 41655 3001 41711
rect 3057 41655 3143 41711
rect 3199 41655 3285 41711
rect 3341 41655 3427 41711
rect 3483 41655 3569 41711
rect 3625 41655 3711 41711
rect 3767 41655 3853 41711
rect 3909 41655 3995 41711
rect 4051 41655 4137 41711
rect 4193 41655 4279 41711
rect 4335 41655 4421 41711
rect 4477 41655 4563 41711
rect 4619 41655 4705 41711
rect 4761 41655 4847 41711
rect 4903 41655 4989 41711
rect 5045 41655 5131 41711
rect 5187 41655 5273 41711
rect 5329 41655 5415 41711
rect 5471 41655 5557 41711
rect 5613 41655 5699 41711
rect 5755 41655 5841 41711
rect 5897 41655 5983 41711
rect 6039 41655 6125 41711
rect 6181 41655 6267 41711
rect 6323 41655 6409 41711
rect 6465 41655 6551 41711
rect 6607 41655 6693 41711
rect 6749 41655 6835 41711
rect 6891 41655 6977 41711
rect 7033 41655 7119 41711
rect 7175 41655 7261 41711
rect 7317 41655 7403 41711
rect 7459 41655 7545 41711
rect 7601 41655 7687 41711
rect 7743 41655 7829 41711
rect 7885 41655 7971 41711
rect 8027 41655 8113 41711
rect 8169 41655 8255 41711
rect 8311 41655 8397 41711
rect 8453 41655 8539 41711
rect 8595 41655 8681 41711
rect 8737 41655 8823 41711
rect 8879 41655 8965 41711
rect 9021 41655 9107 41711
rect 9163 41655 9249 41711
rect 9305 41655 9391 41711
rect 9447 41655 9533 41711
rect 9589 41655 9675 41711
rect 9731 41655 9817 41711
rect 9873 41655 9959 41711
rect 10015 41655 10101 41711
rect 10157 41655 10243 41711
rect 10299 41655 10385 41711
rect 10441 41655 10527 41711
rect 10583 41655 10669 41711
rect 10725 41655 10811 41711
rect 10867 41655 10953 41711
rect 11009 41655 11095 41711
rect 11151 41655 11237 41711
rect 11293 41655 11379 41711
rect 11435 41655 11521 41711
rect 11577 41655 11663 41711
rect 11719 41655 11805 41711
rect 11861 41655 11947 41711
rect 12003 41655 12089 41711
rect 12145 41655 12231 41711
rect 12287 41655 12373 41711
rect 12429 41655 12515 41711
rect 12571 41655 12657 41711
rect 12713 41655 12799 41711
rect 12855 41655 12941 41711
rect 12997 41655 13083 41711
rect 13139 41655 13225 41711
rect 13281 41655 13367 41711
rect 13423 41655 13509 41711
rect 13565 41655 13651 41711
rect 13707 41655 13793 41711
rect 13849 41655 13935 41711
rect 13991 41655 14077 41711
rect 14133 41655 14219 41711
rect 14275 41655 14361 41711
rect 14417 41655 14503 41711
rect 14559 41655 14645 41711
rect 14701 41655 14787 41711
rect 14843 41655 14853 41711
rect 151 41569 14853 41655
rect 151 41513 161 41569
rect 217 41513 303 41569
rect 359 41513 445 41569
rect 501 41513 587 41569
rect 643 41513 729 41569
rect 785 41513 871 41569
rect 927 41513 1013 41569
rect 1069 41513 1155 41569
rect 1211 41513 1297 41569
rect 1353 41513 1439 41569
rect 1495 41513 1581 41569
rect 1637 41513 1723 41569
rect 1779 41513 1865 41569
rect 1921 41513 2007 41569
rect 2063 41513 2149 41569
rect 2205 41513 2291 41569
rect 2347 41513 2433 41569
rect 2489 41513 2575 41569
rect 2631 41513 2717 41569
rect 2773 41513 2859 41569
rect 2915 41513 3001 41569
rect 3057 41513 3143 41569
rect 3199 41513 3285 41569
rect 3341 41513 3427 41569
rect 3483 41513 3569 41569
rect 3625 41513 3711 41569
rect 3767 41513 3853 41569
rect 3909 41513 3995 41569
rect 4051 41513 4137 41569
rect 4193 41513 4279 41569
rect 4335 41513 4421 41569
rect 4477 41513 4563 41569
rect 4619 41513 4705 41569
rect 4761 41513 4847 41569
rect 4903 41513 4989 41569
rect 5045 41513 5131 41569
rect 5187 41513 5273 41569
rect 5329 41513 5415 41569
rect 5471 41513 5557 41569
rect 5613 41513 5699 41569
rect 5755 41513 5841 41569
rect 5897 41513 5983 41569
rect 6039 41513 6125 41569
rect 6181 41513 6267 41569
rect 6323 41513 6409 41569
rect 6465 41513 6551 41569
rect 6607 41513 6693 41569
rect 6749 41513 6835 41569
rect 6891 41513 6977 41569
rect 7033 41513 7119 41569
rect 7175 41513 7261 41569
rect 7317 41513 7403 41569
rect 7459 41513 7545 41569
rect 7601 41513 7687 41569
rect 7743 41513 7829 41569
rect 7885 41513 7971 41569
rect 8027 41513 8113 41569
rect 8169 41513 8255 41569
rect 8311 41513 8397 41569
rect 8453 41513 8539 41569
rect 8595 41513 8681 41569
rect 8737 41513 8823 41569
rect 8879 41513 8965 41569
rect 9021 41513 9107 41569
rect 9163 41513 9249 41569
rect 9305 41513 9391 41569
rect 9447 41513 9533 41569
rect 9589 41513 9675 41569
rect 9731 41513 9817 41569
rect 9873 41513 9959 41569
rect 10015 41513 10101 41569
rect 10157 41513 10243 41569
rect 10299 41513 10385 41569
rect 10441 41513 10527 41569
rect 10583 41513 10669 41569
rect 10725 41513 10811 41569
rect 10867 41513 10953 41569
rect 11009 41513 11095 41569
rect 11151 41513 11237 41569
rect 11293 41513 11379 41569
rect 11435 41513 11521 41569
rect 11577 41513 11663 41569
rect 11719 41513 11805 41569
rect 11861 41513 11947 41569
rect 12003 41513 12089 41569
rect 12145 41513 12231 41569
rect 12287 41513 12373 41569
rect 12429 41513 12515 41569
rect 12571 41513 12657 41569
rect 12713 41513 12799 41569
rect 12855 41513 12941 41569
rect 12997 41513 13083 41569
rect 13139 41513 13225 41569
rect 13281 41513 13367 41569
rect 13423 41513 13509 41569
rect 13565 41513 13651 41569
rect 13707 41513 13793 41569
rect 13849 41513 13935 41569
rect 13991 41513 14077 41569
rect 14133 41513 14219 41569
rect 14275 41513 14361 41569
rect 14417 41513 14503 41569
rect 14559 41513 14645 41569
rect 14701 41513 14787 41569
rect 14843 41513 14853 41569
rect 151 41427 14853 41513
rect 151 41371 161 41427
rect 217 41371 303 41427
rect 359 41371 445 41427
rect 501 41371 587 41427
rect 643 41371 729 41427
rect 785 41371 871 41427
rect 927 41371 1013 41427
rect 1069 41371 1155 41427
rect 1211 41371 1297 41427
rect 1353 41371 1439 41427
rect 1495 41371 1581 41427
rect 1637 41371 1723 41427
rect 1779 41371 1865 41427
rect 1921 41371 2007 41427
rect 2063 41371 2149 41427
rect 2205 41371 2291 41427
rect 2347 41371 2433 41427
rect 2489 41371 2575 41427
rect 2631 41371 2717 41427
rect 2773 41371 2859 41427
rect 2915 41371 3001 41427
rect 3057 41371 3143 41427
rect 3199 41371 3285 41427
rect 3341 41371 3427 41427
rect 3483 41371 3569 41427
rect 3625 41371 3711 41427
rect 3767 41371 3853 41427
rect 3909 41371 3995 41427
rect 4051 41371 4137 41427
rect 4193 41371 4279 41427
rect 4335 41371 4421 41427
rect 4477 41371 4563 41427
rect 4619 41371 4705 41427
rect 4761 41371 4847 41427
rect 4903 41371 4989 41427
rect 5045 41371 5131 41427
rect 5187 41371 5273 41427
rect 5329 41371 5415 41427
rect 5471 41371 5557 41427
rect 5613 41371 5699 41427
rect 5755 41371 5841 41427
rect 5897 41371 5983 41427
rect 6039 41371 6125 41427
rect 6181 41371 6267 41427
rect 6323 41371 6409 41427
rect 6465 41371 6551 41427
rect 6607 41371 6693 41427
rect 6749 41371 6835 41427
rect 6891 41371 6977 41427
rect 7033 41371 7119 41427
rect 7175 41371 7261 41427
rect 7317 41371 7403 41427
rect 7459 41371 7545 41427
rect 7601 41371 7687 41427
rect 7743 41371 7829 41427
rect 7885 41371 7971 41427
rect 8027 41371 8113 41427
rect 8169 41371 8255 41427
rect 8311 41371 8397 41427
rect 8453 41371 8539 41427
rect 8595 41371 8681 41427
rect 8737 41371 8823 41427
rect 8879 41371 8965 41427
rect 9021 41371 9107 41427
rect 9163 41371 9249 41427
rect 9305 41371 9391 41427
rect 9447 41371 9533 41427
rect 9589 41371 9675 41427
rect 9731 41371 9817 41427
rect 9873 41371 9959 41427
rect 10015 41371 10101 41427
rect 10157 41371 10243 41427
rect 10299 41371 10385 41427
rect 10441 41371 10527 41427
rect 10583 41371 10669 41427
rect 10725 41371 10811 41427
rect 10867 41371 10953 41427
rect 11009 41371 11095 41427
rect 11151 41371 11237 41427
rect 11293 41371 11379 41427
rect 11435 41371 11521 41427
rect 11577 41371 11663 41427
rect 11719 41371 11805 41427
rect 11861 41371 11947 41427
rect 12003 41371 12089 41427
rect 12145 41371 12231 41427
rect 12287 41371 12373 41427
rect 12429 41371 12515 41427
rect 12571 41371 12657 41427
rect 12713 41371 12799 41427
rect 12855 41371 12941 41427
rect 12997 41371 13083 41427
rect 13139 41371 13225 41427
rect 13281 41371 13367 41427
rect 13423 41371 13509 41427
rect 13565 41371 13651 41427
rect 13707 41371 13793 41427
rect 13849 41371 13935 41427
rect 13991 41371 14077 41427
rect 14133 41371 14219 41427
rect 14275 41371 14361 41427
rect 14417 41371 14503 41427
rect 14559 41371 14645 41427
rect 14701 41371 14787 41427
rect 14843 41371 14853 41427
rect 151 41285 14853 41371
rect 151 41229 161 41285
rect 217 41229 303 41285
rect 359 41229 445 41285
rect 501 41229 587 41285
rect 643 41229 729 41285
rect 785 41229 871 41285
rect 927 41229 1013 41285
rect 1069 41229 1155 41285
rect 1211 41229 1297 41285
rect 1353 41229 1439 41285
rect 1495 41229 1581 41285
rect 1637 41229 1723 41285
rect 1779 41229 1865 41285
rect 1921 41229 2007 41285
rect 2063 41229 2149 41285
rect 2205 41229 2291 41285
rect 2347 41229 2433 41285
rect 2489 41229 2575 41285
rect 2631 41229 2717 41285
rect 2773 41229 2859 41285
rect 2915 41229 3001 41285
rect 3057 41229 3143 41285
rect 3199 41229 3285 41285
rect 3341 41229 3427 41285
rect 3483 41229 3569 41285
rect 3625 41229 3711 41285
rect 3767 41229 3853 41285
rect 3909 41229 3995 41285
rect 4051 41229 4137 41285
rect 4193 41229 4279 41285
rect 4335 41229 4421 41285
rect 4477 41229 4563 41285
rect 4619 41229 4705 41285
rect 4761 41229 4847 41285
rect 4903 41229 4989 41285
rect 5045 41229 5131 41285
rect 5187 41229 5273 41285
rect 5329 41229 5415 41285
rect 5471 41229 5557 41285
rect 5613 41229 5699 41285
rect 5755 41229 5841 41285
rect 5897 41229 5983 41285
rect 6039 41229 6125 41285
rect 6181 41229 6267 41285
rect 6323 41229 6409 41285
rect 6465 41229 6551 41285
rect 6607 41229 6693 41285
rect 6749 41229 6835 41285
rect 6891 41229 6977 41285
rect 7033 41229 7119 41285
rect 7175 41229 7261 41285
rect 7317 41229 7403 41285
rect 7459 41229 7545 41285
rect 7601 41229 7687 41285
rect 7743 41229 7829 41285
rect 7885 41229 7971 41285
rect 8027 41229 8113 41285
rect 8169 41229 8255 41285
rect 8311 41229 8397 41285
rect 8453 41229 8539 41285
rect 8595 41229 8681 41285
rect 8737 41229 8823 41285
rect 8879 41229 8965 41285
rect 9021 41229 9107 41285
rect 9163 41229 9249 41285
rect 9305 41229 9391 41285
rect 9447 41229 9533 41285
rect 9589 41229 9675 41285
rect 9731 41229 9817 41285
rect 9873 41229 9959 41285
rect 10015 41229 10101 41285
rect 10157 41229 10243 41285
rect 10299 41229 10385 41285
rect 10441 41229 10527 41285
rect 10583 41229 10669 41285
rect 10725 41229 10811 41285
rect 10867 41229 10953 41285
rect 11009 41229 11095 41285
rect 11151 41229 11237 41285
rect 11293 41229 11379 41285
rect 11435 41229 11521 41285
rect 11577 41229 11663 41285
rect 11719 41229 11805 41285
rect 11861 41229 11947 41285
rect 12003 41229 12089 41285
rect 12145 41229 12231 41285
rect 12287 41229 12373 41285
rect 12429 41229 12515 41285
rect 12571 41229 12657 41285
rect 12713 41229 12799 41285
rect 12855 41229 12941 41285
rect 12997 41229 13083 41285
rect 13139 41229 13225 41285
rect 13281 41229 13367 41285
rect 13423 41229 13509 41285
rect 13565 41229 13651 41285
rect 13707 41229 13793 41285
rect 13849 41229 13935 41285
rect 13991 41229 14077 41285
rect 14133 41229 14219 41285
rect 14275 41229 14361 41285
rect 14417 41229 14503 41285
rect 14559 41229 14645 41285
rect 14701 41229 14787 41285
rect 14843 41229 14853 41285
rect 151 41219 14853 41229
rect 151 40963 14853 40973
rect 151 40907 161 40963
rect 217 40907 303 40963
rect 359 40907 445 40963
rect 501 40907 587 40963
rect 643 40907 729 40963
rect 785 40907 871 40963
rect 927 40907 1013 40963
rect 1069 40907 1155 40963
rect 1211 40907 1297 40963
rect 1353 40907 1439 40963
rect 1495 40907 1581 40963
rect 1637 40907 1723 40963
rect 1779 40907 1865 40963
rect 1921 40907 2007 40963
rect 2063 40907 2149 40963
rect 2205 40907 2291 40963
rect 2347 40907 2433 40963
rect 2489 40907 2575 40963
rect 2631 40907 2717 40963
rect 2773 40907 2859 40963
rect 2915 40907 3001 40963
rect 3057 40907 3143 40963
rect 3199 40907 3285 40963
rect 3341 40907 3427 40963
rect 3483 40907 3569 40963
rect 3625 40907 3711 40963
rect 3767 40907 3853 40963
rect 3909 40907 3995 40963
rect 4051 40907 4137 40963
rect 4193 40907 4279 40963
rect 4335 40907 4421 40963
rect 4477 40907 4563 40963
rect 4619 40907 4705 40963
rect 4761 40907 4847 40963
rect 4903 40907 4989 40963
rect 5045 40907 5131 40963
rect 5187 40907 5273 40963
rect 5329 40907 5415 40963
rect 5471 40907 5557 40963
rect 5613 40907 5699 40963
rect 5755 40907 5841 40963
rect 5897 40907 5983 40963
rect 6039 40907 6125 40963
rect 6181 40907 6267 40963
rect 6323 40907 6409 40963
rect 6465 40907 6551 40963
rect 6607 40907 6693 40963
rect 6749 40907 6835 40963
rect 6891 40907 6977 40963
rect 7033 40907 7119 40963
rect 7175 40907 7261 40963
rect 7317 40907 7403 40963
rect 7459 40907 7545 40963
rect 7601 40907 7687 40963
rect 7743 40907 7829 40963
rect 7885 40907 7971 40963
rect 8027 40907 8113 40963
rect 8169 40907 8255 40963
rect 8311 40907 8397 40963
rect 8453 40907 8539 40963
rect 8595 40907 8681 40963
rect 8737 40907 8823 40963
rect 8879 40907 8965 40963
rect 9021 40907 9107 40963
rect 9163 40907 9249 40963
rect 9305 40907 9391 40963
rect 9447 40907 9533 40963
rect 9589 40907 9675 40963
rect 9731 40907 9817 40963
rect 9873 40907 9959 40963
rect 10015 40907 10101 40963
rect 10157 40907 10243 40963
rect 10299 40907 10385 40963
rect 10441 40907 10527 40963
rect 10583 40907 10669 40963
rect 10725 40907 10811 40963
rect 10867 40907 10953 40963
rect 11009 40907 11095 40963
rect 11151 40907 11237 40963
rect 11293 40907 11379 40963
rect 11435 40907 11521 40963
rect 11577 40907 11663 40963
rect 11719 40907 11805 40963
rect 11861 40907 11947 40963
rect 12003 40907 12089 40963
rect 12145 40907 12231 40963
rect 12287 40907 12373 40963
rect 12429 40907 12515 40963
rect 12571 40907 12657 40963
rect 12713 40907 12799 40963
rect 12855 40907 12941 40963
rect 12997 40907 13083 40963
rect 13139 40907 13225 40963
rect 13281 40907 13367 40963
rect 13423 40907 13509 40963
rect 13565 40907 13651 40963
rect 13707 40907 13793 40963
rect 13849 40907 13935 40963
rect 13991 40907 14077 40963
rect 14133 40907 14219 40963
rect 14275 40907 14361 40963
rect 14417 40907 14503 40963
rect 14559 40907 14645 40963
rect 14701 40907 14787 40963
rect 14843 40907 14853 40963
rect 151 40821 14853 40907
rect 151 40765 161 40821
rect 217 40765 303 40821
rect 359 40765 445 40821
rect 501 40765 587 40821
rect 643 40765 729 40821
rect 785 40765 871 40821
rect 927 40765 1013 40821
rect 1069 40765 1155 40821
rect 1211 40765 1297 40821
rect 1353 40765 1439 40821
rect 1495 40765 1581 40821
rect 1637 40765 1723 40821
rect 1779 40765 1865 40821
rect 1921 40765 2007 40821
rect 2063 40765 2149 40821
rect 2205 40765 2291 40821
rect 2347 40765 2433 40821
rect 2489 40765 2575 40821
rect 2631 40765 2717 40821
rect 2773 40765 2859 40821
rect 2915 40765 3001 40821
rect 3057 40765 3143 40821
rect 3199 40765 3285 40821
rect 3341 40765 3427 40821
rect 3483 40765 3569 40821
rect 3625 40765 3711 40821
rect 3767 40765 3853 40821
rect 3909 40765 3995 40821
rect 4051 40765 4137 40821
rect 4193 40765 4279 40821
rect 4335 40765 4421 40821
rect 4477 40765 4563 40821
rect 4619 40765 4705 40821
rect 4761 40765 4847 40821
rect 4903 40765 4989 40821
rect 5045 40765 5131 40821
rect 5187 40765 5273 40821
rect 5329 40765 5415 40821
rect 5471 40765 5557 40821
rect 5613 40765 5699 40821
rect 5755 40765 5841 40821
rect 5897 40765 5983 40821
rect 6039 40765 6125 40821
rect 6181 40765 6267 40821
rect 6323 40765 6409 40821
rect 6465 40765 6551 40821
rect 6607 40765 6693 40821
rect 6749 40765 6835 40821
rect 6891 40765 6977 40821
rect 7033 40765 7119 40821
rect 7175 40765 7261 40821
rect 7317 40765 7403 40821
rect 7459 40765 7545 40821
rect 7601 40765 7687 40821
rect 7743 40765 7829 40821
rect 7885 40765 7971 40821
rect 8027 40765 8113 40821
rect 8169 40765 8255 40821
rect 8311 40765 8397 40821
rect 8453 40765 8539 40821
rect 8595 40765 8681 40821
rect 8737 40765 8823 40821
rect 8879 40765 8965 40821
rect 9021 40765 9107 40821
rect 9163 40765 9249 40821
rect 9305 40765 9391 40821
rect 9447 40765 9533 40821
rect 9589 40765 9675 40821
rect 9731 40765 9817 40821
rect 9873 40765 9959 40821
rect 10015 40765 10101 40821
rect 10157 40765 10243 40821
rect 10299 40765 10385 40821
rect 10441 40765 10527 40821
rect 10583 40765 10669 40821
rect 10725 40765 10811 40821
rect 10867 40765 10953 40821
rect 11009 40765 11095 40821
rect 11151 40765 11237 40821
rect 11293 40765 11379 40821
rect 11435 40765 11521 40821
rect 11577 40765 11663 40821
rect 11719 40765 11805 40821
rect 11861 40765 11947 40821
rect 12003 40765 12089 40821
rect 12145 40765 12231 40821
rect 12287 40765 12373 40821
rect 12429 40765 12515 40821
rect 12571 40765 12657 40821
rect 12713 40765 12799 40821
rect 12855 40765 12941 40821
rect 12997 40765 13083 40821
rect 13139 40765 13225 40821
rect 13281 40765 13367 40821
rect 13423 40765 13509 40821
rect 13565 40765 13651 40821
rect 13707 40765 13793 40821
rect 13849 40765 13935 40821
rect 13991 40765 14077 40821
rect 14133 40765 14219 40821
rect 14275 40765 14361 40821
rect 14417 40765 14503 40821
rect 14559 40765 14645 40821
rect 14701 40765 14787 40821
rect 14843 40765 14853 40821
rect 151 40679 14853 40765
rect 151 40623 161 40679
rect 217 40623 303 40679
rect 359 40623 445 40679
rect 501 40623 587 40679
rect 643 40623 729 40679
rect 785 40623 871 40679
rect 927 40623 1013 40679
rect 1069 40623 1155 40679
rect 1211 40623 1297 40679
rect 1353 40623 1439 40679
rect 1495 40623 1581 40679
rect 1637 40623 1723 40679
rect 1779 40623 1865 40679
rect 1921 40623 2007 40679
rect 2063 40623 2149 40679
rect 2205 40623 2291 40679
rect 2347 40623 2433 40679
rect 2489 40623 2575 40679
rect 2631 40623 2717 40679
rect 2773 40623 2859 40679
rect 2915 40623 3001 40679
rect 3057 40623 3143 40679
rect 3199 40623 3285 40679
rect 3341 40623 3427 40679
rect 3483 40623 3569 40679
rect 3625 40623 3711 40679
rect 3767 40623 3853 40679
rect 3909 40623 3995 40679
rect 4051 40623 4137 40679
rect 4193 40623 4279 40679
rect 4335 40623 4421 40679
rect 4477 40623 4563 40679
rect 4619 40623 4705 40679
rect 4761 40623 4847 40679
rect 4903 40623 4989 40679
rect 5045 40623 5131 40679
rect 5187 40623 5273 40679
rect 5329 40623 5415 40679
rect 5471 40623 5557 40679
rect 5613 40623 5699 40679
rect 5755 40623 5841 40679
rect 5897 40623 5983 40679
rect 6039 40623 6125 40679
rect 6181 40623 6267 40679
rect 6323 40623 6409 40679
rect 6465 40623 6551 40679
rect 6607 40623 6693 40679
rect 6749 40623 6835 40679
rect 6891 40623 6977 40679
rect 7033 40623 7119 40679
rect 7175 40623 7261 40679
rect 7317 40623 7403 40679
rect 7459 40623 7545 40679
rect 7601 40623 7687 40679
rect 7743 40623 7829 40679
rect 7885 40623 7971 40679
rect 8027 40623 8113 40679
rect 8169 40623 8255 40679
rect 8311 40623 8397 40679
rect 8453 40623 8539 40679
rect 8595 40623 8681 40679
rect 8737 40623 8823 40679
rect 8879 40623 8965 40679
rect 9021 40623 9107 40679
rect 9163 40623 9249 40679
rect 9305 40623 9391 40679
rect 9447 40623 9533 40679
rect 9589 40623 9675 40679
rect 9731 40623 9817 40679
rect 9873 40623 9959 40679
rect 10015 40623 10101 40679
rect 10157 40623 10243 40679
rect 10299 40623 10385 40679
rect 10441 40623 10527 40679
rect 10583 40623 10669 40679
rect 10725 40623 10811 40679
rect 10867 40623 10953 40679
rect 11009 40623 11095 40679
rect 11151 40623 11237 40679
rect 11293 40623 11379 40679
rect 11435 40623 11521 40679
rect 11577 40623 11663 40679
rect 11719 40623 11805 40679
rect 11861 40623 11947 40679
rect 12003 40623 12089 40679
rect 12145 40623 12231 40679
rect 12287 40623 12373 40679
rect 12429 40623 12515 40679
rect 12571 40623 12657 40679
rect 12713 40623 12799 40679
rect 12855 40623 12941 40679
rect 12997 40623 13083 40679
rect 13139 40623 13225 40679
rect 13281 40623 13367 40679
rect 13423 40623 13509 40679
rect 13565 40623 13651 40679
rect 13707 40623 13793 40679
rect 13849 40623 13935 40679
rect 13991 40623 14077 40679
rect 14133 40623 14219 40679
rect 14275 40623 14361 40679
rect 14417 40623 14503 40679
rect 14559 40623 14645 40679
rect 14701 40623 14787 40679
rect 14843 40623 14853 40679
rect 151 40537 14853 40623
rect 151 40481 161 40537
rect 217 40481 303 40537
rect 359 40481 445 40537
rect 501 40481 587 40537
rect 643 40481 729 40537
rect 785 40481 871 40537
rect 927 40481 1013 40537
rect 1069 40481 1155 40537
rect 1211 40481 1297 40537
rect 1353 40481 1439 40537
rect 1495 40481 1581 40537
rect 1637 40481 1723 40537
rect 1779 40481 1865 40537
rect 1921 40481 2007 40537
rect 2063 40481 2149 40537
rect 2205 40481 2291 40537
rect 2347 40481 2433 40537
rect 2489 40481 2575 40537
rect 2631 40481 2717 40537
rect 2773 40481 2859 40537
rect 2915 40481 3001 40537
rect 3057 40481 3143 40537
rect 3199 40481 3285 40537
rect 3341 40481 3427 40537
rect 3483 40481 3569 40537
rect 3625 40481 3711 40537
rect 3767 40481 3853 40537
rect 3909 40481 3995 40537
rect 4051 40481 4137 40537
rect 4193 40481 4279 40537
rect 4335 40481 4421 40537
rect 4477 40481 4563 40537
rect 4619 40481 4705 40537
rect 4761 40481 4847 40537
rect 4903 40481 4989 40537
rect 5045 40481 5131 40537
rect 5187 40481 5273 40537
rect 5329 40481 5415 40537
rect 5471 40481 5557 40537
rect 5613 40481 5699 40537
rect 5755 40481 5841 40537
rect 5897 40481 5983 40537
rect 6039 40481 6125 40537
rect 6181 40481 6267 40537
rect 6323 40481 6409 40537
rect 6465 40481 6551 40537
rect 6607 40481 6693 40537
rect 6749 40481 6835 40537
rect 6891 40481 6977 40537
rect 7033 40481 7119 40537
rect 7175 40481 7261 40537
rect 7317 40481 7403 40537
rect 7459 40481 7545 40537
rect 7601 40481 7687 40537
rect 7743 40481 7829 40537
rect 7885 40481 7971 40537
rect 8027 40481 8113 40537
rect 8169 40481 8255 40537
rect 8311 40481 8397 40537
rect 8453 40481 8539 40537
rect 8595 40481 8681 40537
rect 8737 40481 8823 40537
rect 8879 40481 8965 40537
rect 9021 40481 9107 40537
rect 9163 40481 9249 40537
rect 9305 40481 9391 40537
rect 9447 40481 9533 40537
rect 9589 40481 9675 40537
rect 9731 40481 9817 40537
rect 9873 40481 9959 40537
rect 10015 40481 10101 40537
rect 10157 40481 10243 40537
rect 10299 40481 10385 40537
rect 10441 40481 10527 40537
rect 10583 40481 10669 40537
rect 10725 40481 10811 40537
rect 10867 40481 10953 40537
rect 11009 40481 11095 40537
rect 11151 40481 11237 40537
rect 11293 40481 11379 40537
rect 11435 40481 11521 40537
rect 11577 40481 11663 40537
rect 11719 40481 11805 40537
rect 11861 40481 11947 40537
rect 12003 40481 12089 40537
rect 12145 40481 12231 40537
rect 12287 40481 12373 40537
rect 12429 40481 12515 40537
rect 12571 40481 12657 40537
rect 12713 40481 12799 40537
rect 12855 40481 12941 40537
rect 12997 40481 13083 40537
rect 13139 40481 13225 40537
rect 13281 40481 13367 40537
rect 13423 40481 13509 40537
rect 13565 40481 13651 40537
rect 13707 40481 13793 40537
rect 13849 40481 13935 40537
rect 13991 40481 14077 40537
rect 14133 40481 14219 40537
rect 14275 40481 14361 40537
rect 14417 40481 14503 40537
rect 14559 40481 14645 40537
rect 14701 40481 14787 40537
rect 14843 40481 14853 40537
rect 151 40395 14853 40481
rect 151 40339 161 40395
rect 217 40339 303 40395
rect 359 40339 445 40395
rect 501 40339 587 40395
rect 643 40339 729 40395
rect 785 40339 871 40395
rect 927 40339 1013 40395
rect 1069 40339 1155 40395
rect 1211 40339 1297 40395
rect 1353 40339 1439 40395
rect 1495 40339 1581 40395
rect 1637 40339 1723 40395
rect 1779 40339 1865 40395
rect 1921 40339 2007 40395
rect 2063 40339 2149 40395
rect 2205 40339 2291 40395
rect 2347 40339 2433 40395
rect 2489 40339 2575 40395
rect 2631 40339 2717 40395
rect 2773 40339 2859 40395
rect 2915 40339 3001 40395
rect 3057 40339 3143 40395
rect 3199 40339 3285 40395
rect 3341 40339 3427 40395
rect 3483 40339 3569 40395
rect 3625 40339 3711 40395
rect 3767 40339 3853 40395
rect 3909 40339 3995 40395
rect 4051 40339 4137 40395
rect 4193 40339 4279 40395
rect 4335 40339 4421 40395
rect 4477 40339 4563 40395
rect 4619 40339 4705 40395
rect 4761 40339 4847 40395
rect 4903 40339 4989 40395
rect 5045 40339 5131 40395
rect 5187 40339 5273 40395
rect 5329 40339 5415 40395
rect 5471 40339 5557 40395
rect 5613 40339 5699 40395
rect 5755 40339 5841 40395
rect 5897 40339 5983 40395
rect 6039 40339 6125 40395
rect 6181 40339 6267 40395
rect 6323 40339 6409 40395
rect 6465 40339 6551 40395
rect 6607 40339 6693 40395
rect 6749 40339 6835 40395
rect 6891 40339 6977 40395
rect 7033 40339 7119 40395
rect 7175 40339 7261 40395
rect 7317 40339 7403 40395
rect 7459 40339 7545 40395
rect 7601 40339 7687 40395
rect 7743 40339 7829 40395
rect 7885 40339 7971 40395
rect 8027 40339 8113 40395
rect 8169 40339 8255 40395
rect 8311 40339 8397 40395
rect 8453 40339 8539 40395
rect 8595 40339 8681 40395
rect 8737 40339 8823 40395
rect 8879 40339 8965 40395
rect 9021 40339 9107 40395
rect 9163 40339 9249 40395
rect 9305 40339 9391 40395
rect 9447 40339 9533 40395
rect 9589 40339 9675 40395
rect 9731 40339 9817 40395
rect 9873 40339 9959 40395
rect 10015 40339 10101 40395
rect 10157 40339 10243 40395
rect 10299 40339 10385 40395
rect 10441 40339 10527 40395
rect 10583 40339 10669 40395
rect 10725 40339 10811 40395
rect 10867 40339 10953 40395
rect 11009 40339 11095 40395
rect 11151 40339 11237 40395
rect 11293 40339 11379 40395
rect 11435 40339 11521 40395
rect 11577 40339 11663 40395
rect 11719 40339 11805 40395
rect 11861 40339 11947 40395
rect 12003 40339 12089 40395
rect 12145 40339 12231 40395
rect 12287 40339 12373 40395
rect 12429 40339 12515 40395
rect 12571 40339 12657 40395
rect 12713 40339 12799 40395
rect 12855 40339 12941 40395
rect 12997 40339 13083 40395
rect 13139 40339 13225 40395
rect 13281 40339 13367 40395
rect 13423 40339 13509 40395
rect 13565 40339 13651 40395
rect 13707 40339 13793 40395
rect 13849 40339 13935 40395
rect 13991 40339 14077 40395
rect 14133 40339 14219 40395
rect 14275 40339 14361 40395
rect 14417 40339 14503 40395
rect 14559 40339 14645 40395
rect 14701 40339 14787 40395
rect 14843 40339 14853 40395
rect 151 40253 14853 40339
rect 151 40197 161 40253
rect 217 40197 303 40253
rect 359 40197 445 40253
rect 501 40197 587 40253
rect 643 40197 729 40253
rect 785 40197 871 40253
rect 927 40197 1013 40253
rect 1069 40197 1155 40253
rect 1211 40197 1297 40253
rect 1353 40197 1439 40253
rect 1495 40197 1581 40253
rect 1637 40197 1723 40253
rect 1779 40197 1865 40253
rect 1921 40197 2007 40253
rect 2063 40197 2149 40253
rect 2205 40197 2291 40253
rect 2347 40197 2433 40253
rect 2489 40197 2575 40253
rect 2631 40197 2717 40253
rect 2773 40197 2859 40253
rect 2915 40197 3001 40253
rect 3057 40197 3143 40253
rect 3199 40197 3285 40253
rect 3341 40197 3427 40253
rect 3483 40197 3569 40253
rect 3625 40197 3711 40253
rect 3767 40197 3853 40253
rect 3909 40197 3995 40253
rect 4051 40197 4137 40253
rect 4193 40197 4279 40253
rect 4335 40197 4421 40253
rect 4477 40197 4563 40253
rect 4619 40197 4705 40253
rect 4761 40197 4847 40253
rect 4903 40197 4989 40253
rect 5045 40197 5131 40253
rect 5187 40197 5273 40253
rect 5329 40197 5415 40253
rect 5471 40197 5557 40253
rect 5613 40197 5699 40253
rect 5755 40197 5841 40253
rect 5897 40197 5983 40253
rect 6039 40197 6125 40253
rect 6181 40197 6267 40253
rect 6323 40197 6409 40253
rect 6465 40197 6551 40253
rect 6607 40197 6693 40253
rect 6749 40197 6835 40253
rect 6891 40197 6977 40253
rect 7033 40197 7119 40253
rect 7175 40197 7261 40253
rect 7317 40197 7403 40253
rect 7459 40197 7545 40253
rect 7601 40197 7687 40253
rect 7743 40197 7829 40253
rect 7885 40197 7971 40253
rect 8027 40197 8113 40253
rect 8169 40197 8255 40253
rect 8311 40197 8397 40253
rect 8453 40197 8539 40253
rect 8595 40197 8681 40253
rect 8737 40197 8823 40253
rect 8879 40197 8965 40253
rect 9021 40197 9107 40253
rect 9163 40197 9249 40253
rect 9305 40197 9391 40253
rect 9447 40197 9533 40253
rect 9589 40197 9675 40253
rect 9731 40197 9817 40253
rect 9873 40197 9959 40253
rect 10015 40197 10101 40253
rect 10157 40197 10243 40253
rect 10299 40197 10385 40253
rect 10441 40197 10527 40253
rect 10583 40197 10669 40253
rect 10725 40197 10811 40253
rect 10867 40197 10953 40253
rect 11009 40197 11095 40253
rect 11151 40197 11237 40253
rect 11293 40197 11379 40253
rect 11435 40197 11521 40253
rect 11577 40197 11663 40253
rect 11719 40197 11805 40253
rect 11861 40197 11947 40253
rect 12003 40197 12089 40253
rect 12145 40197 12231 40253
rect 12287 40197 12373 40253
rect 12429 40197 12515 40253
rect 12571 40197 12657 40253
rect 12713 40197 12799 40253
rect 12855 40197 12941 40253
rect 12997 40197 13083 40253
rect 13139 40197 13225 40253
rect 13281 40197 13367 40253
rect 13423 40197 13509 40253
rect 13565 40197 13651 40253
rect 13707 40197 13793 40253
rect 13849 40197 13935 40253
rect 13991 40197 14077 40253
rect 14133 40197 14219 40253
rect 14275 40197 14361 40253
rect 14417 40197 14503 40253
rect 14559 40197 14645 40253
rect 14701 40197 14787 40253
rect 14843 40197 14853 40253
rect 151 40111 14853 40197
rect 151 40055 161 40111
rect 217 40055 303 40111
rect 359 40055 445 40111
rect 501 40055 587 40111
rect 643 40055 729 40111
rect 785 40055 871 40111
rect 927 40055 1013 40111
rect 1069 40055 1155 40111
rect 1211 40055 1297 40111
rect 1353 40055 1439 40111
rect 1495 40055 1581 40111
rect 1637 40055 1723 40111
rect 1779 40055 1865 40111
rect 1921 40055 2007 40111
rect 2063 40055 2149 40111
rect 2205 40055 2291 40111
rect 2347 40055 2433 40111
rect 2489 40055 2575 40111
rect 2631 40055 2717 40111
rect 2773 40055 2859 40111
rect 2915 40055 3001 40111
rect 3057 40055 3143 40111
rect 3199 40055 3285 40111
rect 3341 40055 3427 40111
rect 3483 40055 3569 40111
rect 3625 40055 3711 40111
rect 3767 40055 3853 40111
rect 3909 40055 3995 40111
rect 4051 40055 4137 40111
rect 4193 40055 4279 40111
rect 4335 40055 4421 40111
rect 4477 40055 4563 40111
rect 4619 40055 4705 40111
rect 4761 40055 4847 40111
rect 4903 40055 4989 40111
rect 5045 40055 5131 40111
rect 5187 40055 5273 40111
rect 5329 40055 5415 40111
rect 5471 40055 5557 40111
rect 5613 40055 5699 40111
rect 5755 40055 5841 40111
rect 5897 40055 5983 40111
rect 6039 40055 6125 40111
rect 6181 40055 6267 40111
rect 6323 40055 6409 40111
rect 6465 40055 6551 40111
rect 6607 40055 6693 40111
rect 6749 40055 6835 40111
rect 6891 40055 6977 40111
rect 7033 40055 7119 40111
rect 7175 40055 7261 40111
rect 7317 40055 7403 40111
rect 7459 40055 7545 40111
rect 7601 40055 7687 40111
rect 7743 40055 7829 40111
rect 7885 40055 7971 40111
rect 8027 40055 8113 40111
rect 8169 40055 8255 40111
rect 8311 40055 8397 40111
rect 8453 40055 8539 40111
rect 8595 40055 8681 40111
rect 8737 40055 8823 40111
rect 8879 40055 8965 40111
rect 9021 40055 9107 40111
rect 9163 40055 9249 40111
rect 9305 40055 9391 40111
rect 9447 40055 9533 40111
rect 9589 40055 9675 40111
rect 9731 40055 9817 40111
rect 9873 40055 9959 40111
rect 10015 40055 10101 40111
rect 10157 40055 10243 40111
rect 10299 40055 10385 40111
rect 10441 40055 10527 40111
rect 10583 40055 10669 40111
rect 10725 40055 10811 40111
rect 10867 40055 10953 40111
rect 11009 40055 11095 40111
rect 11151 40055 11237 40111
rect 11293 40055 11379 40111
rect 11435 40055 11521 40111
rect 11577 40055 11663 40111
rect 11719 40055 11805 40111
rect 11861 40055 11947 40111
rect 12003 40055 12089 40111
rect 12145 40055 12231 40111
rect 12287 40055 12373 40111
rect 12429 40055 12515 40111
rect 12571 40055 12657 40111
rect 12713 40055 12799 40111
rect 12855 40055 12941 40111
rect 12997 40055 13083 40111
rect 13139 40055 13225 40111
rect 13281 40055 13367 40111
rect 13423 40055 13509 40111
rect 13565 40055 13651 40111
rect 13707 40055 13793 40111
rect 13849 40055 13935 40111
rect 13991 40055 14077 40111
rect 14133 40055 14219 40111
rect 14275 40055 14361 40111
rect 14417 40055 14503 40111
rect 14559 40055 14645 40111
rect 14701 40055 14787 40111
rect 14843 40055 14853 40111
rect 151 39969 14853 40055
rect 151 39913 161 39969
rect 217 39913 303 39969
rect 359 39913 445 39969
rect 501 39913 587 39969
rect 643 39913 729 39969
rect 785 39913 871 39969
rect 927 39913 1013 39969
rect 1069 39913 1155 39969
rect 1211 39913 1297 39969
rect 1353 39913 1439 39969
rect 1495 39913 1581 39969
rect 1637 39913 1723 39969
rect 1779 39913 1865 39969
rect 1921 39913 2007 39969
rect 2063 39913 2149 39969
rect 2205 39913 2291 39969
rect 2347 39913 2433 39969
rect 2489 39913 2575 39969
rect 2631 39913 2717 39969
rect 2773 39913 2859 39969
rect 2915 39913 3001 39969
rect 3057 39913 3143 39969
rect 3199 39913 3285 39969
rect 3341 39913 3427 39969
rect 3483 39913 3569 39969
rect 3625 39913 3711 39969
rect 3767 39913 3853 39969
rect 3909 39913 3995 39969
rect 4051 39913 4137 39969
rect 4193 39913 4279 39969
rect 4335 39913 4421 39969
rect 4477 39913 4563 39969
rect 4619 39913 4705 39969
rect 4761 39913 4847 39969
rect 4903 39913 4989 39969
rect 5045 39913 5131 39969
rect 5187 39913 5273 39969
rect 5329 39913 5415 39969
rect 5471 39913 5557 39969
rect 5613 39913 5699 39969
rect 5755 39913 5841 39969
rect 5897 39913 5983 39969
rect 6039 39913 6125 39969
rect 6181 39913 6267 39969
rect 6323 39913 6409 39969
rect 6465 39913 6551 39969
rect 6607 39913 6693 39969
rect 6749 39913 6835 39969
rect 6891 39913 6977 39969
rect 7033 39913 7119 39969
rect 7175 39913 7261 39969
rect 7317 39913 7403 39969
rect 7459 39913 7545 39969
rect 7601 39913 7687 39969
rect 7743 39913 7829 39969
rect 7885 39913 7971 39969
rect 8027 39913 8113 39969
rect 8169 39913 8255 39969
rect 8311 39913 8397 39969
rect 8453 39913 8539 39969
rect 8595 39913 8681 39969
rect 8737 39913 8823 39969
rect 8879 39913 8965 39969
rect 9021 39913 9107 39969
rect 9163 39913 9249 39969
rect 9305 39913 9391 39969
rect 9447 39913 9533 39969
rect 9589 39913 9675 39969
rect 9731 39913 9817 39969
rect 9873 39913 9959 39969
rect 10015 39913 10101 39969
rect 10157 39913 10243 39969
rect 10299 39913 10385 39969
rect 10441 39913 10527 39969
rect 10583 39913 10669 39969
rect 10725 39913 10811 39969
rect 10867 39913 10953 39969
rect 11009 39913 11095 39969
rect 11151 39913 11237 39969
rect 11293 39913 11379 39969
rect 11435 39913 11521 39969
rect 11577 39913 11663 39969
rect 11719 39913 11805 39969
rect 11861 39913 11947 39969
rect 12003 39913 12089 39969
rect 12145 39913 12231 39969
rect 12287 39913 12373 39969
rect 12429 39913 12515 39969
rect 12571 39913 12657 39969
rect 12713 39913 12799 39969
rect 12855 39913 12941 39969
rect 12997 39913 13083 39969
rect 13139 39913 13225 39969
rect 13281 39913 13367 39969
rect 13423 39913 13509 39969
rect 13565 39913 13651 39969
rect 13707 39913 13793 39969
rect 13849 39913 13935 39969
rect 13991 39913 14077 39969
rect 14133 39913 14219 39969
rect 14275 39913 14361 39969
rect 14417 39913 14503 39969
rect 14559 39913 14645 39969
rect 14701 39913 14787 39969
rect 14843 39913 14853 39969
rect 151 39827 14853 39913
rect 151 39771 161 39827
rect 217 39771 303 39827
rect 359 39771 445 39827
rect 501 39771 587 39827
rect 643 39771 729 39827
rect 785 39771 871 39827
rect 927 39771 1013 39827
rect 1069 39771 1155 39827
rect 1211 39771 1297 39827
rect 1353 39771 1439 39827
rect 1495 39771 1581 39827
rect 1637 39771 1723 39827
rect 1779 39771 1865 39827
rect 1921 39771 2007 39827
rect 2063 39771 2149 39827
rect 2205 39771 2291 39827
rect 2347 39771 2433 39827
rect 2489 39771 2575 39827
rect 2631 39771 2717 39827
rect 2773 39771 2859 39827
rect 2915 39771 3001 39827
rect 3057 39771 3143 39827
rect 3199 39771 3285 39827
rect 3341 39771 3427 39827
rect 3483 39771 3569 39827
rect 3625 39771 3711 39827
rect 3767 39771 3853 39827
rect 3909 39771 3995 39827
rect 4051 39771 4137 39827
rect 4193 39771 4279 39827
rect 4335 39771 4421 39827
rect 4477 39771 4563 39827
rect 4619 39771 4705 39827
rect 4761 39771 4847 39827
rect 4903 39771 4989 39827
rect 5045 39771 5131 39827
rect 5187 39771 5273 39827
rect 5329 39771 5415 39827
rect 5471 39771 5557 39827
rect 5613 39771 5699 39827
rect 5755 39771 5841 39827
rect 5897 39771 5983 39827
rect 6039 39771 6125 39827
rect 6181 39771 6267 39827
rect 6323 39771 6409 39827
rect 6465 39771 6551 39827
rect 6607 39771 6693 39827
rect 6749 39771 6835 39827
rect 6891 39771 6977 39827
rect 7033 39771 7119 39827
rect 7175 39771 7261 39827
rect 7317 39771 7403 39827
rect 7459 39771 7545 39827
rect 7601 39771 7687 39827
rect 7743 39771 7829 39827
rect 7885 39771 7971 39827
rect 8027 39771 8113 39827
rect 8169 39771 8255 39827
rect 8311 39771 8397 39827
rect 8453 39771 8539 39827
rect 8595 39771 8681 39827
rect 8737 39771 8823 39827
rect 8879 39771 8965 39827
rect 9021 39771 9107 39827
rect 9163 39771 9249 39827
rect 9305 39771 9391 39827
rect 9447 39771 9533 39827
rect 9589 39771 9675 39827
rect 9731 39771 9817 39827
rect 9873 39771 9959 39827
rect 10015 39771 10101 39827
rect 10157 39771 10243 39827
rect 10299 39771 10385 39827
rect 10441 39771 10527 39827
rect 10583 39771 10669 39827
rect 10725 39771 10811 39827
rect 10867 39771 10953 39827
rect 11009 39771 11095 39827
rect 11151 39771 11237 39827
rect 11293 39771 11379 39827
rect 11435 39771 11521 39827
rect 11577 39771 11663 39827
rect 11719 39771 11805 39827
rect 11861 39771 11947 39827
rect 12003 39771 12089 39827
rect 12145 39771 12231 39827
rect 12287 39771 12373 39827
rect 12429 39771 12515 39827
rect 12571 39771 12657 39827
rect 12713 39771 12799 39827
rect 12855 39771 12941 39827
rect 12997 39771 13083 39827
rect 13139 39771 13225 39827
rect 13281 39771 13367 39827
rect 13423 39771 13509 39827
rect 13565 39771 13651 39827
rect 13707 39771 13793 39827
rect 13849 39771 13935 39827
rect 13991 39771 14077 39827
rect 14133 39771 14219 39827
rect 14275 39771 14361 39827
rect 14417 39771 14503 39827
rect 14559 39771 14645 39827
rect 14701 39771 14787 39827
rect 14843 39771 14853 39827
rect 151 39685 14853 39771
rect 151 39629 161 39685
rect 217 39629 303 39685
rect 359 39629 445 39685
rect 501 39629 587 39685
rect 643 39629 729 39685
rect 785 39629 871 39685
rect 927 39629 1013 39685
rect 1069 39629 1155 39685
rect 1211 39629 1297 39685
rect 1353 39629 1439 39685
rect 1495 39629 1581 39685
rect 1637 39629 1723 39685
rect 1779 39629 1865 39685
rect 1921 39629 2007 39685
rect 2063 39629 2149 39685
rect 2205 39629 2291 39685
rect 2347 39629 2433 39685
rect 2489 39629 2575 39685
rect 2631 39629 2717 39685
rect 2773 39629 2859 39685
rect 2915 39629 3001 39685
rect 3057 39629 3143 39685
rect 3199 39629 3285 39685
rect 3341 39629 3427 39685
rect 3483 39629 3569 39685
rect 3625 39629 3711 39685
rect 3767 39629 3853 39685
rect 3909 39629 3995 39685
rect 4051 39629 4137 39685
rect 4193 39629 4279 39685
rect 4335 39629 4421 39685
rect 4477 39629 4563 39685
rect 4619 39629 4705 39685
rect 4761 39629 4847 39685
rect 4903 39629 4989 39685
rect 5045 39629 5131 39685
rect 5187 39629 5273 39685
rect 5329 39629 5415 39685
rect 5471 39629 5557 39685
rect 5613 39629 5699 39685
rect 5755 39629 5841 39685
rect 5897 39629 5983 39685
rect 6039 39629 6125 39685
rect 6181 39629 6267 39685
rect 6323 39629 6409 39685
rect 6465 39629 6551 39685
rect 6607 39629 6693 39685
rect 6749 39629 6835 39685
rect 6891 39629 6977 39685
rect 7033 39629 7119 39685
rect 7175 39629 7261 39685
rect 7317 39629 7403 39685
rect 7459 39629 7545 39685
rect 7601 39629 7687 39685
rect 7743 39629 7829 39685
rect 7885 39629 7971 39685
rect 8027 39629 8113 39685
rect 8169 39629 8255 39685
rect 8311 39629 8397 39685
rect 8453 39629 8539 39685
rect 8595 39629 8681 39685
rect 8737 39629 8823 39685
rect 8879 39629 8965 39685
rect 9021 39629 9107 39685
rect 9163 39629 9249 39685
rect 9305 39629 9391 39685
rect 9447 39629 9533 39685
rect 9589 39629 9675 39685
rect 9731 39629 9817 39685
rect 9873 39629 9959 39685
rect 10015 39629 10101 39685
rect 10157 39629 10243 39685
rect 10299 39629 10385 39685
rect 10441 39629 10527 39685
rect 10583 39629 10669 39685
rect 10725 39629 10811 39685
rect 10867 39629 10953 39685
rect 11009 39629 11095 39685
rect 11151 39629 11237 39685
rect 11293 39629 11379 39685
rect 11435 39629 11521 39685
rect 11577 39629 11663 39685
rect 11719 39629 11805 39685
rect 11861 39629 11947 39685
rect 12003 39629 12089 39685
rect 12145 39629 12231 39685
rect 12287 39629 12373 39685
rect 12429 39629 12515 39685
rect 12571 39629 12657 39685
rect 12713 39629 12799 39685
rect 12855 39629 12941 39685
rect 12997 39629 13083 39685
rect 13139 39629 13225 39685
rect 13281 39629 13367 39685
rect 13423 39629 13509 39685
rect 13565 39629 13651 39685
rect 13707 39629 13793 39685
rect 13849 39629 13935 39685
rect 13991 39629 14077 39685
rect 14133 39629 14219 39685
rect 14275 39629 14361 39685
rect 14417 39629 14503 39685
rect 14559 39629 14645 39685
rect 14701 39629 14787 39685
rect 14843 39629 14853 39685
rect 151 39619 14853 39629
rect 151 39342 14853 39352
rect 151 39286 161 39342
rect 217 39286 303 39342
rect 359 39286 445 39342
rect 501 39286 587 39342
rect 643 39286 729 39342
rect 785 39286 871 39342
rect 927 39286 1013 39342
rect 1069 39286 1155 39342
rect 1211 39286 1297 39342
rect 1353 39286 1439 39342
rect 1495 39286 1581 39342
rect 1637 39286 1723 39342
rect 1779 39286 1865 39342
rect 1921 39286 2007 39342
rect 2063 39286 2149 39342
rect 2205 39286 2291 39342
rect 2347 39286 2433 39342
rect 2489 39286 2575 39342
rect 2631 39286 2717 39342
rect 2773 39286 2859 39342
rect 2915 39286 3001 39342
rect 3057 39286 3143 39342
rect 3199 39286 3285 39342
rect 3341 39286 3427 39342
rect 3483 39286 3569 39342
rect 3625 39286 3711 39342
rect 3767 39286 3853 39342
rect 3909 39286 3995 39342
rect 4051 39286 4137 39342
rect 4193 39286 4279 39342
rect 4335 39286 4421 39342
rect 4477 39286 4563 39342
rect 4619 39286 4705 39342
rect 4761 39286 4847 39342
rect 4903 39286 4989 39342
rect 5045 39286 5131 39342
rect 5187 39286 5273 39342
rect 5329 39286 5415 39342
rect 5471 39286 5557 39342
rect 5613 39286 5699 39342
rect 5755 39286 5841 39342
rect 5897 39286 5983 39342
rect 6039 39286 6125 39342
rect 6181 39286 6267 39342
rect 6323 39286 6409 39342
rect 6465 39286 6551 39342
rect 6607 39286 6693 39342
rect 6749 39286 6835 39342
rect 6891 39286 6977 39342
rect 7033 39286 7119 39342
rect 7175 39286 7261 39342
rect 7317 39286 7403 39342
rect 7459 39286 7545 39342
rect 7601 39286 7687 39342
rect 7743 39286 7829 39342
rect 7885 39286 7971 39342
rect 8027 39286 8113 39342
rect 8169 39286 8255 39342
rect 8311 39286 8397 39342
rect 8453 39286 8539 39342
rect 8595 39286 8681 39342
rect 8737 39286 8823 39342
rect 8879 39286 8965 39342
rect 9021 39286 9107 39342
rect 9163 39286 9249 39342
rect 9305 39286 9391 39342
rect 9447 39286 9533 39342
rect 9589 39286 9675 39342
rect 9731 39286 9817 39342
rect 9873 39286 9959 39342
rect 10015 39286 10101 39342
rect 10157 39286 10243 39342
rect 10299 39286 10385 39342
rect 10441 39286 10527 39342
rect 10583 39286 10669 39342
rect 10725 39286 10811 39342
rect 10867 39286 10953 39342
rect 11009 39286 11095 39342
rect 11151 39286 11237 39342
rect 11293 39286 11379 39342
rect 11435 39286 11521 39342
rect 11577 39286 11663 39342
rect 11719 39286 11805 39342
rect 11861 39286 11947 39342
rect 12003 39286 12089 39342
rect 12145 39286 12231 39342
rect 12287 39286 12373 39342
rect 12429 39286 12515 39342
rect 12571 39286 12657 39342
rect 12713 39286 12799 39342
rect 12855 39286 12941 39342
rect 12997 39286 13083 39342
rect 13139 39286 13225 39342
rect 13281 39286 13367 39342
rect 13423 39286 13509 39342
rect 13565 39286 13651 39342
rect 13707 39286 13793 39342
rect 13849 39286 13935 39342
rect 13991 39286 14077 39342
rect 14133 39286 14219 39342
rect 14275 39286 14361 39342
rect 14417 39286 14503 39342
rect 14559 39286 14645 39342
rect 14701 39286 14787 39342
rect 14843 39286 14853 39342
rect 151 39200 14853 39286
rect 151 39144 161 39200
rect 217 39144 303 39200
rect 359 39144 445 39200
rect 501 39144 587 39200
rect 643 39144 729 39200
rect 785 39144 871 39200
rect 927 39144 1013 39200
rect 1069 39144 1155 39200
rect 1211 39144 1297 39200
rect 1353 39144 1439 39200
rect 1495 39144 1581 39200
rect 1637 39144 1723 39200
rect 1779 39144 1865 39200
rect 1921 39144 2007 39200
rect 2063 39144 2149 39200
rect 2205 39144 2291 39200
rect 2347 39144 2433 39200
rect 2489 39144 2575 39200
rect 2631 39144 2717 39200
rect 2773 39144 2859 39200
rect 2915 39144 3001 39200
rect 3057 39144 3143 39200
rect 3199 39144 3285 39200
rect 3341 39144 3427 39200
rect 3483 39144 3569 39200
rect 3625 39144 3711 39200
rect 3767 39144 3853 39200
rect 3909 39144 3995 39200
rect 4051 39144 4137 39200
rect 4193 39144 4279 39200
rect 4335 39144 4421 39200
rect 4477 39144 4563 39200
rect 4619 39144 4705 39200
rect 4761 39144 4847 39200
rect 4903 39144 4989 39200
rect 5045 39144 5131 39200
rect 5187 39144 5273 39200
rect 5329 39144 5415 39200
rect 5471 39144 5557 39200
rect 5613 39144 5699 39200
rect 5755 39144 5841 39200
rect 5897 39144 5983 39200
rect 6039 39144 6125 39200
rect 6181 39144 6267 39200
rect 6323 39144 6409 39200
rect 6465 39144 6551 39200
rect 6607 39144 6693 39200
rect 6749 39144 6835 39200
rect 6891 39144 6977 39200
rect 7033 39144 7119 39200
rect 7175 39144 7261 39200
rect 7317 39144 7403 39200
rect 7459 39144 7545 39200
rect 7601 39144 7687 39200
rect 7743 39144 7829 39200
rect 7885 39144 7971 39200
rect 8027 39144 8113 39200
rect 8169 39144 8255 39200
rect 8311 39144 8397 39200
rect 8453 39144 8539 39200
rect 8595 39144 8681 39200
rect 8737 39144 8823 39200
rect 8879 39144 8965 39200
rect 9021 39144 9107 39200
rect 9163 39144 9249 39200
rect 9305 39144 9391 39200
rect 9447 39144 9533 39200
rect 9589 39144 9675 39200
rect 9731 39144 9817 39200
rect 9873 39144 9959 39200
rect 10015 39144 10101 39200
rect 10157 39144 10243 39200
rect 10299 39144 10385 39200
rect 10441 39144 10527 39200
rect 10583 39144 10669 39200
rect 10725 39144 10811 39200
rect 10867 39144 10953 39200
rect 11009 39144 11095 39200
rect 11151 39144 11237 39200
rect 11293 39144 11379 39200
rect 11435 39144 11521 39200
rect 11577 39144 11663 39200
rect 11719 39144 11805 39200
rect 11861 39144 11947 39200
rect 12003 39144 12089 39200
rect 12145 39144 12231 39200
rect 12287 39144 12373 39200
rect 12429 39144 12515 39200
rect 12571 39144 12657 39200
rect 12713 39144 12799 39200
rect 12855 39144 12941 39200
rect 12997 39144 13083 39200
rect 13139 39144 13225 39200
rect 13281 39144 13367 39200
rect 13423 39144 13509 39200
rect 13565 39144 13651 39200
rect 13707 39144 13793 39200
rect 13849 39144 13935 39200
rect 13991 39144 14077 39200
rect 14133 39144 14219 39200
rect 14275 39144 14361 39200
rect 14417 39144 14503 39200
rect 14559 39144 14645 39200
rect 14701 39144 14787 39200
rect 14843 39144 14853 39200
rect 151 39058 14853 39144
rect 151 39002 161 39058
rect 217 39002 303 39058
rect 359 39002 445 39058
rect 501 39002 587 39058
rect 643 39002 729 39058
rect 785 39002 871 39058
rect 927 39002 1013 39058
rect 1069 39002 1155 39058
rect 1211 39002 1297 39058
rect 1353 39002 1439 39058
rect 1495 39002 1581 39058
rect 1637 39002 1723 39058
rect 1779 39002 1865 39058
rect 1921 39002 2007 39058
rect 2063 39002 2149 39058
rect 2205 39002 2291 39058
rect 2347 39002 2433 39058
rect 2489 39002 2575 39058
rect 2631 39002 2717 39058
rect 2773 39002 2859 39058
rect 2915 39002 3001 39058
rect 3057 39002 3143 39058
rect 3199 39002 3285 39058
rect 3341 39002 3427 39058
rect 3483 39002 3569 39058
rect 3625 39002 3711 39058
rect 3767 39002 3853 39058
rect 3909 39002 3995 39058
rect 4051 39002 4137 39058
rect 4193 39002 4279 39058
rect 4335 39002 4421 39058
rect 4477 39002 4563 39058
rect 4619 39002 4705 39058
rect 4761 39002 4847 39058
rect 4903 39002 4989 39058
rect 5045 39002 5131 39058
rect 5187 39002 5273 39058
rect 5329 39002 5415 39058
rect 5471 39002 5557 39058
rect 5613 39002 5699 39058
rect 5755 39002 5841 39058
rect 5897 39002 5983 39058
rect 6039 39002 6125 39058
rect 6181 39002 6267 39058
rect 6323 39002 6409 39058
rect 6465 39002 6551 39058
rect 6607 39002 6693 39058
rect 6749 39002 6835 39058
rect 6891 39002 6977 39058
rect 7033 39002 7119 39058
rect 7175 39002 7261 39058
rect 7317 39002 7403 39058
rect 7459 39002 7545 39058
rect 7601 39002 7687 39058
rect 7743 39002 7829 39058
rect 7885 39002 7971 39058
rect 8027 39002 8113 39058
rect 8169 39002 8255 39058
rect 8311 39002 8397 39058
rect 8453 39002 8539 39058
rect 8595 39002 8681 39058
rect 8737 39002 8823 39058
rect 8879 39002 8965 39058
rect 9021 39002 9107 39058
rect 9163 39002 9249 39058
rect 9305 39002 9391 39058
rect 9447 39002 9533 39058
rect 9589 39002 9675 39058
rect 9731 39002 9817 39058
rect 9873 39002 9959 39058
rect 10015 39002 10101 39058
rect 10157 39002 10243 39058
rect 10299 39002 10385 39058
rect 10441 39002 10527 39058
rect 10583 39002 10669 39058
rect 10725 39002 10811 39058
rect 10867 39002 10953 39058
rect 11009 39002 11095 39058
rect 11151 39002 11237 39058
rect 11293 39002 11379 39058
rect 11435 39002 11521 39058
rect 11577 39002 11663 39058
rect 11719 39002 11805 39058
rect 11861 39002 11947 39058
rect 12003 39002 12089 39058
rect 12145 39002 12231 39058
rect 12287 39002 12373 39058
rect 12429 39002 12515 39058
rect 12571 39002 12657 39058
rect 12713 39002 12799 39058
rect 12855 39002 12941 39058
rect 12997 39002 13083 39058
rect 13139 39002 13225 39058
rect 13281 39002 13367 39058
rect 13423 39002 13509 39058
rect 13565 39002 13651 39058
rect 13707 39002 13793 39058
rect 13849 39002 13935 39058
rect 13991 39002 14077 39058
rect 14133 39002 14219 39058
rect 14275 39002 14361 39058
rect 14417 39002 14503 39058
rect 14559 39002 14645 39058
rect 14701 39002 14787 39058
rect 14843 39002 14853 39058
rect 151 38916 14853 39002
rect 151 38860 161 38916
rect 217 38860 303 38916
rect 359 38860 445 38916
rect 501 38860 587 38916
rect 643 38860 729 38916
rect 785 38860 871 38916
rect 927 38860 1013 38916
rect 1069 38860 1155 38916
rect 1211 38860 1297 38916
rect 1353 38860 1439 38916
rect 1495 38860 1581 38916
rect 1637 38860 1723 38916
rect 1779 38860 1865 38916
rect 1921 38860 2007 38916
rect 2063 38860 2149 38916
rect 2205 38860 2291 38916
rect 2347 38860 2433 38916
rect 2489 38860 2575 38916
rect 2631 38860 2717 38916
rect 2773 38860 2859 38916
rect 2915 38860 3001 38916
rect 3057 38860 3143 38916
rect 3199 38860 3285 38916
rect 3341 38860 3427 38916
rect 3483 38860 3569 38916
rect 3625 38860 3711 38916
rect 3767 38860 3853 38916
rect 3909 38860 3995 38916
rect 4051 38860 4137 38916
rect 4193 38860 4279 38916
rect 4335 38860 4421 38916
rect 4477 38860 4563 38916
rect 4619 38860 4705 38916
rect 4761 38860 4847 38916
rect 4903 38860 4989 38916
rect 5045 38860 5131 38916
rect 5187 38860 5273 38916
rect 5329 38860 5415 38916
rect 5471 38860 5557 38916
rect 5613 38860 5699 38916
rect 5755 38860 5841 38916
rect 5897 38860 5983 38916
rect 6039 38860 6125 38916
rect 6181 38860 6267 38916
rect 6323 38860 6409 38916
rect 6465 38860 6551 38916
rect 6607 38860 6693 38916
rect 6749 38860 6835 38916
rect 6891 38860 6977 38916
rect 7033 38860 7119 38916
rect 7175 38860 7261 38916
rect 7317 38860 7403 38916
rect 7459 38860 7545 38916
rect 7601 38860 7687 38916
rect 7743 38860 7829 38916
rect 7885 38860 7971 38916
rect 8027 38860 8113 38916
rect 8169 38860 8255 38916
rect 8311 38860 8397 38916
rect 8453 38860 8539 38916
rect 8595 38860 8681 38916
rect 8737 38860 8823 38916
rect 8879 38860 8965 38916
rect 9021 38860 9107 38916
rect 9163 38860 9249 38916
rect 9305 38860 9391 38916
rect 9447 38860 9533 38916
rect 9589 38860 9675 38916
rect 9731 38860 9817 38916
rect 9873 38860 9959 38916
rect 10015 38860 10101 38916
rect 10157 38860 10243 38916
rect 10299 38860 10385 38916
rect 10441 38860 10527 38916
rect 10583 38860 10669 38916
rect 10725 38860 10811 38916
rect 10867 38860 10953 38916
rect 11009 38860 11095 38916
rect 11151 38860 11237 38916
rect 11293 38860 11379 38916
rect 11435 38860 11521 38916
rect 11577 38860 11663 38916
rect 11719 38860 11805 38916
rect 11861 38860 11947 38916
rect 12003 38860 12089 38916
rect 12145 38860 12231 38916
rect 12287 38860 12373 38916
rect 12429 38860 12515 38916
rect 12571 38860 12657 38916
rect 12713 38860 12799 38916
rect 12855 38860 12941 38916
rect 12997 38860 13083 38916
rect 13139 38860 13225 38916
rect 13281 38860 13367 38916
rect 13423 38860 13509 38916
rect 13565 38860 13651 38916
rect 13707 38860 13793 38916
rect 13849 38860 13935 38916
rect 13991 38860 14077 38916
rect 14133 38860 14219 38916
rect 14275 38860 14361 38916
rect 14417 38860 14503 38916
rect 14559 38860 14645 38916
rect 14701 38860 14787 38916
rect 14843 38860 14853 38916
rect 151 38774 14853 38860
rect 151 38718 161 38774
rect 217 38718 303 38774
rect 359 38718 445 38774
rect 501 38718 587 38774
rect 643 38718 729 38774
rect 785 38718 871 38774
rect 927 38718 1013 38774
rect 1069 38718 1155 38774
rect 1211 38718 1297 38774
rect 1353 38718 1439 38774
rect 1495 38718 1581 38774
rect 1637 38718 1723 38774
rect 1779 38718 1865 38774
rect 1921 38718 2007 38774
rect 2063 38718 2149 38774
rect 2205 38718 2291 38774
rect 2347 38718 2433 38774
rect 2489 38718 2575 38774
rect 2631 38718 2717 38774
rect 2773 38718 2859 38774
rect 2915 38718 3001 38774
rect 3057 38718 3143 38774
rect 3199 38718 3285 38774
rect 3341 38718 3427 38774
rect 3483 38718 3569 38774
rect 3625 38718 3711 38774
rect 3767 38718 3853 38774
rect 3909 38718 3995 38774
rect 4051 38718 4137 38774
rect 4193 38718 4279 38774
rect 4335 38718 4421 38774
rect 4477 38718 4563 38774
rect 4619 38718 4705 38774
rect 4761 38718 4847 38774
rect 4903 38718 4989 38774
rect 5045 38718 5131 38774
rect 5187 38718 5273 38774
rect 5329 38718 5415 38774
rect 5471 38718 5557 38774
rect 5613 38718 5699 38774
rect 5755 38718 5841 38774
rect 5897 38718 5983 38774
rect 6039 38718 6125 38774
rect 6181 38718 6267 38774
rect 6323 38718 6409 38774
rect 6465 38718 6551 38774
rect 6607 38718 6693 38774
rect 6749 38718 6835 38774
rect 6891 38718 6977 38774
rect 7033 38718 7119 38774
rect 7175 38718 7261 38774
rect 7317 38718 7403 38774
rect 7459 38718 7545 38774
rect 7601 38718 7687 38774
rect 7743 38718 7829 38774
rect 7885 38718 7971 38774
rect 8027 38718 8113 38774
rect 8169 38718 8255 38774
rect 8311 38718 8397 38774
rect 8453 38718 8539 38774
rect 8595 38718 8681 38774
rect 8737 38718 8823 38774
rect 8879 38718 8965 38774
rect 9021 38718 9107 38774
rect 9163 38718 9249 38774
rect 9305 38718 9391 38774
rect 9447 38718 9533 38774
rect 9589 38718 9675 38774
rect 9731 38718 9817 38774
rect 9873 38718 9959 38774
rect 10015 38718 10101 38774
rect 10157 38718 10243 38774
rect 10299 38718 10385 38774
rect 10441 38718 10527 38774
rect 10583 38718 10669 38774
rect 10725 38718 10811 38774
rect 10867 38718 10953 38774
rect 11009 38718 11095 38774
rect 11151 38718 11237 38774
rect 11293 38718 11379 38774
rect 11435 38718 11521 38774
rect 11577 38718 11663 38774
rect 11719 38718 11805 38774
rect 11861 38718 11947 38774
rect 12003 38718 12089 38774
rect 12145 38718 12231 38774
rect 12287 38718 12373 38774
rect 12429 38718 12515 38774
rect 12571 38718 12657 38774
rect 12713 38718 12799 38774
rect 12855 38718 12941 38774
rect 12997 38718 13083 38774
rect 13139 38718 13225 38774
rect 13281 38718 13367 38774
rect 13423 38718 13509 38774
rect 13565 38718 13651 38774
rect 13707 38718 13793 38774
rect 13849 38718 13935 38774
rect 13991 38718 14077 38774
rect 14133 38718 14219 38774
rect 14275 38718 14361 38774
rect 14417 38718 14503 38774
rect 14559 38718 14645 38774
rect 14701 38718 14787 38774
rect 14843 38718 14853 38774
rect 151 38632 14853 38718
rect 151 38576 161 38632
rect 217 38576 303 38632
rect 359 38576 445 38632
rect 501 38576 587 38632
rect 643 38576 729 38632
rect 785 38576 871 38632
rect 927 38576 1013 38632
rect 1069 38576 1155 38632
rect 1211 38576 1297 38632
rect 1353 38576 1439 38632
rect 1495 38576 1581 38632
rect 1637 38576 1723 38632
rect 1779 38576 1865 38632
rect 1921 38576 2007 38632
rect 2063 38576 2149 38632
rect 2205 38576 2291 38632
rect 2347 38576 2433 38632
rect 2489 38576 2575 38632
rect 2631 38576 2717 38632
rect 2773 38576 2859 38632
rect 2915 38576 3001 38632
rect 3057 38576 3143 38632
rect 3199 38576 3285 38632
rect 3341 38576 3427 38632
rect 3483 38576 3569 38632
rect 3625 38576 3711 38632
rect 3767 38576 3853 38632
rect 3909 38576 3995 38632
rect 4051 38576 4137 38632
rect 4193 38576 4279 38632
rect 4335 38576 4421 38632
rect 4477 38576 4563 38632
rect 4619 38576 4705 38632
rect 4761 38576 4847 38632
rect 4903 38576 4989 38632
rect 5045 38576 5131 38632
rect 5187 38576 5273 38632
rect 5329 38576 5415 38632
rect 5471 38576 5557 38632
rect 5613 38576 5699 38632
rect 5755 38576 5841 38632
rect 5897 38576 5983 38632
rect 6039 38576 6125 38632
rect 6181 38576 6267 38632
rect 6323 38576 6409 38632
rect 6465 38576 6551 38632
rect 6607 38576 6693 38632
rect 6749 38576 6835 38632
rect 6891 38576 6977 38632
rect 7033 38576 7119 38632
rect 7175 38576 7261 38632
rect 7317 38576 7403 38632
rect 7459 38576 7545 38632
rect 7601 38576 7687 38632
rect 7743 38576 7829 38632
rect 7885 38576 7971 38632
rect 8027 38576 8113 38632
rect 8169 38576 8255 38632
rect 8311 38576 8397 38632
rect 8453 38576 8539 38632
rect 8595 38576 8681 38632
rect 8737 38576 8823 38632
rect 8879 38576 8965 38632
rect 9021 38576 9107 38632
rect 9163 38576 9249 38632
rect 9305 38576 9391 38632
rect 9447 38576 9533 38632
rect 9589 38576 9675 38632
rect 9731 38576 9817 38632
rect 9873 38576 9959 38632
rect 10015 38576 10101 38632
rect 10157 38576 10243 38632
rect 10299 38576 10385 38632
rect 10441 38576 10527 38632
rect 10583 38576 10669 38632
rect 10725 38576 10811 38632
rect 10867 38576 10953 38632
rect 11009 38576 11095 38632
rect 11151 38576 11237 38632
rect 11293 38576 11379 38632
rect 11435 38576 11521 38632
rect 11577 38576 11663 38632
rect 11719 38576 11805 38632
rect 11861 38576 11947 38632
rect 12003 38576 12089 38632
rect 12145 38576 12231 38632
rect 12287 38576 12373 38632
rect 12429 38576 12515 38632
rect 12571 38576 12657 38632
rect 12713 38576 12799 38632
rect 12855 38576 12941 38632
rect 12997 38576 13083 38632
rect 13139 38576 13225 38632
rect 13281 38576 13367 38632
rect 13423 38576 13509 38632
rect 13565 38576 13651 38632
rect 13707 38576 13793 38632
rect 13849 38576 13935 38632
rect 13991 38576 14077 38632
rect 14133 38576 14219 38632
rect 14275 38576 14361 38632
rect 14417 38576 14503 38632
rect 14559 38576 14645 38632
rect 14701 38576 14787 38632
rect 14843 38576 14853 38632
rect 151 38490 14853 38576
rect 151 38434 161 38490
rect 217 38434 303 38490
rect 359 38434 445 38490
rect 501 38434 587 38490
rect 643 38434 729 38490
rect 785 38434 871 38490
rect 927 38434 1013 38490
rect 1069 38434 1155 38490
rect 1211 38434 1297 38490
rect 1353 38434 1439 38490
rect 1495 38434 1581 38490
rect 1637 38434 1723 38490
rect 1779 38434 1865 38490
rect 1921 38434 2007 38490
rect 2063 38434 2149 38490
rect 2205 38434 2291 38490
rect 2347 38434 2433 38490
rect 2489 38434 2575 38490
rect 2631 38434 2717 38490
rect 2773 38434 2859 38490
rect 2915 38434 3001 38490
rect 3057 38434 3143 38490
rect 3199 38434 3285 38490
rect 3341 38434 3427 38490
rect 3483 38434 3569 38490
rect 3625 38434 3711 38490
rect 3767 38434 3853 38490
rect 3909 38434 3995 38490
rect 4051 38434 4137 38490
rect 4193 38434 4279 38490
rect 4335 38434 4421 38490
rect 4477 38434 4563 38490
rect 4619 38434 4705 38490
rect 4761 38434 4847 38490
rect 4903 38434 4989 38490
rect 5045 38434 5131 38490
rect 5187 38434 5273 38490
rect 5329 38434 5415 38490
rect 5471 38434 5557 38490
rect 5613 38434 5699 38490
rect 5755 38434 5841 38490
rect 5897 38434 5983 38490
rect 6039 38434 6125 38490
rect 6181 38434 6267 38490
rect 6323 38434 6409 38490
rect 6465 38434 6551 38490
rect 6607 38434 6693 38490
rect 6749 38434 6835 38490
rect 6891 38434 6977 38490
rect 7033 38434 7119 38490
rect 7175 38434 7261 38490
rect 7317 38434 7403 38490
rect 7459 38434 7545 38490
rect 7601 38434 7687 38490
rect 7743 38434 7829 38490
rect 7885 38434 7971 38490
rect 8027 38434 8113 38490
rect 8169 38434 8255 38490
rect 8311 38434 8397 38490
rect 8453 38434 8539 38490
rect 8595 38434 8681 38490
rect 8737 38434 8823 38490
rect 8879 38434 8965 38490
rect 9021 38434 9107 38490
rect 9163 38434 9249 38490
rect 9305 38434 9391 38490
rect 9447 38434 9533 38490
rect 9589 38434 9675 38490
rect 9731 38434 9817 38490
rect 9873 38434 9959 38490
rect 10015 38434 10101 38490
rect 10157 38434 10243 38490
rect 10299 38434 10385 38490
rect 10441 38434 10527 38490
rect 10583 38434 10669 38490
rect 10725 38434 10811 38490
rect 10867 38434 10953 38490
rect 11009 38434 11095 38490
rect 11151 38434 11237 38490
rect 11293 38434 11379 38490
rect 11435 38434 11521 38490
rect 11577 38434 11663 38490
rect 11719 38434 11805 38490
rect 11861 38434 11947 38490
rect 12003 38434 12089 38490
rect 12145 38434 12231 38490
rect 12287 38434 12373 38490
rect 12429 38434 12515 38490
rect 12571 38434 12657 38490
rect 12713 38434 12799 38490
rect 12855 38434 12941 38490
rect 12997 38434 13083 38490
rect 13139 38434 13225 38490
rect 13281 38434 13367 38490
rect 13423 38434 13509 38490
rect 13565 38434 13651 38490
rect 13707 38434 13793 38490
rect 13849 38434 13935 38490
rect 13991 38434 14077 38490
rect 14133 38434 14219 38490
rect 14275 38434 14361 38490
rect 14417 38434 14503 38490
rect 14559 38434 14645 38490
rect 14701 38434 14787 38490
rect 14843 38434 14853 38490
rect 151 38348 14853 38434
rect 151 38292 161 38348
rect 217 38292 303 38348
rect 359 38292 445 38348
rect 501 38292 587 38348
rect 643 38292 729 38348
rect 785 38292 871 38348
rect 927 38292 1013 38348
rect 1069 38292 1155 38348
rect 1211 38292 1297 38348
rect 1353 38292 1439 38348
rect 1495 38292 1581 38348
rect 1637 38292 1723 38348
rect 1779 38292 1865 38348
rect 1921 38292 2007 38348
rect 2063 38292 2149 38348
rect 2205 38292 2291 38348
rect 2347 38292 2433 38348
rect 2489 38292 2575 38348
rect 2631 38292 2717 38348
rect 2773 38292 2859 38348
rect 2915 38292 3001 38348
rect 3057 38292 3143 38348
rect 3199 38292 3285 38348
rect 3341 38292 3427 38348
rect 3483 38292 3569 38348
rect 3625 38292 3711 38348
rect 3767 38292 3853 38348
rect 3909 38292 3995 38348
rect 4051 38292 4137 38348
rect 4193 38292 4279 38348
rect 4335 38292 4421 38348
rect 4477 38292 4563 38348
rect 4619 38292 4705 38348
rect 4761 38292 4847 38348
rect 4903 38292 4989 38348
rect 5045 38292 5131 38348
rect 5187 38292 5273 38348
rect 5329 38292 5415 38348
rect 5471 38292 5557 38348
rect 5613 38292 5699 38348
rect 5755 38292 5841 38348
rect 5897 38292 5983 38348
rect 6039 38292 6125 38348
rect 6181 38292 6267 38348
rect 6323 38292 6409 38348
rect 6465 38292 6551 38348
rect 6607 38292 6693 38348
rect 6749 38292 6835 38348
rect 6891 38292 6977 38348
rect 7033 38292 7119 38348
rect 7175 38292 7261 38348
rect 7317 38292 7403 38348
rect 7459 38292 7545 38348
rect 7601 38292 7687 38348
rect 7743 38292 7829 38348
rect 7885 38292 7971 38348
rect 8027 38292 8113 38348
rect 8169 38292 8255 38348
rect 8311 38292 8397 38348
rect 8453 38292 8539 38348
rect 8595 38292 8681 38348
rect 8737 38292 8823 38348
rect 8879 38292 8965 38348
rect 9021 38292 9107 38348
rect 9163 38292 9249 38348
rect 9305 38292 9391 38348
rect 9447 38292 9533 38348
rect 9589 38292 9675 38348
rect 9731 38292 9817 38348
rect 9873 38292 9959 38348
rect 10015 38292 10101 38348
rect 10157 38292 10243 38348
rect 10299 38292 10385 38348
rect 10441 38292 10527 38348
rect 10583 38292 10669 38348
rect 10725 38292 10811 38348
rect 10867 38292 10953 38348
rect 11009 38292 11095 38348
rect 11151 38292 11237 38348
rect 11293 38292 11379 38348
rect 11435 38292 11521 38348
rect 11577 38292 11663 38348
rect 11719 38292 11805 38348
rect 11861 38292 11947 38348
rect 12003 38292 12089 38348
rect 12145 38292 12231 38348
rect 12287 38292 12373 38348
rect 12429 38292 12515 38348
rect 12571 38292 12657 38348
rect 12713 38292 12799 38348
rect 12855 38292 12941 38348
rect 12997 38292 13083 38348
rect 13139 38292 13225 38348
rect 13281 38292 13367 38348
rect 13423 38292 13509 38348
rect 13565 38292 13651 38348
rect 13707 38292 13793 38348
rect 13849 38292 13935 38348
rect 13991 38292 14077 38348
rect 14133 38292 14219 38348
rect 14275 38292 14361 38348
rect 14417 38292 14503 38348
rect 14559 38292 14645 38348
rect 14701 38292 14787 38348
rect 14843 38292 14853 38348
rect 151 38206 14853 38292
rect 151 38150 161 38206
rect 217 38150 303 38206
rect 359 38150 445 38206
rect 501 38150 587 38206
rect 643 38150 729 38206
rect 785 38150 871 38206
rect 927 38150 1013 38206
rect 1069 38150 1155 38206
rect 1211 38150 1297 38206
rect 1353 38150 1439 38206
rect 1495 38150 1581 38206
rect 1637 38150 1723 38206
rect 1779 38150 1865 38206
rect 1921 38150 2007 38206
rect 2063 38150 2149 38206
rect 2205 38150 2291 38206
rect 2347 38150 2433 38206
rect 2489 38150 2575 38206
rect 2631 38150 2717 38206
rect 2773 38150 2859 38206
rect 2915 38150 3001 38206
rect 3057 38150 3143 38206
rect 3199 38150 3285 38206
rect 3341 38150 3427 38206
rect 3483 38150 3569 38206
rect 3625 38150 3711 38206
rect 3767 38150 3853 38206
rect 3909 38150 3995 38206
rect 4051 38150 4137 38206
rect 4193 38150 4279 38206
rect 4335 38150 4421 38206
rect 4477 38150 4563 38206
rect 4619 38150 4705 38206
rect 4761 38150 4847 38206
rect 4903 38150 4989 38206
rect 5045 38150 5131 38206
rect 5187 38150 5273 38206
rect 5329 38150 5415 38206
rect 5471 38150 5557 38206
rect 5613 38150 5699 38206
rect 5755 38150 5841 38206
rect 5897 38150 5983 38206
rect 6039 38150 6125 38206
rect 6181 38150 6267 38206
rect 6323 38150 6409 38206
rect 6465 38150 6551 38206
rect 6607 38150 6693 38206
rect 6749 38150 6835 38206
rect 6891 38150 6977 38206
rect 7033 38150 7119 38206
rect 7175 38150 7261 38206
rect 7317 38150 7403 38206
rect 7459 38150 7545 38206
rect 7601 38150 7687 38206
rect 7743 38150 7829 38206
rect 7885 38150 7971 38206
rect 8027 38150 8113 38206
rect 8169 38150 8255 38206
rect 8311 38150 8397 38206
rect 8453 38150 8539 38206
rect 8595 38150 8681 38206
rect 8737 38150 8823 38206
rect 8879 38150 8965 38206
rect 9021 38150 9107 38206
rect 9163 38150 9249 38206
rect 9305 38150 9391 38206
rect 9447 38150 9533 38206
rect 9589 38150 9675 38206
rect 9731 38150 9817 38206
rect 9873 38150 9959 38206
rect 10015 38150 10101 38206
rect 10157 38150 10243 38206
rect 10299 38150 10385 38206
rect 10441 38150 10527 38206
rect 10583 38150 10669 38206
rect 10725 38150 10811 38206
rect 10867 38150 10953 38206
rect 11009 38150 11095 38206
rect 11151 38150 11237 38206
rect 11293 38150 11379 38206
rect 11435 38150 11521 38206
rect 11577 38150 11663 38206
rect 11719 38150 11805 38206
rect 11861 38150 11947 38206
rect 12003 38150 12089 38206
rect 12145 38150 12231 38206
rect 12287 38150 12373 38206
rect 12429 38150 12515 38206
rect 12571 38150 12657 38206
rect 12713 38150 12799 38206
rect 12855 38150 12941 38206
rect 12997 38150 13083 38206
rect 13139 38150 13225 38206
rect 13281 38150 13367 38206
rect 13423 38150 13509 38206
rect 13565 38150 13651 38206
rect 13707 38150 13793 38206
rect 13849 38150 13935 38206
rect 13991 38150 14077 38206
rect 14133 38150 14219 38206
rect 14275 38150 14361 38206
rect 14417 38150 14503 38206
rect 14559 38150 14645 38206
rect 14701 38150 14787 38206
rect 14843 38150 14853 38206
rect 151 38064 14853 38150
rect 151 38008 161 38064
rect 217 38008 303 38064
rect 359 38008 445 38064
rect 501 38008 587 38064
rect 643 38008 729 38064
rect 785 38008 871 38064
rect 927 38008 1013 38064
rect 1069 38008 1155 38064
rect 1211 38008 1297 38064
rect 1353 38008 1439 38064
rect 1495 38008 1581 38064
rect 1637 38008 1723 38064
rect 1779 38008 1865 38064
rect 1921 38008 2007 38064
rect 2063 38008 2149 38064
rect 2205 38008 2291 38064
rect 2347 38008 2433 38064
rect 2489 38008 2575 38064
rect 2631 38008 2717 38064
rect 2773 38008 2859 38064
rect 2915 38008 3001 38064
rect 3057 38008 3143 38064
rect 3199 38008 3285 38064
rect 3341 38008 3427 38064
rect 3483 38008 3569 38064
rect 3625 38008 3711 38064
rect 3767 38008 3853 38064
rect 3909 38008 3995 38064
rect 4051 38008 4137 38064
rect 4193 38008 4279 38064
rect 4335 38008 4421 38064
rect 4477 38008 4563 38064
rect 4619 38008 4705 38064
rect 4761 38008 4847 38064
rect 4903 38008 4989 38064
rect 5045 38008 5131 38064
rect 5187 38008 5273 38064
rect 5329 38008 5415 38064
rect 5471 38008 5557 38064
rect 5613 38008 5699 38064
rect 5755 38008 5841 38064
rect 5897 38008 5983 38064
rect 6039 38008 6125 38064
rect 6181 38008 6267 38064
rect 6323 38008 6409 38064
rect 6465 38008 6551 38064
rect 6607 38008 6693 38064
rect 6749 38008 6835 38064
rect 6891 38008 6977 38064
rect 7033 38008 7119 38064
rect 7175 38008 7261 38064
rect 7317 38008 7403 38064
rect 7459 38008 7545 38064
rect 7601 38008 7687 38064
rect 7743 38008 7829 38064
rect 7885 38008 7971 38064
rect 8027 38008 8113 38064
rect 8169 38008 8255 38064
rect 8311 38008 8397 38064
rect 8453 38008 8539 38064
rect 8595 38008 8681 38064
rect 8737 38008 8823 38064
rect 8879 38008 8965 38064
rect 9021 38008 9107 38064
rect 9163 38008 9249 38064
rect 9305 38008 9391 38064
rect 9447 38008 9533 38064
rect 9589 38008 9675 38064
rect 9731 38008 9817 38064
rect 9873 38008 9959 38064
rect 10015 38008 10101 38064
rect 10157 38008 10243 38064
rect 10299 38008 10385 38064
rect 10441 38008 10527 38064
rect 10583 38008 10669 38064
rect 10725 38008 10811 38064
rect 10867 38008 10953 38064
rect 11009 38008 11095 38064
rect 11151 38008 11237 38064
rect 11293 38008 11379 38064
rect 11435 38008 11521 38064
rect 11577 38008 11663 38064
rect 11719 38008 11805 38064
rect 11861 38008 11947 38064
rect 12003 38008 12089 38064
rect 12145 38008 12231 38064
rect 12287 38008 12373 38064
rect 12429 38008 12515 38064
rect 12571 38008 12657 38064
rect 12713 38008 12799 38064
rect 12855 38008 12941 38064
rect 12997 38008 13083 38064
rect 13139 38008 13225 38064
rect 13281 38008 13367 38064
rect 13423 38008 13509 38064
rect 13565 38008 13651 38064
rect 13707 38008 13793 38064
rect 13849 38008 13935 38064
rect 13991 38008 14077 38064
rect 14133 38008 14219 38064
rect 14275 38008 14361 38064
rect 14417 38008 14503 38064
rect 14559 38008 14645 38064
rect 14701 38008 14787 38064
rect 14843 38008 14853 38064
rect 151 37922 14853 38008
rect 151 37866 161 37922
rect 217 37866 303 37922
rect 359 37866 445 37922
rect 501 37866 587 37922
rect 643 37866 729 37922
rect 785 37866 871 37922
rect 927 37866 1013 37922
rect 1069 37866 1155 37922
rect 1211 37866 1297 37922
rect 1353 37866 1439 37922
rect 1495 37866 1581 37922
rect 1637 37866 1723 37922
rect 1779 37866 1865 37922
rect 1921 37866 2007 37922
rect 2063 37866 2149 37922
rect 2205 37866 2291 37922
rect 2347 37866 2433 37922
rect 2489 37866 2575 37922
rect 2631 37866 2717 37922
rect 2773 37866 2859 37922
rect 2915 37866 3001 37922
rect 3057 37866 3143 37922
rect 3199 37866 3285 37922
rect 3341 37866 3427 37922
rect 3483 37866 3569 37922
rect 3625 37866 3711 37922
rect 3767 37866 3853 37922
rect 3909 37866 3995 37922
rect 4051 37866 4137 37922
rect 4193 37866 4279 37922
rect 4335 37866 4421 37922
rect 4477 37866 4563 37922
rect 4619 37866 4705 37922
rect 4761 37866 4847 37922
rect 4903 37866 4989 37922
rect 5045 37866 5131 37922
rect 5187 37866 5273 37922
rect 5329 37866 5415 37922
rect 5471 37866 5557 37922
rect 5613 37866 5699 37922
rect 5755 37866 5841 37922
rect 5897 37866 5983 37922
rect 6039 37866 6125 37922
rect 6181 37866 6267 37922
rect 6323 37866 6409 37922
rect 6465 37866 6551 37922
rect 6607 37866 6693 37922
rect 6749 37866 6835 37922
rect 6891 37866 6977 37922
rect 7033 37866 7119 37922
rect 7175 37866 7261 37922
rect 7317 37866 7403 37922
rect 7459 37866 7545 37922
rect 7601 37866 7687 37922
rect 7743 37866 7829 37922
rect 7885 37866 7971 37922
rect 8027 37866 8113 37922
rect 8169 37866 8255 37922
rect 8311 37866 8397 37922
rect 8453 37866 8539 37922
rect 8595 37866 8681 37922
rect 8737 37866 8823 37922
rect 8879 37866 8965 37922
rect 9021 37866 9107 37922
rect 9163 37866 9249 37922
rect 9305 37866 9391 37922
rect 9447 37866 9533 37922
rect 9589 37866 9675 37922
rect 9731 37866 9817 37922
rect 9873 37866 9959 37922
rect 10015 37866 10101 37922
rect 10157 37866 10243 37922
rect 10299 37866 10385 37922
rect 10441 37866 10527 37922
rect 10583 37866 10669 37922
rect 10725 37866 10811 37922
rect 10867 37866 10953 37922
rect 11009 37866 11095 37922
rect 11151 37866 11237 37922
rect 11293 37866 11379 37922
rect 11435 37866 11521 37922
rect 11577 37866 11663 37922
rect 11719 37866 11805 37922
rect 11861 37866 11947 37922
rect 12003 37866 12089 37922
rect 12145 37866 12231 37922
rect 12287 37866 12373 37922
rect 12429 37866 12515 37922
rect 12571 37866 12657 37922
rect 12713 37866 12799 37922
rect 12855 37866 12941 37922
rect 12997 37866 13083 37922
rect 13139 37866 13225 37922
rect 13281 37866 13367 37922
rect 13423 37866 13509 37922
rect 13565 37866 13651 37922
rect 13707 37866 13793 37922
rect 13849 37866 13935 37922
rect 13991 37866 14077 37922
rect 14133 37866 14219 37922
rect 14275 37866 14361 37922
rect 14417 37866 14503 37922
rect 14559 37866 14645 37922
rect 14701 37866 14787 37922
rect 14843 37866 14853 37922
rect 151 37780 14853 37866
rect 151 37724 161 37780
rect 217 37724 303 37780
rect 359 37724 445 37780
rect 501 37724 587 37780
rect 643 37724 729 37780
rect 785 37724 871 37780
rect 927 37724 1013 37780
rect 1069 37724 1155 37780
rect 1211 37724 1297 37780
rect 1353 37724 1439 37780
rect 1495 37724 1581 37780
rect 1637 37724 1723 37780
rect 1779 37724 1865 37780
rect 1921 37724 2007 37780
rect 2063 37724 2149 37780
rect 2205 37724 2291 37780
rect 2347 37724 2433 37780
rect 2489 37724 2575 37780
rect 2631 37724 2717 37780
rect 2773 37724 2859 37780
rect 2915 37724 3001 37780
rect 3057 37724 3143 37780
rect 3199 37724 3285 37780
rect 3341 37724 3427 37780
rect 3483 37724 3569 37780
rect 3625 37724 3711 37780
rect 3767 37724 3853 37780
rect 3909 37724 3995 37780
rect 4051 37724 4137 37780
rect 4193 37724 4279 37780
rect 4335 37724 4421 37780
rect 4477 37724 4563 37780
rect 4619 37724 4705 37780
rect 4761 37724 4847 37780
rect 4903 37724 4989 37780
rect 5045 37724 5131 37780
rect 5187 37724 5273 37780
rect 5329 37724 5415 37780
rect 5471 37724 5557 37780
rect 5613 37724 5699 37780
rect 5755 37724 5841 37780
rect 5897 37724 5983 37780
rect 6039 37724 6125 37780
rect 6181 37724 6267 37780
rect 6323 37724 6409 37780
rect 6465 37724 6551 37780
rect 6607 37724 6693 37780
rect 6749 37724 6835 37780
rect 6891 37724 6977 37780
rect 7033 37724 7119 37780
rect 7175 37724 7261 37780
rect 7317 37724 7403 37780
rect 7459 37724 7545 37780
rect 7601 37724 7687 37780
rect 7743 37724 7829 37780
rect 7885 37724 7971 37780
rect 8027 37724 8113 37780
rect 8169 37724 8255 37780
rect 8311 37724 8397 37780
rect 8453 37724 8539 37780
rect 8595 37724 8681 37780
rect 8737 37724 8823 37780
rect 8879 37724 8965 37780
rect 9021 37724 9107 37780
rect 9163 37724 9249 37780
rect 9305 37724 9391 37780
rect 9447 37724 9533 37780
rect 9589 37724 9675 37780
rect 9731 37724 9817 37780
rect 9873 37724 9959 37780
rect 10015 37724 10101 37780
rect 10157 37724 10243 37780
rect 10299 37724 10385 37780
rect 10441 37724 10527 37780
rect 10583 37724 10669 37780
rect 10725 37724 10811 37780
rect 10867 37724 10953 37780
rect 11009 37724 11095 37780
rect 11151 37724 11237 37780
rect 11293 37724 11379 37780
rect 11435 37724 11521 37780
rect 11577 37724 11663 37780
rect 11719 37724 11805 37780
rect 11861 37724 11947 37780
rect 12003 37724 12089 37780
rect 12145 37724 12231 37780
rect 12287 37724 12373 37780
rect 12429 37724 12515 37780
rect 12571 37724 12657 37780
rect 12713 37724 12799 37780
rect 12855 37724 12941 37780
rect 12997 37724 13083 37780
rect 13139 37724 13225 37780
rect 13281 37724 13367 37780
rect 13423 37724 13509 37780
rect 13565 37724 13651 37780
rect 13707 37724 13793 37780
rect 13849 37724 13935 37780
rect 13991 37724 14077 37780
rect 14133 37724 14219 37780
rect 14275 37724 14361 37780
rect 14417 37724 14503 37780
rect 14559 37724 14645 37780
rect 14701 37724 14787 37780
rect 14843 37724 14853 37780
rect 151 37638 14853 37724
rect 151 37582 161 37638
rect 217 37582 303 37638
rect 359 37582 445 37638
rect 501 37582 587 37638
rect 643 37582 729 37638
rect 785 37582 871 37638
rect 927 37582 1013 37638
rect 1069 37582 1155 37638
rect 1211 37582 1297 37638
rect 1353 37582 1439 37638
rect 1495 37582 1581 37638
rect 1637 37582 1723 37638
rect 1779 37582 1865 37638
rect 1921 37582 2007 37638
rect 2063 37582 2149 37638
rect 2205 37582 2291 37638
rect 2347 37582 2433 37638
rect 2489 37582 2575 37638
rect 2631 37582 2717 37638
rect 2773 37582 2859 37638
rect 2915 37582 3001 37638
rect 3057 37582 3143 37638
rect 3199 37582 3285 37638
rect 3341 37582 3427 37638
rect 3483 37582 3569 37638
rect 3625 37582 3711 37638
rect 3767 37582 3853 37638
rect 3909 37582 3995 37638
rect 4051 37582 4137 37638
rect 4193 37582 4279 37638
rect 4335 37582 4421 37638
rect 4477 37582 4563 37638
rect 4619 37582 4705 37638
rect 4761 37582 4847 37638
rect 4903 37582 4989 37638
rect 5045 37582 5131 37638
rect 5187 37582 5273 37638
rect 5329 37582 5415 37638
rect 5471 37582 5557 37638
rect 5613 37582 5699 37638
rect 5755 37582 5841 37638
rect 5897 37582 5983 37638
rect 6039 37582 6125 37638
rect 6181 37582 6267 37638
rect 6323 37582 6409 37638
rect 6465 37582 6551 37638
rect 6607 37582 6693 37638
rect 6749 37582 6835 37638
rect 6891 37582 6977 37638
rect 7033 37582 7119 37638
rect 7175 37582 7261 37638
rect 7317 37582 7403 37638
rect 7459 37582 7545 37638
rect 7601 37582 7687 37638
rect 7743 37582 7829 37638
rect 7885 37582 7971 37638
rect 8027 37582 8113 37638
rect 8169 37582 8255 37638
rect 8311 37582 8397 37638
rect 8453 37582 8539 37638
rect 8595 37582 8681 37638
rect 8737 37582 8823 37638
rect 8879 37582 8965 37638
rect 9021 37582 9107 37638
rect 9163 37582 9249 37638
rect 9305 37582 9391 37638
rect 9447 37582 9533 37638
rect 9589 37582 9675 37638
rect 9731 37582 9817 37638
rect 9873 37582 9959 37638
rect 10015 37582 10101 37638
rect 10157 37582 10243 37638
rect 10299 37582 10385 37638
rect 10441 37582 10527 37638
rect 10583 37582 10669 37638
rect 10725 37582 10811 37638
rect 10867 37582 10953 37638
rect 11009 37582 11095 37638
rect 11151 37582 11237 37638
rect 11293 37582 11379 37638
rect 11435 37582 11521 37638
rect 11577 37582 11663 37638
rect 11719 37582 11805 37638
rect 11861 37582 11947 37638
rect 12003 37582 12089 37638
rect 12145 37582 12231 37638
rect 12287 37582 12373 37638
rect 12429 37582 12515 37638
rect 12571 37582 12657 37638
rect 12713 37582 12799 37638
rect 12855 37582 12941 37638
rect 12997 37582 13083 37638
rect 13139 37582 13225 37638
rect 13281 37582 13367 37638
rect 13423 37582 13509 37638
rect 13565 37582 13651 37638
rect 13707 37582 13793 37638
rect 13849 37582 13935 37638
rect 13991 37582 14077 37638
rect 14133 37582 14219 37638
rect 14275 37582 14361 37638
rect 14417 37582 14503 37638
rect 14559 37582 14645 37638
rect 14701 37582 14787 37638
rect 14843 37582 14853 37638
rect 151 37496 14853 37582
rect 151 37440 161 37496
rect 217 37440 303 37496
rect 359 37440 445 37496
rect 501 37440 587 37496
rect 643 37440 729 37496
rect 785 37440 871 37496
rect 927 37440 1013 37496
rect 1069 37440 1155 37496
rect 1211 37440 1297 37496
rect 1353 37440 1439 37496
rect 1495 37440 1581 37496
rect 1637 37440 1723 37496
rect 1779 37440 1865 37496
rect 1921 37440 2007 37496
rect 2063 37440 2149 37496
rect 2205 37440 2291 37496
rect 2347 37440 2433 37496
rect 2489 37440 2575 37496
rect 2631 37440 2717 37496
rect 2773 37440 2859 37496
rect 2915 37440 3001 37496
rect 3057 37440 3143 37496
rect 3199 37440 3285 37496
rect 3341 37440 3427 37496
rect 3483 37440 3569 37496
rect 3625 37440 3711 37496
rect 3767 37440 3853 37496
rect 3909 37440 3995 37496
rect 4051 37440 4137 37496
rect 4193 37440 4279 37496
rect 4335 37440 4421 37496
rect 4477 37440 4563 37496
rect 4619 37440 4705 37496
rect 4761 37440 4847 37496
rect 4903 37440 4989 37496
rect 5045 37440 5131 37496
rect 5187 37440 5273 37496
rect 5329 37440 5415 37496
rect 5471 37440 5557 37496
rect 5613 37440 5699 37496
rect 5755 37440 5841 37496
rect 5897 37440 5983 37496
rect 6039 37440 6125 37496
rect 6181 37440 6267 37496
rect 6323 37440 6409 37496
rect 6465 37440 6551 37496
rect 6607 37440 6693 37496
rect 6749 37440 6835 37496
rect 6891 37440 6977 37496
rect 7033 37440 7119 37496
rect 7175 37440 7261 37496
rect 7317 37440 7403 37496
rect 7459 37440 7545 37496
rect 7601 37440 7687 37496
rect 7743 37440 7829 37496
rect 7885 37440 7971 37496
rect 8027 37440 8113 37496
rect 8169 37440 8255 37496
rect 8311 37440 8397 37496
rect 8453 37440 8539 37496
rect 8595 37440 8681 37496
rect 8737 37440 8823 37496
rect 8879 37440 8965 37496
rect 9021 37440 9107 37496
rect 9163 37440 9249 37496
rect 9305 37440 9391 37496
rect 9447 37440 9533 37496
rect 9589 37440 9675 37496
rect 9731 37440 9817 37496
rect 9873 37440 9959 37496
rect 10015 37440 10101 37496
rect 10157 37440 10243 37496
rect 10299 37440 10385 37496
rect 10441 37440 10527 37496
rect 10583 37440 10669 37496
rect 10725 37440 10811 37496
rect 10867 37440 10953 37496
rect 11009 37440 11095 37496
rect 11151 37440 11237 37496
rect 11293 37440 11379 37496
rect 11435 37440 11521 37496
rect 11577 37440 11663 37496
rect 11719 37440 11805 37496
rect 11861 37440 11947 37496
rect 12003 37440 12089 37496
rect 12145 37440 12231 37496
rect 12287 37440 12373 37496
rect 12429 37440 12515 37496
rect 12571 37440 12657 37496
rect 12713 37440 12799 37496
rect 12855 37440 12941 37496
rect 12997 37440 13083 37496
rect 13139 37440 13225 37496
rect 13281 37440 13367 37496
rect 13423 37440 13509 37496
rect 13565 37440 13651 37496
rect 13707 37440 13793 37496
rect 13849 37440 13935 37496
rect 13991 37440 14077 37496
rect 14133 37440 14219 37496
rect 14275 37440 14361 37496
rect 14417 37440 14503 37496
rect 14559 37440 14645 37496
rect 14701 37440 14787 37496
rect 14843 37440 14853 37496
rect 151 37354 14853 37440
rect 151 37298 161 37354
rect 217 37298 303 37354
rect 359 37298 445 37354
rect 501 37298 587 37354
rect 643 37298 729 37354
rect 785 37298 871 37354
rect 927 37298 1013 37354
rect 1069 37298 1155 37354
rect 1211 37298 1297 37354
rect 1353 37298 1439 37354
rect 1495 37298 1581 37354
rect 1637 37298 1723 37354
rect 1779 37298 1865 37354
rect 1921 37298 2007 37354
rect 2063 37298 2149 37354
rect 2205 37298 2291 37354
rect 2347 37298 2433 37354
rect 2489 37298 2575 37354
rect 2631 37298 2717 37354
rect 2773 37298 2859 37354
rect 2915 37298 3001 37354
rect 3057 37298 3143 37354
rect 3199 37298 3285 37354
rect 3341 37298 3427 37354
rect 3483 37298 3569 37354
rect 3625 37298 3711 37354
rect 3767 37298 3853 37354
rect 3909 37298 3995 37354
rect 4051 37298 4137 37354
rect 4193 37298 4279 37354
rect 4335 37298 4421 37354
rect 4477 37298 4563 37354
rect 4619 37298 4705 37354
rect 4761 37298 4847 37354
rect 4903 37298 4989 37354
rect 5045 37298 5131 37354
rect 5187 37298 5273 37354
rect 5329 37298 5415 37354
rect 5471 37298 5557 37354
rect 5613 37298 5699 37354
rect 5755 37298 5841 37354
rect 5897 37298 5983 37354
rect 6039 37298 6125 37354
rect 6181 37298 6267 37354
rect 6323 37298 6409 37354
rect 6465 37298 6551 37354
rect 6607 37298 6693 37354
rect 6749 37298 6835 37354
rect 6891 37298 6977 37354
rect 7033 37298 7119 37354
rect 7175 37298 7261 37354
rect 7317 37298 7403 37354
rect 7459 37298 7545 37354
rect 7601 37298 7687 37354
rect 7743 37298 7829 37354
rect 7885 37298 7971 37354
rect 8027 37298 8113 37354
rect 8169 37298 8255 37354
rect 8311 37298 8397 37354
rect 8453 37298 8539 37354
rect 8595 37298 8681 37354
rect 8737 37298 8823 37354
rect 8879 37298 8965 37354
rect 9021 37298 9107 37354
rect 9163 37298 9249 37354
rect 9305 37298 9391 37354
rect 9447 37298 9533 37354
rect 9589 37298 9675 37354
rect 9731 37298 9817 37354
rect 9873 37298 9959 37354
rect 10015 37298 10101 37354
rect 10157 37298 10243 37354
rect 10299 37298 10385 37354
rect 10441 37298 10527 37354
rect 10583 37298 10669 37354
rect 10725 37298 10811 37354
rect 10867 37298 10953 37354
rect 11009 37298 11095 37354
rect 11151 37298 11237 37354
rect 11293 37298 11379 37354
rect 11435 37298 11521 37354
rect 11577 37298 11663 37354
rect 11719 37298 11805 37354
rect 11861 37298 11947 37354
rect 12003 37298 12089 37354
rect 12145 37298 12231 37354
rect 12287 37298 12373 37354
rect 12429 37298 12515 37354
rect 12571 37298 12657 37354
rect 12713 37298 12799 37354
rect 12855 37298 12941 37354
rect 12997 37298 13083 37354
rect 13139 37298 13225 37354
rect 13281 37298 13367 37354
rect 13423 37298 13509 37354
rect 13565 37298 13651 37354
rect 13707 37298 13793 37354
rect 13849 37298 13935 37354
rect 13991 37298 14077 37354
rect 14133 37298 14219 37354
rect 14275 37298 14361 37354
rect 14417 37298 14503 37354
rect 14559 37298 14645 37354
rect 14701 37298 14787 37354
rect 14843 37298 14853 37354
rect 151 37212 14853 37298
rect 151 37156 161 37212
rect 217 37156 303 37212
rect 359 37156 445 37212
rect 501 37156 587 37212
rect 643 37156 729 37212
rect 785 37156 871 37212
rect 927 37156 1013 37212
rect 1069 37156 1155 37212
rect 1211 37156 1297 37212
rect 1353 37156 1439 37212
rect 1495 37156 1581 37212
rect 1637 37156 1723 37212
rect 1779 37156 1865 37212
rect 1921 37156 2007 37212
rect 2063 37156 2149 37212
rect 2205 37156 2291 37212
rect 2347 37156 2433 37212
rect 2489 37156 2575 37212
rect 2631 37156 2717 37212
rect 2773 37156 2859 37212
rect 2915 37156 3001 37212
rect 3057 37156 3143 37212
rect 3199 37156 3285 37212
rect 3341 37156 3427 37212
rect 3483 37156 3569 37212
rect 3625 37156 3711 37212
rect 3767 37156 3853 37212
rect 3909 37156 3995 37212
rect 4051 37156 4137 37212
rect 4193 37156 4279 37212
rect 4335 37156 4421 37212
rect 4477 37156 4563 37212
rect 4619 37156 4705 37212
rect 4761 37156 4847 37212
rect 4903 37156 4989 37212
rect 5045 37156 5131 37212
rect 5187 37156 5273 37212
rect 5329 37156 5415 37212
rect 5471 37156 5557 37212
rect 5613 37156 5699 37212
rect 5755 37156 5841 37212
rect 5897 37156 5983 37212
rect 6039 37156 6125 37212
rect 6181 37156 6267 37212
rect 6323 37156 6409 37212
rect 6465 37156 6551 37212
rect 6607 37156 6693 37212
rect 6749 37156 6835 37212
rect 6891 37156 6977 37212
rect 7033 37156 7119 37212
rect 7175 37156 7261 37212
rect 7317 37156 7403 37212
rect 7459 37156 7545 37212
rect 7601 37156 7687 37212
rect 7743 37156 7829 37212
rect 7885 37156 7971 37212
rect 8027 37156 8113 37212
rect 8169 37156 8255 37212
rect 8311 37156 8397 37212
rect 8453 37156 8539 37212
rect 8595 37156 8681 37212
rect 8737 37156 8823 37212
rect 8879 37156 8965 37212
rect 9021 37156 9107 37212
rect 9163 37156 9249 37212
rect 9305 37156 9391 37212
rect 9447 37156 9533 37212
rect 9589 37156 9675 37212
rect 9731 37156 9817 37212
rect 9873 37156 9959 37212
rect 10015 37156 10101 37212
rect 10157 37156 10243 37212
rect 10299 37156 10385 37212
rect 10441 37156 10527 37212
rect 10583 37156 10669 37212
rect 10725 37156 10811 37212
rect 10867 37156 10953 37212
rect 11009 37156 11095 37212
rect 11151 37156 11237 37212
rect 11293 37156 11379 37212
rect 11435 37156 11521 37212
rect 11577 37156 11663 37212
rect 11719 37156 11805 37212
rect 11861 37156 11947 37212
rect 12003 37156 12089 37212
rect 12145 37156 12231 37212
rect 12287 37156 12373 37212
rect 12429 37156 12515 37212
rect 12571 37156 12657 37212
rect 12713 37156 12799 37212
rect 12855 37156 12941 37212
rect 12997 37156 13083 37212
rect 13139 37156 13225 37212
rect 13281 37156 13367 37212
rect 13423 37156 13509 37212
rect 13565 37156 13651 37212
rect 13707 37156 13793 37212
rect 13849 37156 13935 37212
rect 13991 37156 14077 37212
rect 14133 37156 14219 37212
rect 14275 37156 14361 37212
rect 14417 37156 14503 37212
rect 14559 37156 14645 37212
rect 14701 37156 14787 37212
rect 14843 37156 14853 37212
rect 151 37070 14853 37156
rect 151 37014 161 37070
rect 217 37014 303 37070
rect 359 37014 445 37070
rect 501 37014 587 37070
rect 643 37014 729 37070
rect 785 37014 871 37070
rect 927 37014 1013 37070
rect 1069 37014 1155 37070
rect 1211 37014 1297 37070
rect 1353 37014 1439 37070
rect 1495 37014 1581 37070
rect 1637 37014 1723 37070
rect 1779 37014 1865 37070
rect 1921 37014 2007 37070
rect 2063 37014 2149 37070
rect 2205 37014 2291 37070
rect 2347 37014 2433 37070
rect 2489 37014 2575 37070
rect 2631 37014 2717 37070
rect 2773 37014 2859 37070
rect 2915 37014 3001 37070
rect 3057 37014 3143 37070
rect 3199 37014 3285 37070
rect 3341 37014 3427 37070
rect 3483 37014 3569 37070
rect 3625 37014 3711 37070
rect 3767 37014 3853 37070
rect 3909 37014 3995 37070
rect 4051 37014 4137 37070
rect 4193 37014 4279 37070
rect 4335 37014 4421 37070
rect 4477 37014 4563 37070
rect 4619 37014 4705 37070
rect 4761 37014 4847 37070
rect 4903 37014 4989 37070
rect 5045 37014 5131 37070
rect 5187 37014 5273 37070
rect 5329 37014 5415 37070
rect 5471 37014 5557 37070
rect 5613 37014 5699 37070
rect 5755 37014 5841 37070
rect 5897 37014 5983 37070
rect 6039 37014 6125 37070
rect 6181 37014 6267 37070
rect 6323 37014 6409 37070
rect 6465 37014 6551 37070
rect 6607 37014 6693 37070
rect 6749 37014 6835 37070
rect 6891 37014 6977 37070
rect 7033 37014 7119 37070
rect 7175 37014 7261 37070
rect 7317 37014 7403 37070
rect 7459 37014 7545 37070
rect 7601 37014 7687 37070
rect 7743 37014 7829 37070
rect 7885 37014 7971 37070
rect 8027 37014 8113 37070
rect 8169 37014 8255 37070
rect 8311 37014 8397 37070
rect 8453 37014 8539 37070
rect 8595 37014 8681 37070
rect 8737 37014 8823 37070
rect 8879 37014 8965 37070
rect 9021 37014 9107 37070
rect 9163 37014 9249 37070
rect 9305 37014 9391 37070
rect 9447 37014 9533 37070
rect 9589 37014 9675 37070
rect 9731 37014 9817 37070
rect 9873 37014 9959 37070
rect 10015 37014 10101 37070
rect 10157 37014 10243 37070
rect 10299 37014 10385 37070
rect 10441 37014 10527 37070
rect 10583 37014 10669 37070
rect 10725 37014 10811 37070
rect 10867 37014 10953 37070
rect 11009 37014 11095 37070
rect 11151 37014 11237 37070
rect 11293 37014 11379 37070
rect 11435 37014 11521 37070
rect 11577 37014 11663 37070
rect 11719 37014 11805 37070
rect 11861 37014 11947 37070
rect 12003 37014 12089 37070
rect 12145 37014 12231 37070
rect 12287 37014 12373 37070
rect 12429 37014 12515 37070
rect 12571 37014 12657 37070
rect 12713 37014 12799 37070
rect 12855 37014 12941 37070
rect 12997 37014 13083 37070
rect 13139 37014 13225 37070
rect 13281 37014 13367 37070
rect 13423 37014 13509 37070
rect 13565 37014 13651 37070
rect 13707 37014 13793 37070
rect 13849 37014 13935 37070
rect 13991 37014 14077 37070
rect 14133 37014 14219 37070
rect 14275 37014 14361 37070
rect 14417 37014 14503 37070
rect 14559 37014 14645 37070
rect 14701 37014 14787 37070
rect 14843 37014 14853 37070
rect 151 36928 14853 37014
rect 151 36872 161 36928
rect 217 36872 303 36928
rect 359 36872 445 36928
rect 501 36872 587 36928
rect 643 36872 729 36928
rect 785 36872 871 36928
rect 927 36872 1013 36928
rect 1069 36872 1155 36928
rect 1211 36872 1297 36928
rect 1353 36872 1439 36928
rect 1495 36872 1581 36928
rect 1637 36872 1723 36928
rect 1779 36872 1865 36928
rect 1921 36872 2007 36928
rect 2063 36872 2149 36928
rect 2205 36872 2291 36928
rect 2347 36872 2433 36928
rect 2489 36872 2575 36928
rect 2631 36872 2717 36928
rect 2773 36872 2859 36928
rect 2915 36872 3001 36928
rect 3057 36872 3143 36928
rect 3199 36872 3285 36928
rect 3341 36872 3427 36928
rect 3483 36872 3569 36928
rect 3625 36872 3711 36928
rect 3767 36872 3853 36928
rect 3909 36872 3995 36928
rect 4051 36872 4137 36928
rect 4193 36872 4279 36928
rect 4335 36872 4421 36928
rect 4477 36872 4563 36928
rect 4619 36872 4705 36928
rect 4761 36872 4847 36928
rect 4903 36872 4989 36928
rect 5045 36872 5131 36928
rect 5187 36872 5273 36928
rect 5329 36872 5415 36928
rect 5471 36872 5557 36928
rect 5613 36872 5699 36928
rect 5755 36872 5841 36928
rect 5897 36872 5983 36928
rect 6039 36872 6125 36928
rect 6181 36872 6267 36928
rect 6323 36872 6409 36928
rect 6465 36872 6551 36928
rect 6607 36872 6693 36928
rect 6749 36872 6835 36928
rect 6891 36872 6977 36928
rect 7033 36872 7119 36928
rect 7175 36872 7261 36928
rect 7317 36872 7403 36928
rect 7459 36872 7545 36928
rect 7601 36872 7687 36928
rect 7743 36872 7829 36928
rect 7885 36872 7971 36928
rect 8027 36872 8113 36928
rect 8169 36872 8255 36928
rect 8311 36872 8397 36928
rect 8453 36872 8539 36928
rect 8595 36872 8681 36928
rect 8737 36872 8823 36928
rect 8879 36872 8965 36928
rect 9021 36872 9107 36928
rect 9163 36872 9249 36928
rect 9305 36872 9391 36928
rect 9447 36872 9533 36928
rect 9589 36872 9675 36928
rect 9731 36872 9817 36928
rect 9873 36872 9959 36928
rect 10015 36872 10101 36928
rect 10157 36872 10243 36928
rect 10299 36872 10385 36928
rect 10441 36872 10527 36928
rect 10583 36872 10669 36928
rect 10725 36872 10811 36928
rect 10867 36872 10953 36928
rect 11009 36872 11095 36928
rect 11151 36872 11237 36928
rect 11293 36872 11379 36928
rect 11435 36872 11521 36928
rect 11577 36872 11663 36928
rect 11719 36872 11805 36928
rect 11861 36872 11947 36928
rect 12003 36872 12089 36928
rect 12145 36872 12231 36928
rect 12287 36872 12373 36928
rect 12429 36872 12515 36928
rect 12571 36872 12657 36928
rect 12713 36872 12799 36928
rect 12855 36872 12941 36928
rect 12997 36872 13083 36928
rect 13139 36872 13225 36928
rect 13281 36872 13367 36928
rect 13423 36872 13509 36928
rect 13565 36872 13651 36928
rect 13707 36872 13793 36928
rect 13849 36872 13935 36928
rect 13991 36872 14077 36928
rect 14133 36872 14219 36928
rect 14275 36872 14361 36928
rect 14417 36872 14503 36928
rect 14559 36872 14645 36928
rect 14701 36872 14787 36928
rect 14843 36872 14853 36928
rect 151 36786 14853 36872
rect 151 36730 161 36786
rect 217 36730 303 36786
rect 359 36730 445 36786
rect 501 36730 587 36786
rect 643 36730 729 36786
rect 785 36730 871 36786
rect 927 36730 1013 36786
rect 1069 36730 1155 36786
rect 1211 36730 1297 36786
rect 1353 36730 1439 36786
rect 1495 36730 1581 36786
rect 1637 36730 1723 36786
rect 1779 36730 1865 36786
rect 1921 36730 2007 36786
rect 2063 36730 2149 36786
rect 2205 36730 2291 36786
rect 2347 36730 2433 36786
rect 2489 36730 2575 36786
rect 2631 36730 2717 36786
rect 2773 36730 2859 36786
rect 2915 36730 3001 36786
rect 3057 36730 3143 36786
rect 3199 36730 3285 36786
rect 3341 36730 3427 36786
rect 3483 36730 3569 36786
rect 3625 36730 3711 36786
rect 3767 36730 3853 36786
rect 3909 36730 3995 36786
rect 4051 36730 4137 36786
rect 4193 36730 4279 36786
rect 4335 36730 4421 36786
rect 4477 36730 4563 36786
rect 4619 36730 4705 36786
rect 4761 36730 4847 36786
rect 4903 36730 4989 36786
rect 5045 36730 5131 36786
rect 5187 36730 5273 36786
rect 5329 36730 5415 36786
rect 5471 36730 5557 36786
rect 5613 36730 5699 36786
rect 5755 36730 5841 36786
rect 5897 36730 5983 36786
rect 6039 36730 6125 36786
rect 6181 36730 6267 36786
rect 6323 36730 6409 36786
rect 6465 36730 6551 36786
rect 6607 36730 6693 36786
rect 6749 36730 6835 36786
rect 6891 36730 6977 36786
rect 7033 36730 7119 36786
rect 7175 36730 7261 36786
rect 7317 36730 7403 36786
rect 7459 36730 7545 36786
rect 7601 36730 7687 36786
rect 7743 36730 7829 36786
rect 7885 36730 7971 36786
rect 8027 36730 8113 36786
rect 8169 36730 8255 36786
rect 8311 36730 8397 36786
rect 8453 36730 8539 36786
rect 8595 36730 8681 36786
rect 8737 36730 8823 36786
rect 8879 36730 8965 36786
rect 9021 36730 9107 36786
rect 9163 36730 9249 36786
rect 9305 36730 9391 36786
rect 9447 36730 9533 36786
rect 9589 36730 9675 36786
rect 9731 36730 9817 36786
rect 9873 36730 9959 36786
rect 10015 36730 10101 36786
rect 10157 36730 10243 36786
rect 10299 36730 10385 36786
rect 10441 36730 10527 36786
rect 10583 36730 10669 36786
rect 10725 36730 10811 36786
rect 10867 36730 10953 36786
rect 11009 36730 11095 36786
rect 11151 36730 11237 36786
rect 11293 36730 11379 36786
rect 11435 36730 11521 36786
rect 11577 36730 11663 36786
rect 11719 36730 11805 36786
rect 11861 36730 11947 36786
rect 12003 36730 12089 36786
rect 12145 36730 12231 36786
rect 12287 36730 12373 36786
rect 12429 36730 12515 36786
rect 12571 36730 12657 36786
rect 12713 36730 12799 36786
rect 12855 36730 12941 36786
rect 12997 36730 13083 36786
rect 13139 36730 13225 36786
rect 13281 36730 13367 36786
rect 13423 36730 13509 36786
rect 13565 36730 13651 36786
rect 13707 36730 13793 36786
rect 13849 36730 13935 36786
rect 13991 36730 14077 36786
rect 14133 36730 14219 36786
rect 14275 36730 14361 36786
rect 14417 36730 14503 36786
rect 14559 36730 14645 36786
rect 14701 36730 14787 36786
rect 14843 36730 14853 36786
rect 151 36644 14853 36730
rect 151 36588 161 36644
rect 217 36588 303 36644
rect 359 36588 445 36644
rect 501 36588 587 36644
rect 643 36588 729 36644
rect 785 36588 871 36644
rect 927 36588 1013 36644
rect 1069 36588 1155 36644
rect 1211 36588 1297 36644
rect 1353 36588 1439 36644
rect 1495 36588 1581 36644
rect 1637 36588 1723 36644
rect 1779 36588 1865 36644
rect 1921 36588 2007 36644
rect 2063 36588 2149 36644
rect 2205 36588 2291 36644
rect 2347 36588 2433 36644
rect 2489 36588 2575 36644
rect 2631 36588 2717 36644
rect 2773 36588 2859 36644
rect 2915 36588 3001 36644
rect 3057 36588 3143 36644
rect 3199 36588 3285 36644
rect 3341 36588 3427 36644
rect 3483 36588 3569 36644
rect 3625 36588 3711 36644
rect 3767 36588 3853 36644
rect 3909 36588 3995 36644
rect 4051 36588 4137 36644
rect 4193 36588 4279 36644
rect 4335 36588 4421 36644
rect 4477 36588 4563 36644
rect 4619 36588 4705 36644
rect 4761 36588 4847 36644
rect 4903 36588 4989 36644
rect 5045 36588 5131 36644
rect 5187 36588 5273 36644
rect 5329 36588 5415 36644
rect 5471 36588 5557 36644
rect 5613 36588 5699 36644
rect 5755 36588 5841 36644
rect 5897 36588 5983 36644
rect 6039 36588 6125 36644
rect 6181 36588 6267 36644
rect 6323 36588 6409 36644
rect 6465 36588 6551 36644
rect 6607 36588 6693 36644
rect 6749 36588 6835 36644
rect 6891 36588 6977 36644
rect 7033 36588 7119 36644
rect 7175 36588 7261 36644
rect 7317 36588 7403 36644
rect 7459 36588 7545 36644
rect 7601 36588 7687 36644
rect 7743 36588 7829 36644
rect 7885 36588 7971 36644
rect 8027 36588 8113 36644
rect 8169 36588 8255 36644
rect 8311 36588 8397 36644
rect 8453 36588 8539 36644
rect 8595 36588 8681 36644
rect 8737 36588 8823 36644
rect 8879 36588 8965 36644
rect 9021 36588 9107 36644
rect 9163 36588 9249 36644
rect 9305 36588 9391 36644
rect 9447 36588 9533 36644
rect 9589 36588 9675 36644
rect 9731 36588 9817 36644
rect 9873 36588 9959 36644
rect 10015 36588 10101 36644
rect 10157 36588 10243 36644
rect 10299 36588 10385 36644
rect 10441 36588 10527 36644
rect 10583 36588 10669 36644
rect 10725 36588 10811 36644
rect 10867 36588 10953 36644
rect 11009 36588 11095 36644
rect 11151 36588 11237 36644
rect 11293 36588 11379 36644
rect 11435 36588 11521 36644
rect 11577 36588 11663 36644
rect 11719 36588 11805 36644
rect 11861 36588 11947 36644
rect 12003 36588 12089 36644
rect 12145 36588 12231 36644
rect 12287 36588 12373 36644
rect 12429 36588 12515 36644
rect 12571 36588 12657 36644
rect 12713 36588 12799 36644
rect 12855 36588 12941 36644
rect 12997 36588 13083 36644
rect 13139 36588 13225 36644
rect 13281 36588 13367 36644
rect 13423 36588 13509 36644
rect 13565 36588 13651 36644
rect 13707 36588 13793 36644
rect 13849 36588 13935 36644
rect 13991 36588 14077 36644
rect 14133 36588 14219 36644
rect 14275 36588 14361 36644
rect 14417 36588 14503 36644
rect 14559 36588 14645 36644
rect 14701 36588 14787 36644
rect 14843 36588 14853 36644
rect 151 36502 14853 36588
rect 151 36446 161 36502
rect 217 36446 303 36502
rect 359 36446 445 36502
rect 501 36446 587 36502
rect 643 36446 729 36502
rect 785 36446 871 36502
rect 927 36446 1013 36502
rect 1069 36446 1155 36502
rect 1211 36446 1297 36502
rect 1353 36446 1439 36502
rect 1495 36446 1581 36502
rect 1637 36446 1723 36502
rect 1779 36446 1865 36502
rect 1921 36446 2007 36502
rect 2063 36446 2149 36502
rect 2205 36446 2291 36502
rect 2347 36446 2433 36502
rect 2489 36446 2575 36502
rect 2631 36446 2717 36502
rect 2773 36446 2859 36502
rect 2915 36446 3001 36502
rect 3057 36446 3143 36502
rect 3199 36446 3285 36502
rect 3341 36446 3427 36502
rect 3483 36446 3569 36502
rect 3625 36446 3711 36502
rect 3767 36446 3853 36502
rect 3909 36446 3995 36502
rect 4051 36446 4137 36502
rect 4193 36446 4279 36502
rect 4335 36446 4421 36502
rect 4477 36446 4563 36502
rect 4619 36446 4705 36502
rect 4761 36446 4847 36502
rect 4903 36446 4989 36502
rect 5045 36446 5131 36502
rect 5187 36446 5273 36502
rect 5329 36446 5415 36502
rect 5471 36446 5557 36502
rect 5613 36446 5699 36502
rect 5755 36446 5841 36502
rect 5897 36446 5983 36502
rect 6039 36446 6125 36502
rect 6181 36446 6267 36502
rect 6323 36446 6409 36502
rect 6465 36446 6551 36502
rect 6607 36446 6693 36502
rect 6749 36446 6835 36502
rect 6891 36446 6977 36502
rect 7033 36446 7119 36502
rect 7175 36446 7261 36502
rect 7317 36446 7403 36502
rect 7459 36446 7545 36502
rect 7601 36446 7687 36502
rect 7743 36446 7829 36502
rect 7885 36446 7971 36502
rect 8027 36446 8113 36502
rect 8169 36446 8255 36502
rect 8311 36446 8397 36502
rect 8453 36446 8539 36502
rect 8595 36446 8681 36502
rect 8737 36446 8823 36502
rect 8879 36446 8965 36502
rect 9021 36446 9107 36502
rect 9163 36446 9249 36502
rect 9305 36446 9391 36502
rect 9447 36446 9533 36502
rect 9589 36446 9675 36502
rect 9731 36446 9817 36502
rect 9873 36446 9959 36502
rect 10015 36446 10101 36502
rect 10157 36446 10243 36502
rect 10299 36446 10385 36502
rect 10441 36446 10527 36502
rect 10583 36446 10669 36502
rect 10725 36446 10811 36502
rect 10867 36446 10953 36502
rect 11009 36446 11095 36502
rect 11151 36446 11237 36502
rect 11293 36446 11379 36502
rect 11435 36446 11521 36502
rect 11577 36446 11663 36502
rect 11719 36446 11805 36502
rect 11861 36446 11947 36502
rect 12003 36446 12089 36502
rect 12145 36446 12231 36502
rect 12287 36446 12373 36502
rect 12429 36446 12515 36502
rect 12571 36446 12657 36502
rect 12713 36446 12799 36502
rect 12855 36446 12941 36502
rect 12997 36446 13083 36502
rect 13139 36446 13225 36502
rect 13281 36446 13367 36502
rect 13423 36446 13509 36502
rect 13565 36446 13651 36502
rect 13707 36446 13793 36502
rect 13849 36446 13935 36502
rect 13991 36446 14077 36502
rect 14133 36446 14219 36502
rect 14275 36446 14361 36502
rect 14417 36446 14503 36502
rect 14559 36446 14645 36502
rect 14701 36446 14787 36502
rect 14843 36446 14853 36502
rect 151 36436 14853 36446
rect 151 36142 14853 36152
rect 151 36086 161 36142
rect 217 36086 303 36142
rect 359 36086 445 36142
rect 501 36086 587 36142
rect 643 36086 729 36142
rect 785 36086 871 36142
rect 927 36086 1013 36142
rect 1069 36086 1155 36142
rect 1211 36086 1297 36142
rect 1353 36086 1439 36142
rect 1495 36086 1581 36142
rect 1637 36086 1723 36142
rect 1779 36086 1865 36142
rect 1921 36086 2007 36142
rect 2063 36086 2149 36142
rect 2205 36086 2291 36142
rect 2347 36086 2433 36142
rect 2489 36086 2575 36142
rect 2631 36086 2717 36142
rect 2773 36086 2859 36142
rect 2915 36086 3001 36142
rect 3057 36086 3143 36142
rect 3199 36086 3285 36142
rect 3341 36086 3427 36142
rect 3483 36086 3569 36142
rect 3625 36086 3711 36142
rect 3767 36086 3853 36142
rect 3909 36086 3995 36142
rect 4051 36086 4137 36142
rect 4193 36086 4279 36142
rect 4335 36086 4421 36142
rect 4477 36086 4563 36142
rect 4619 36086 4705 36142
rect 4761 36086 4847 36142
rect 4903 36086 4989 36142
rect 5045 36086 5131 36142
rect 5187 36086 5273 36142
rect 5329 36086 5415 36142
rect 5471 36086 5557 36142
rect 5613 36086 5699 36142
rect 5755 36086 5841 36142
rect 5897 36086 5983 36142
rect 6039 36086 6125 36142
rect 6181 36086 6267 36142
rect 6323 36086 6409 36142
rect 6465 36086 6551 36142
rect 6607 36086 6693 36142
rect 6749 36086 6835 36142
rect 6891 36086 6977 36142
rect 7033 36086 7119 36142
rect 7175 36086 7261 36142
rect 7317 36086 7403 36142
rect 7459 36086 7545 36142
rect 7601 36086 7687 36142
rect 7743 36086 7829 36142
rect 7885 36086 7971 36142
rect 8027 36086 8113 36142
rect 8169 36086 8255 36142
rect 8311 36086 8397 36142
rect 8453 36086 8539 36142
rect 8595 36086 8681 36142
rect 8737 36086 8823 36142
rect 8879 36086 8965 36142
rect 9021 36086 9107 36142
rect 9163 36086 9249 36142
rect 9305 36086 9391 36142
rect 9447 36086 9533 36142
rect 9589 36086 9675 36142
rect 9731 36086 9817 36142
rect 9873 36086 9959 36142
rect 10015 36086 10101 36142
rect 10157 36086 10243 36142
rect 10299 36086 10385 36142
rect 10441 36086 10527 36142
rect 10583 36086 10669 36142
rect 10725 36086 10811 36142
rect 10867 36086 10953 36142
rect 11009 36086 11095 36142
rect 11151 36086 11237 36142
rect 11293 36086 11379 36142
rect 11435 36086 11521 36142
rect 11577 36086 11663 36142
rect 11719 36086 11805 36142
rect 11861 36086 11947 36142
rect 12003 36086 12089 36142
rect 12145 36086 12231 36142
rect 12287 36086 12373 36142
rect 12429 36086 12515 36142
rect 12571 36086 12657 36142
rect 12713 36086 12799 36142
rect 12855 36086 12941 36142
rect 12997 36086 13083 36142
rect 13139 36086 13225 36142
rect 13281 36086 13367 36142
rect 13423 36086 13509 36142
rect 13565 36086 13651 36142
rect 13707 36086 13793 36142
rect 13849 36086 13935 36142
rect 13991 36086 14077 36142
rect 14133 36086 14219 36142
rect 14275 36086 14361 36142
rect 14417 36086 14503 36142
rect 14559 36086 14645 36142
rect 14701 36086 14787 36142
rect 14843 36086 14853 36142
rect 151 36000 14853 36086
rect 151 35944 161 36000
rect 217 35944 303 36000
rect 359 35944 445 36000
rect 501 35944 587 36000
rect 643 35944 729 36000
rect 785 35944 871 36000
rect 927 35944 1013 36000
rect 1069 35944 1155 36000
rect 1211 35944 1297 36000
rect 1353 35944 1439 36000
rect 1495 35944 1581 36000
rect 1637 35944 1723 36000
rect 1779 35944 1865 36000
rect 1921 35944 2007 36000
rect 2063 35944 2149 36000
rect 2205 35944 2291 36000
rect 2347 35944 2433 36000
rect 2489 35944 2575 36000
rect 2631 35944 2717 36000
rect 2773 35944 2859 36000
rect 2915 35944 3001 36000
rect 3057 35944 3143 36000
rect 3199 35944 3285 36000
rect 3341 35944 3427 36000
rect 3483 35944 3569 36000
rect 3625 35944 3711 36000
rect 3767 35944 3853 36000
rect 3909 35944 3995 36000
rect 4051 35944 4137 36000
rect 4193 35944 4279 36000
rect 4335 35944 4421 36000
rect 4477 35944 4563 36000
rect 4619 35944 4705 36000
rect 4761 35944 4847 36000
rect 4903 35944 4989 36000
rect 5045 35944 5131 36000
rect 5187 35944 5273 36000
rect 5329 35944 5415 36000
rect 5471 35944 5557 36000
rect 5613 35944 5699 36000
rect 5755 35944 5841 36000
rect 5897 35944 5983 36000
rect 6039 35944 6125 36000
rect 6181 35944 6267 36000
rect 6323 35944 6409 36000
rect 6465 35944 6551 36000
rect 6607 35944 6693 36000
rect 6749 35944 6835 36000
rect 6891 35944 6977 36000
rect 7033 35944 7119 36000
rect 7175 35944 7261 36000
rect 7317 35944 7403 36000
rect 7459 35944 7545 36000
rect 7601 35944 7687 36000
rect 7743 35944 7829 36000
rect 7885 35944 7971 36000
rect 8027 35944 8113 36000
rect 8169 35944 8255 36000
rect 8311 35944 8397 36000
rect 8453 35944 8539 36000
rect 8595 35944 8681 36000
rect 8737 35944 8823 36000
rect 8879 35944 8965 36000
rect 9021 35944 9107 36000
rect 9163 35944 9249 36000
rect 9305 35944 9391 36000
rect 9447 35944 9533 36000
rect 9589 35944 9675 36000
rect 9731 35944 9817 36000
rect 9873 35944 9959 36000
rect 10015 35944 10101 36000
rect 10157 35944 10243 36000
rect 10299 35944 10385 36000
rect 10441 35944 10527 36000
rect 10583 35944 10669 36000
rect 10725 35944 10811 36000
rect 10867 35944 10953 36000
rect 11009 35944 11095 36000
rect 11151 35944 11237 36000
rect 11293 35944 11379 36000
rect 11435 35944 11521 36000
rect 11577 35944 11663 36000
rect 11719 35944 11805 36000
rect 11861 35944 11947 36000
rect 12003 35944 12089 36000
rect 12145 35944 12231 36000
rect 12287 35944 12373 36000
rect 12429 35944 12515 36000
rect 12571 35944 12657 36000
rect 12713 35944 12799 36000
rect 12855 35944 12941 36000
rect 12997 35944 13083 36000
rect 13139 35944 13225 36000
rect 13281 35944 13367 36000
rect 13423 35944 13509 36000
rect 13565 35944 13651 36000
rect 13707 35944 13793 36000
rect 13849 35944 13935 36000
rect 13991 35944 14077 36000
rect 14133 35944 14219 36000
rect 14275 35944 14361 36000
rect 14417 35944 14503 36000
rect 14559 35944 14645 36000
rect 14701 35944 14787 36000
rect 14843 35944 14853 36000
rect 151 35858 14853 35944
rect 151 35802 161 35858
rect 217 35802 303 35858
rect 359 35802 445 35858
rect 501 35802 587 35858
rect 643 35802 729 35858
rect 785 35802 871 35858
rect 927 35802 1013 35858
rect 1069 35802 1155 35858
rect 1211 35802 1297 35858
rect 1353 35802 1439 35858
rect 1495 35802 1581 35858
rect 1637 35802 1723 35858
rect 1779 35802 1865 35858
rect 1921 35802 2007 35858
rect 2063 35802 2149 35858
rect 2205 35802 2291 35858
rect 2347 35802 2433 35858
rect 2489 35802 2575 35858
rect 2631 35802 2717 35858
rect 2773 35802 2859 35858
rect 2915 35802 3001 35858
rect 3057 35802 3143 35858
rect 3199 35802 3285 35858
rect 3341 35802 3427 35858
rect 3483 35802 3569 35858
rect 3625 35802 3711 35858
rect 3767 35802 3853 35858
rect 3909 35802 3995 35858
rect 4051 35802 4137 35858
rect 4193 35802 4279 35858
rect 4335 35802 4421 35858
rect 4477 35802 4563 35858
rect 4619 35802 4705 35858
rect 4761 35802 4847 35858
rect 4903 35802 4989 35858
rect 5045 35802 5131 35858
rect 5187 35802 5273 35858
rect 5329 35802 5415 35858
rect 5471 35802 5557 35858
rect 5613 35802 5699 35858
rect 5755 35802 5841 35858
rect 5897 35802 5983 35858
rect 6039 35802 6125 35858
rect 6181 35802 6267 35858
rect 6323 35802 6409 35858
rect 6465 35802 6551 35858
rect 6607 35802 6693 35858
rect 6749 35802 6835 35858
rect 6891 35802 6977 35858
rect 7033 35802 7119 35858
rect 7175 35802 7261 35858
rect 7317 35802 7403 35858
rect 7459 35802 7545 35858
rect 7601 35802 7687 35858
rect 7743 35802 7829 35858
rect 7885 35802 7971 35858
rect 8027 35802 8113 35858
rect 8169 35802 8255 35858
rect 8311 35802 8397 35858
rect 8453 35802 8539 35858
rect 8595 35802 8681 35858
rect 8737 35802 8823 35858
rect 8879 35802 8965 35858
rect 9021 35802 9107 35858
rect 9163 35802 9249 35858
rect 9305 35802 9391 35858
rect 9447 35802 9533 35858
rect 9589 35802 9675 35858
rect 9731 35802 9817 35858
rect 9873 35802 9959 35858
rect 10015 35802 10101 35858
rect 10157 35802 10243 35858
rect 10299 35802 10385 35858
rect 10441 35802 10527 35858
rect 10583 35802 10669 35858
rect 10725 35802 10811 35858
rect 10867 35802 10953 35858
rect 11009 35802 11095 35858
rect 11151 35802 11237 35858
rect 11293 35802 11379 35858
rect 11435 35802 11521 35858
rect 11577 35802 11663 35858
rect 11719 35802 11805 35858
rect 11861 35802 11947 35858
rect 12003 35802 12089 35858
rect 12145 35802 12231 35858
rect 12287 35802 12373 35858
rect 12429 35802 12515 35858
rect 12571 35802 12657 35858
rect 12713 35802 12799 35858
rect 12855 35802 12941 35858
rect 12997 35802 13083 35858
rect 13139 35802 13225 35858
rect 13281 35802 13367 35858
rect 13423 35802 13509 35858
rect 13565 35802 13651 35858
rect 13707 35802 13793 35858
rect 13849 35802 13935 35858
rect 13991 35802 14077 35858
rect 14133 35802 14219 35858
rect 14275 35802 14361 35858
rect 14417 35802 14503 35858
rect 14559 35802 14645 35858
rect 14701 35802 14787 35858
rect 14843 35802 14853 35858
rect 151 35716 14853 35802
rect 151 35660 161 35716
rect 217 35660 303 35716
rect 359 35660 445 35716
rect 501 35660 587 35716
rect 643 35660 729 35716
rect 785 35660 871 35716
rect 927 35660 1013 35716
rect 1069 35660 1155 35716
rect 1211 35660 1297 35716
rect 1353 35660 1439 35716
rect 1495 35660 1581 35716
rect 1637 35660 1723 35716
rect 1779 35660 1865 35716
rect 1921 35660 2007 35716
rect 2063 35660 2149 35716
rect 2205 35660 2291 35716
rect 2347 35660 2433 35716
rect 2489 35660 2575 35716
rect 2631 35660 2717 35716
rect 2773 35660 2859 35716
rect 2915 35660 3001 35716
rect 3057 35660 3143 35716
rect 3199 35660 3285 35716
rect 3341 35660 3427 35716
rect 3483 35660 3569 35716
rect 3625 35660 3711 35716
rect 3767 35660 3853 35716
rect 3909 35660 3995 35716
rect 4051 35660 4137 35716
rect 4193 35660 4279 35716
rect 4335 35660 4421 35716
rect 4477 35660 4563 35716
rect 4619 35660 4705 35716
rect 4761 35660 4847 35716
rect 4903 35660 4989 35716
rect 5045 35660 5131 35716
rect 5187 35660 5273 35716
rect 5329 35660 5415 35716
rect 5471 35660 5557 35716
rect 5613 35660 5699 35716
rect 5755 35660 5841 35716
rect 5897 35660 5983 35716
rect 6039 35660 6125 35716
rect 6181 35660 6267 35716
rect 6323 35660 6409 35716
rect 6465 35660 6551 35716
rect 6607 35660 6693 35716
rect 6749 35660 6835 35716
rect 6891 35660 6977 35716
rect 7033 35660 7119 35716
rect 7175 35660 7261 35716
rect 7317 35660 7403 35716
rect 7459 35660 7545 35716
rect 7601 35660 7687 35716
rect 7743 35660 7829 35716
rect 7885 35660 7971 35716
rect 8027 35660 8113 35716
rect 8169 35660 8255 35716
rect 8311 35660 8397 35716
rect 8453 35660 8539 35716
rect 8595 35660 8681 35716
rect 8737 35660 8823 35716
rect 8879 35660 8965 35716
rect 9021 35660 9107 35716
rect 9163 35660 9249 35716
rect 9305 35660 9391 35716
rect 9447 35660 9533 35716
rect 9589 35660 9675 35716
rect 9731 35660 9817 35716
rect 9873 35660 9959 35716
rect 10015 35660 10101 35716
rect 10157 35660 10243 35716
rect 10299 35660 10385 35716
rect 10441 35660 10527 35716
rect 10583 35660 10669 35716
rect 10725 35660 10811 35716
rect 10867 35660 10953 35716
rect 11009 35660 11095 35716
rect 11151 35660 11237 35716
rect 11293 35660 11379 35716
rect 11435 35660 11521 35716
rect 11577 35660 11663 35716
rect 11719 35660 11805 35716
rect 11861 35660 11947 35716
rect 12003 35660 12089 35716
rect 12145 35660 12231 35716
rect 12287 35660 12373 35716
rect 12429 35660 12515 35716
rect 12571 35660 12657 35716
rect 12713 35660 12799 35716
rect 12855 35660 12941 35716
rect 12997 35660 13083 35716
rect 13139 35660 13225 35716
rect 13281 35660 13367 35716
rect 13423 35660 13509 35716
rect 13565 35660 13651 35716
rect 13707 35660 13793 35716
rect 13849 35660 13935 35716
rect 13991 35660 14077 35716
rect 14133 35660 14219 35716
rect 14275 35660 14361 35716
rect 14417 35660 14503 35716
rect 14559 35660 14645 35716
rect 14701 35660 14787 35716
rect 14843 35660 14853 35716
rect 151 35574 14853 35660
rect 151 35518 161 35574
rect 217 35518 303 35574
rect 359 35518 445 35574
rect 501 35518 587 35574
rect 643 35518 729 35574
rect 785 35518 871 35574
rect 927 35518 1013 35574
rect 1069 35518 1155 35574
rect 1211 35518 1297 35574
rect 1353 35518 1439 35574
rect 1495 35518 1581 35574
rect 1637 35518 1723 35574
rect 1779 35518 1865 35574
rect 1921 35518 2007 35574
rect 2063 35518 2149 35574
rect 2205 35518 2291 35574
rect 2347 35518 2433 35574
rect 2489 35518 2575 35574
rect 2631 35518 2717 35574
rect 2773 35518 2859 35574
rect 2915 35518 3001 35574
rect 3057 35518 3143 35574
rect 3199 35518 3285 35574
rect 3341 35518 3427 35574
rect 3483 35518 3569 35574
rect 3625 35518 3711 35574
rect 3767 35518 3853 35574
rect 3909 35518 3995 35574
rect 4051 35518 4137 35574
rect 4193 35518 4279 35574
rect 4335 35518 4421 35574
rect 4477 35518 4563 35574
rect 4619 35518 4705 35574
rect 4761 35518 4847 35574
rect 4903 35518 4989 35574
rect 5045 35518 5131 35574
rect 5187 35518 5273 35574
rect 5329 35518 5415 35574
rect 5471 35518 5557 35574
rect 5613 35518 5699 35574
rect 5755 35518 5841 35574
rect 5897 35518 5983 35574
rect 6039 35518 6125 35574
rect 6181 35518 6267 35574
rect 6323 35518 6409 35574
rect 6465 35518 6551 35574
rect 6607 35518 6693 35574
rect 6749 35518 6835 35574
rect 6891 35518 6977 35574
rect 7033 35518 7119 35574
rect 7175 35518 7261 35574
rect 7317 35518 7403 35574
rect 7459 35518 7545 35574
rect 7601 35518 7687 35574
rect 7743 35518 7829 35574
rect 7885 35518 7971 35574
rect 8027 35518 8113 35574
rect 8169 35518 8255 35574
rect 8311 35518 8397 35574
rect 8453 35518 8539 35574
rect 8595 35518 8681 35574
rect 8737 35518 8823 35574
rect 8879 35518 8965 35574
rect 9021 35518 9107 35574
rect 9163 35518 9249 35574
rect 9305 35518 9391 35574
rect 9447 35518 9533 35574
rect 9589 35518 9675 35574
rect 9731 35518 9817 35574
rect 9873 35518 9959 35574
rect 10015 35518 10101 35574
rect 10157 35518 10243 35574
rect 10299 35518 10385 35574
rect 10441 35518 10527 35574
rect 10583 35518 10669 35574
rect 10725 35518 10811 35574
rect 10867 35518 10953 35574
rect 11009 35518 11095 35574
rect 11151 35518 11237 35574
rect 11293 35518 11379 35574
rect 11435 35518 11521 35574
rect 11577 35518 11663 35574
rect 11719 35518 11805 35574
rect 11861 35518 11947 35574
rect 12003 35518 12089 35574
rect 12145 35518 12231 35574
rect 12287 35518 12373 35574
rect 12429 35518 12515 35574
rect 12571 35518 12657 35574
rect 12713 35518 12799 35574
rect 12855 35518 12941 35574
rect 12997 35518 13083 35574
rect 13139 35518 13225 35574
rect 13281 35518 13367 35574
rect 13423 35518 13509 35574
rect 13565 35518 13651 35574
rect 13707 35518 13793 35574
rect 13849 35518 13935 35574
rect 13991 35518 14077 35574
rect 14133 35518 14219 35574
rect 14275 35518 14361 35574
rect 14417 35518 14503 35574
rect 14559 35518 14645 35574
rect 14701 35518 14787 35574
rect 14843 35518 14853 35574
rect 151 35432 14853 35518
rect 151 35376 161 35432
rect 217 35376 303 35432
rect 359 35376 445 35432
rect 501 35376 587 35432
rect 643 35376 729 35432
rect 785 35376 871 35432
rect 927 35376 1013 35432
rect 1069 35376 1155 35432
rect 1211 35376 1297 35432
rect 1353 35376 1439 35432
rect 1495 35376 1581 35432
rect 1637 35376 1723 35432
rect 1779 35376 1865 35432
rect 1921 35376 2007 35432
rect 2063 35376 2149 35432
rect 2205 35376 2291 35432
rect 2347 35376 2433 35432
rect 2489 35376 2575 35432
rect 2631 35376 2717 35432
rect 2773 35376 2859 35432
rect 2915 35376 3001 35432
rect 3057 35376 3143 35432
rect 3199 35376 3285 35432
rect 3341 35376 3427 35432
rect 3483 35376 3569 35432
rect 3625 35376 3711 35432
rect 3767 35376 3853 35432
rect 3909 35376 3995 35432
rect 4051 35376 4137 35432
rect 4193 35376 4279 35432
rect 4335 35376 4421 35432
rect 4477 35376 4563 35432
rect 4619 35376 4705 35432
rect 4761 35376 4847 35432
rect 4903 35376 4989 35432
rect 5045 35376 5131 35432
rect 5187 35376 5273 35432
rect 5329 35376 5415 35432
rect 5471 35376 5557 35432
rect 5613 35376 5699 35432
rect 5755 35376 5841 35432
rect 5897 35376 5983 35432
rect 6039 35376 6125 35432
rect 6181 35376 6267 35432
rect 6323 35376 6409 35432
rect 6465 35376 6551 35432
rect 6607 35376 6693 35432
rect 6749 35376 6835 35432
rect 6891 35376 6977 35432
rect 7033 35376 7119 35432
rect 7175 35376 7261 35432
rect 7317 35376 7403 35432
rect 7459 35376 7545 35432
rect 7601 35376 7687 35432
rect 7743 35376 7829 35432
rect 7885 35376 7971 35432
rect 8027 35376 8113 35432
rect 8169 35376 8255 35432
rect 8311 35376 8397 35432
rect 8453 35376 8539 35432
rect 8595 35376 8681 35432
rect 8737 35376 8823 35432
rect 8879 35376 8965 35432
rect 9021 35376 9107 35432
rect 9163 35376 9249 35432
rect 9305 35376 9391 35432
rect 9447 35376 9533 35432
rect 9589 35376 9675 35432
rect 9731 35376 9817 35432
rect 9873 35376 9959 35432
rect 10015 35376 10101 35432
rect 10157 35376 10243 35432
rect 10299 35376 10385 35432
rect 10441 35376 10527 35432
rect 10583 35376 10669 35432
rect 10725 35376 10811 35432
rect 10867 35376 10953 35432
rect 11009 35376 11095 35432
rect 11151 35376 11237 35432
rect 11293 35376 11379 35432
rect 11435 35376 11521 35432
rect 11577 35376 11663 35432
rect 11719 35376 11805 35432
rect 11861 35376 11947 35432
rect 12003 35376 12089 35432
rect 12145 35376 12231 35432
rect 12287 35376 12373 35432
rect 12429 35376 12515 35432
rect 12571 35376 12657 35432
rect 12713 35376 12799 35432
rect 12855 35376 12941 35432
rect 12997 35376 13083 35432
rect 13139 35376 13225 35432
rect 13281 35376 13367 35432
rect 13423 35376 13509 35432
rect 13565 35376 13651 35432
rect 13707 35376 13793 35432
rect 13849 35376 13935 35432
rect 13991 35376 14077 35432
rect 14133 35376 14219 35432
rect 14275 35376 14361 35432
rect 14417 35376 14503 35432
rect 14559 35376 14645 35432
rect 14701 35376 14787 35432
rect 14843 35376 14853 35432
rect 151 35290 14853 35376
rect 151 35234 161 35290
rect 217 35234 303 35290
rect 359 35234 445 35290
rect 501 35234 587 35290
rect 643 35234 729 35290
rect 785 35234 871 35290
rect 927 35234 1013 35290
rect 1069 35234 1155 35290
rect 1211 35234 1297 35290
rect 1353 35234 1439 35290
rect 1495 35234 1581 35290
rect 1637 35234 1723 35290
rect 1779 35234 1865 35290
rect 1921 35234 2007 35290
rect 2063 35234 2149 35290
rect 2205 35234 2291 35290
rect 2347 35234 2433 35290
rect 2489 35234 2575 35290
rect 2631 35234 2717 35290
rect 2773 35234 2859 35290
rect 2915 35234 3001 35290
rect 3057 35234 3143 35290
rect 3199 35234 3285 35290
rect 3341 35234 3427 35290
rect 3483 35234 3569 35290
rect 3625 35234 3711 35290
rect 3767 35234 3853 35290
rect 3909 35234 3995 35290
rect 4051 35234 4137 35290
rect 4193 35234 4279 35290
rect 4335 35234 4421 35290
rect 4477 35234 4563 35290
rect 4619 35234 4705 35290
rect 4761 35234 4847 35290
rect 4903 35234 4989 35290
rect 5045 35234 5131 35290
rect 5187 35234 5273 35290
rect 5329 35234 5415 35290
rect 5471 35234 5557 35290
rect 5613 35234 5699 35290
rect 5755 35234 5841 35290
rect 5897 35234 5983 35290
rect 6039 35234 6125 35290
rect 6181 35234 6267 35290
rect 6323 35234 6409 35290
rect 6465 35234 6551 35290
rect 6607 35234 6693 35290
rect 6749 35234 6835 35290
rect 6891 35234 6977 35290
rect 7033 35234 7119 35290
rect 7175 35234 7261 35290
rect 7317 35234 7403 35290
rect 7459 35234 7545 35290
rect 7601 35234 7687 35290
rect 7743 35234 7829 35290
rect 7885 35234 7971 35290
rect 8027 35234 8113 35290
rect 8169 35234 8255 35290
rect 8311 35234 8397 35290
rect 8453 35234 8539 35290
rect 8595 35234 8681 35290
rect 8737 35234 8823 35290
rect 8879 35234 8965 35290
rect 9021 35234 9107 35290
rect 9163 35234 9249 35290
rect 9305 35234 9391 35290
rect 9447 35234 9533 35290
rect 9589 35234 9675 35290
rect 9731 35234 9817 35290
rect 9873 35234 9959 35290
rect 10015 35234 10101 35290
rect 10157 35234 10243 35290
rect 10299 35234 10385 35290
rect 10441 35234 10527 35290
rect 10583 35234 10669 35290
rect 10725 35234 10811 35290
rect 10867 35234 10953 35290
rect 11009 35234 11095 35290
rect 11151 35234 11237 35290
rect 11293 35234 11379 35290
rect 11435 35234 11521 35290
rect 11577 35234 11663 35290
rect 11719 35234 11805 35290
rect 11861 35234 11947 35290
rect 12003 35234 12089 35290
rect 12145 35234 12231 35290
rect 12287 35234 12373 35290
rect 12429 35234 12515 35290
rect 12571 35234 12657 35290
rect 12713 35234 12799 35290
rect 12855 35234 12941 35290
rect 12997 35234 13083 35290
rect 13139 35234 13225 35290
rect 13281 35234 13367 35290
rect 13423 35234 13509 35290
rect 13565 35234 13651 35290
rect 13707 35234 13793 35290
rect 13849 35234 13935 35290
rect 13991 35234 14077 35290
rect 14133 35234 14219 35290
rect 14275 35234 14361 35290
rect 14417 35234 14503 35290
rect 14559 35234 14645 35290
rect 14701 35234 14787 35290
rect 14843 35234 14853 35290
rect 151 35148 14853 35234
rect 151 35092 161 35148
rect 217 35092 303 35148
rect 359 35092 445 35148
rect 501 35092 587 35148
rect 643 35092 729 35148
rect 785 35092 871 35148
rect 927 35092 1013 35148
rect 1069 35092 1155 35148
rect 1211 35092 1297 35148
rect 1353 35092 1439 35148
rect 1495 35092 1581 35148
rect 1637 35092 1723 35148
rect 1779 35092 1865 35148
rect 1921 35092 2007 35148
rect 2063 35092 2149 35148
rect 2205 35092 2291 35148
rect 2347 35092 2433 35148
rect 2489 35092 2575 35148
rect 2631 35092 2717 35148
rect 2773 35092 2859 35148
rect 2915 35092 3001 35148
rect 3057 35092 3143 35148
rect 3199 35092 3285 35148
rect 3341 35092 3427 35148
rect 3483 35092 3569 35148
rect 3625 35092 3711 35148
rect 3767 35092 3853 35148
rect 3909 35092 3995 35148
rect 4051 35092 4137 35148
rect 4193 35092 4279 35148
rect 4335 35092 4421 35148
rect 4477 35092 4563 35148
rect 4619 35092 4705 35148
rect 4761 35092 4847 35148
rect 4903 35092 4989 35148
rect 5045 35092 5131 35148
rect 5187 35092 5273 35148
rect 5329 35092 5415 35148
rect 5471 35092 5557 35148
rect 5613 35092 5699 35148
rect 5755 35092 5841 35148
rect 5897 35092 5983 35148
rect 6039 35092 6125 35148
rect 6181 35092 6267 35148
rect 6323 35092 6409 35148
rect 6465 35092 6551 35148
rect 6607 35092 6693 35148
rect 6749 35092 6835 35148
rect 6891 35092 6977 35148
rect 7033 35092 7119 35148
rect 7175 35092 7261 35148
rect 7317 35092 7403 35148
rect 7459 35092 7545 35148
rect 7601 35092 7687 35148
rect 7743 35092 7829 35148
rect 7885 35092 7971 35148
rect 8027 35092 8113 35148
rect 8169 35092 8255 35148
rect 8311 35092 8397 35148
rect 8453 35092 8539 35148
rect 8595 35092 8681 35148
rect 8737 35092 8823 35148
rect 8879 35092 8965 35148
rect 9021 35092 9107 35148
rect 9163 35092 9249 35148
rect 9305 35092 9391 35148
rect 9447 35092 9533 35148
rect 9589 35092 9675 35148
rect 9731 35092 9817 35148
rect 9873 35092 9959 35148
rect 10015 35092 10101 35148
rect 10157 35092 10243 35148
rect 10299 35092 10385 35148
rect 10441 35092 10527 35148
rect 10583 35092 10669 35148
rect 10725 35092 10811 35148
rect 10867 35092 10953 35148
rect 11009 35092 11095 35148
rect 11151 35092 11237 35148
rect 11293 35092 11379 35148
rect 11435 35092 11521 35148
rect 11577 35092 11663 35148
rect 11719 35092 11805 35148
rect 11861 35092 11947 35148
rect 12003 35092 12089 35148
rect 12145 35092 12231 35148
rect 12287 35092 12373 35148
rect 12429 35092 12515 35148
rect 12571 35092 12657 35148
rect 12713 35092 12799 35148
rect 12855 35092 12941 35148
rect 12997 35092 13083 35148
rect 13139 35092 13225 35148
rect 13281 35092 13367 35148
rect 13423 35092 13509 35148
rect 13565 35092 13651 35148
rect 13707 35092 13793 35148
rect 13849 35092 13935 35148
rect 13991 35092 14077 35148
rect 14133 35092 14219 35148
rect 14275 35092 14361 35148
rect 14417 35092 14503 35148
rect 14559 35092 14645 35148
rect 14701 35092 14787 35148
rect 14843 35092 14853 35148
rect 151 35006 14853 35092
rect 151 34950 161 35006
rect 217 34950 303 35006
rect 359 34950 445 35006
rect 501 34950 587 35006
rect 643 34950 729 35006
rect 785 34950 871 35006
rect 927 34950 1013 35006
rect 1069 34950 1155 35006
rect 1211 34950 1297 35006
rect 1353 34950 1439 35006
rect 1495 34950 1581 35006
rect 1637 34950 1723 35006
rect 1779 34950 1865 35006
rect 1921 34950 2007 35006
rect 2063 34950 2149 35006
rect 2205 34950 2291 35006
rect 2347 34950 2433 35006
rect 2489 34950 2575 35006
rect 2631 34950 2717 35006
rect 2773 34950 2859 35006
rect 2915 34950 3001 35006
rect 3057 34950 3143 35006
rect 3199 34950 3285 35006
rect 3341 34950 3427 35006
rect 3483 34950 3569 35006
rect 3625 34950 3711 35006
rect 3767 34950 3853 35006
rect 3909 34950 3995 35006
rect 4051 34950 4137 35006
rect 4193 34950 4279 35006
rect 4335 34950 4421 35006
rect 4477 34950 4563 35006
rect 4619 34950 4705 35006
rect 4761 34950 4847 35006
rect 4903 34950 4989 35006
rect 5045 34950 5131 35006
rect 5187 34950 5273 35006
rect 5329 34950 5415 35006
rect 5471 34950 5557 35006
rect 5613 34950 5699 35006
rect 5755 34950 5841 35006
rect 5897 34950 5983 35006
rect 6039 34950 6125 35006
rect 6181 34950 6267 35006
rect 6323 34950 6409 35006
rect 6465 34950 6551 35006
rect 6607 34950 6693 35006
rect 6749 34950 6835 35006
rect 6891 34950 6977 35006
rect 7033 34950 7119 35006
rect 7175 34950 7261 35006
rect 7317 34950 7403 35006
rect 7459 34950 7545 35006
rect 7601 34950 7687 35006
rect 7743 34950 7829 35006
rect 7885 34950 7971 35006
rect 8027 34950 8113 35006
rect 8169 34950 8255 35006
rect 8311 34950 8397 35006
rect 8453 34950 8539 35006
rect 8595 34950 8681 35006
rect 8737 34950 8823 35006
rect 8879 34950 8965 35006
rect 9021 34950 9107 35006
rect 9163 34950 9249 35006
rect 9305 34950 9391 35006
rect 9447 34950 9533 35006
rect 9589 34950 9675 35006
rect 9731 34950 9817 35006
rect 9873 34950 9959 35006
rect 10015 34950 10101 35006
rect 10157 34950 10243 35006
rect 10299 34950 10385 35006
rect 10441 34950 10527 35006
rect 10583 34950 10669 35006
rect 10725 34950 10811 35006
rect 10867 34950 10953 35006
rect 11009 34950 11095 35006
rect 11151 34950 11237 35006
rect 11293 34950 11379 35006
rect 11435 34950 11521 35006
rect 11577 34950 11663 35006
rect 11719 34950 11805 35006
rect 11861 34950 11947 35006
rect 12003 34950 12089 35006
rect 12145 34950 12231 35006
rect 12287 34950 12373 35006
rect 12429 34950 12515 35006
rect 12571 34950 12657 35006
rect 12713 34950 12799 35006
rect 12855 34950 12941 35006
rect 12997 34950 13083 35006
rect 13139 34950 13225 35006
rect 13281 34950 13367 35006
rect 13423 34950 13509 35006
rect 13565 34950 13651 35006
rect 13707 34950 13793 35006
rect 13849 34950 13935 35006
rect 13991 34950 14077 35006
rect 14133 34950 14219 35006
rect 14275 34950 14361 35006
rect 14417 34950 14503 35006
rect 14559 34950 14645 35006
rect 14701 34950 14787 35006
rect 14843 34950 14853 35006
rect 151 34864 14853 34950
rect 151 34808 161 34864
rect 217 34808 303 34864
rect 359 34808 445 34864
rect 501 34808 587 34864
rect 643 34808 729 34864
rect 785 34808 871 34864
rect 927 34808 1013 34864
rect 1069 34808 1155 34864
rect 1211 34808 1297 34864
rect 1353 34808 1439 34864
rect 1495 34808 1581 34864
rect 1637 34808 1723 34864
rect 1779 34808 1865 34864
rect 1921 34808 2007 34864
rect 2063 34808 2149 34864
rect 2205 34808 2291 34864
rect 2347 34808 2433 34864
rect 2489 34808 2575 34864
rect 2631 34808 2717 34864
rect 2773 34808 2859 34864
rect 2915 34808 3001 34864
rect 3057 34808 3143 34864
rect 3199 34808 3285 34864
rect 3341 34808 3427 34864
rect 3483 34808 3569 34864
rect 3625 34808 3711 34864
rect 3767 34808 3853 34864
rect 3909 34808 3995 34864
rect 4051 34808 4137 34864
rect 4193 34808 4279 34864
rect 4335 34808 4421 34864
rect 4477 34808 4563 34864
rect 4619 34808 4705 34864
rect 4761 34808 4847 34864
rect 4903 34808 4989 34864
rect 5045 34808 5131 34864
rect 5187 34808 5273 34864
rect 5329 34808 5415 34864
rect 5471 34808 5557 34864
rect 5613 34808 5699 34864
rect 5755 34808 5841 34864
rect 5897 34808 5983 34864
rect 6039 34808 6125 34864
rect 6181 34808 6267 34864
rect 6323 34808 6409 34864
rect 6465 34808 6551 34864
rect 6607 34808 6693 34864
rect 6749 34808 6835 34864
rect 6891 34808 6977 34864
rect 7033 34808 7119 34864
rect 7175 34808 7261 34864
rect 7317 34808 7403 34864
rect 7459 34808 7545 34864
rect 7601 34808 7687 34864
rect 7743 34808 7829 34864
rect 7885 34808 7971 34864
rect 8027 34808 8113 34864
rect 8169 34808 8255 34864
rect 8311 34808 8397 34864
rect 8453 34808 8539 34864
rect 8595 34808 8681 34864
rect 8737 34808 8823 34864
rect 8879 34808 8965 34864
rect 9021 34808 9107 34864
rect 9163 34808 9249 34864
rect 9305 34808 9391 34864
rect 9447 34808 9533 34864
rect 9589 34808 9675 34864
rect 9731 34808 9817 34864
rect 9873 34808 9959 34864
rect 10015 34808 10101 34864
rect 10157 34808 10243 34864
rect 10299 34808 10385 34864
rect 10441 34808 10527 34864
rect 10583 34808 10669 34864
rect 10725 34808 10811 34864
rect 10867 34808 10953 34864
rect 11009 34808 11095 34864
rect 11151 34808 11237 34864
rect 11293 34808 11379 34864
rect 11435 34808 11521 34864
rect 11577 34808 11663 34864
rect 11719 34808 11805 34864
rect 11861 34808 11947 34864
rect 12003 34808 12089 34864
rect 12145 34808 12231 34864
rect 12287 34808 12373 34864
rect 12429 34808 12515 34864
rect 12571 34808 12657 34864
rect 12713 34808 12799 34864
rect 12855 34808 12941 34864
rect 12997 34808 13083 34864
rect 13139 34808 13225 34864
rect 13281 34808 13367 34864
rect 13423 34808 13509 34864
rect 13565 34808 13651 34864
rect 13707 34808 13793 34864
rect 13849 34808 13935 34864
rect 13991 34808 14077 34864
rect 14133 34808 14219 34864
rect 14275 34808 14361 34864
rect 14417 34808 14503 34864
rect 14559 34808 14645 34864
rect 14701 34808 14787 34864
rect 14843 34808 14853 34864
rect 151 34722 14853 34808
rect 151 34666 161 34722
rect 217 34666 303 34722
rect 359 34666 445 34722
rect 501 34666 587 34722
rect 643 34666 729 34722
rect 785 34666 871 34722
rect 927 34666 1013 34722
rect 1069 34666 1155 34722
rect 1211 34666 1297 34722
rect 1353 34666 1439 34722
rect 1495 34666 1581 34722
rect 1637 34666 1723 34722
rect 1779 34666 1865 34722
rect 1921 34666 2007 34722
rect 2063 34666 2149 34722
rect 2205 34666 2291 34722
rect 2347 34666 2433 34722
rect 2489 34666 2575 34722
rect 2631 34666 2717 34722
rect 2773 34666 2859 34722
rect 2915 34666 3001 34722
rect 3057 34666 3143 34722
rect 3199 34666 3285 34722
rect 3341 34666 3427 34722
rect 3483 34666 3569 34722
rect 3625 34666 3711 34722
rect 3767 34666 3853 34722
rect 3909 34666 3995 34722
rect 4051 34666 4137 34722
rect 4193 34666 4279 34722
rect 4335 34666 4421 34722
rect 4477 34666 4563 34722
rect 4619 34666 4705 34722
rect 4761 34666 4847 34722
rect 4903 34666 4989 34722
rect 5045 34666 5131 34722
rect 5187 34666 5273 34722
rect 5329 34666 5415 34722
rect 5471 34666 5557 34722
rect 5613 34666 5699 34722
rect 5755 34666 5841 34722
rect 5897 34666 5983 34722
rect 6039 34666 6125 34722
rect 6181 34666 6267 34722
rect 6323 34666 6409 34722
rect 6465 34666 6551 34722
rect 6607 34666 6693 34722
rect 6749 34666 6835 34722
rect 6891 34666 6977 34722
rect 7033 34666 7119 34722
rect 7175 34666 7261 34722
rect 7317 34666 7403 34722
rect 7459 34666 7545 34722
rect 7601 34666 7687 34722
rect 7743 34666 7829 34722
rect 7885 34666 7971 34722
rect 8027 34666 8113 34722
rect 8169 34666 8255 34722
rect 8311 34666 8397 34722
rect 8453 34666 8539 34722
rect 8595 34666 8681 34722
rect 8737 34666 8823 34722
rect 8879 34666 8965 34722
rect 9021 34666 9107 34722
rect 9163 34666 9249 34722
rect 9305 34666 9391 34722
rect 9447 34666 9533 34722
rect 9589 34666 9675 34722
rect 9731 34666 9817 34722
rect 9873 34666 9959 34722
rect 10015 34666 10101 34722
rect 10157 34666 10243 34722
rect 10299 34666 10385 34722
rect 10441 34666 10527 34722
rect 10583 34666 10669 34722
rect 10725 34666 10811 34722
rect 10867 34666 10953 34722
rect 11009 34666 11095 34722
rect 11151 34666 11237 34722
rect 11293 34666 11379 34722
rect 11435 34666 11521 34722
rect 11577 34666 11663 34722
rect 11719 34666 11805 34722
rect 11861 34666 11947 34722
rect 12003 34666 12089 34722
rect 12145 34666 12231 34722
rect 12287 34666 12373 34722
rect 12429 34666 12515 34722
rect 12571 34666 12657 34722
rect 12713 34666 12799 34722
rect 12855 34666 12941 34722
rect 12997 34666 13083 34722
rect 13139 34666 13225 34722
rect 13281 34666 13367 34722
rect 13423 34666 13509 34722
rect 13565 34666 13651 34722
rect 13707 34666 13793 34722
rect 13849 34666 13935 34722
rect 13991 34666 14077 34722
rect 14133 34666 14219 34722
rect 14275 34666 14361 34722
rect 14417 34666 14503 34722
rect 14559 34666 14645 34722
rect 14701 34666 14787 34722
rect 14843 34666 14853 34722
rect 151 34580 14853 34666
rect 151 34524 161 34580
rect 217 34524 303 34580
rect 359 34524 445 34580
rect 501 34524 587 34580
rect 643 34524 729 34580
rect 785 34524 871 34580
rect 927 34524 1013 34580
rect 1069 34524 1155 34580
rect 1211 34524 1297 34580
rect 1353 34524 1439 34580
rect 1495 34524 1581 34580
rect 1637 34524 1723 34580
rect 1779 34524 1865 34580
rect 1921 34524 2007 34580
rect 2063 34524 2149 34580
rect 2205 34524 2291 34580
rect 2347 34524 2433 34580
rect 2489 34524 2575 34580
rect 2631 34524 2717 34580
rect 2773 34524 2859 34580
rect 2915 34524 3001 34580
rect 3057 34524 3143 34580
rect 3199 34524 3285 34580
rect 3341 34524 3427 34580
rect 3483 34524 3569 34580
rect 3625 34524 3711 34580
rect 3767 34524 3853 34580
rect 3909 34524 3995 34580
rect 4051 34524 4137 34580
rect 4193 34524 4279 34580
rect 4335 34524 4421 34580
rect 4477 34524 4563 34580
rect 4619 34524 4705 34580
rect 4761 34524 4847 34580
rect 4903 34524 4989 34580
rect 5045 34524 5131 34580
rect 5187 34524 5273 34580
rect 5329 34524 5415 34580
rect 5471 34524 5557 34580
rect 5613 34524 5699 34580
rect 5755 34524 5841 34580
rect 5897 34524 5983 34580
rect 6039 34524 6125 34580
rect 6181 34524 6267 34580
rect 6323 34524 6409 34580
rect 6465 34524 6551 34580
rect 6607 34524 6693 34580
rect 6749 34524 6835 34580
rect 6891 34524 6977 34580
rect 7033 34524 7119 34580
rect 7175 34524 7261 34580
rect 7317 34524 7403 34580
rect 7459 34524 7545 34580
rect 7601 34524 7687 34580
rect 7743 34524 7829 34580
rect 7885 34524 7971 34580
rect 8027 34524 8113 34580
rect 8169 34524 8255 34580
rect 8311 34524 8397 34580
rect 8453 34524 8539 34580
rect 8595 34524 8681 34580
rect 8737 34524 8823 34580
rect 8879 34524 8965 34580
rect 9021 34524 9107 34580
rect 9163 34524 9249 34580
rect 9305 34524 9391 34580
rect 9447 34524 9533 34580
rect 9589 34524 9675 34580
rect 9731 34524 9817 34580
rect 9873 34524 9959 34580
rect 10015 34524 10101 34580
rect 10157 34524 10243 34580
rect 10299 34524 10385 34580
rect 10441 34524 10527 34580
rect 10583 34524 10669 34580
rect 10725 34524 10811 34580
rect 10867 34524 10953 34580
rect 11009 34524 11095 34580
rect 11151 34524 11237 34580
rect 11293 34524 11379 34580
rect 11435 34524 11521 34580
rect 11577 34524 11663 34580
rect 11719 34524 11805 34580
rect 11861 34524 11947 34580
rect 12003 34524 12089 34580
rect 12145 34524 12231 34580
rect 12287 34524 12373 34580
rect 12429 34524 12515 34580
rect 12571 34524 12657 34580
rect 12713 34524 12799 34580
rect 12855 34524 12941 34580
rect 12997 34524 13083 34580
rect 13139 34524 13225 34580
rect 13281 34524 13367 34580
rect 13423 34524 13509 34580
rect 13565 34524 13651 34580
rect 13707 34524 13793 34580
rect 13849 34524 13935 34580
rect 13991 34524 14077 34580
rect 14133 34524 14219 34580
rect 14275 34524 14361 34580
rect 14417 34524 14503 34580
rect 14559 34524 14645 34580
rect 14701 34524 14787 34580
rect 14843 34524 14853 34580
rect 151 34438 14853 34524
rect 151 34382 161 34438
rect 217 34382 303 34438
rect 359 34382 445 34438
rect 501 34382 587 34438
rect 643 34382 729 34438
rect 785 34382 871 34438
rect 927 34382 1013 34438
rect 1069 34382 1155 34438
rect 1211 34382 1297 34438
rect 1353 34382 1439 34438
rect 1495 34382 1581 34438
rect 1637 34382 1723 34438
rect 1779 34382 1865 34438
rect 1921 34382 2007 34438
rect 2063 34382 2149 34438
rect 2205 34382 2291 34438
rect 2347 34382 2433 34438
rect 2489 34382 2575 34438
rect 2631 34382 2717 34438
rect 2773 34382 2859 34438
rect 2915 34382 3001 34438
rect 3057 34382 3143 34438
rect 3199 34382 3285 34438
rect 3341 34382 3427 34438
rect 3483 34382 3569 34438
rect 3625 34382 3711 34438
rect 3767 34382 3853 34438
rect 3909 34382 3995 34438
rect 4051 34382 4137 34438
rect 4193 34382 4279 34438
rect 4335 34382 4421 34438
rect 4477 34382 4563 34438
rect 4619 34382 4705 34438
rect 4761 34382 4847 34438
rect 4903 34382 4989 34438
rect 5045 34382 5131 34438
rect 5187 34382 5273 34438
rect 5329 34382 5415 34438
rect 5471 34382 5557 34438
rect 5613 34382 5699 34438
rect 5755 34382 5841 34438
rect 5897 34382 5983 34438
rect 6039 34382 6125 34438
rect 6181 34382 6267 34438
rect 6323 34382 6409 34438
rect 6465 34382 6551 34438
rect 6607 34382 6693 34438
rect 6749 34382 6835 34438
rect 6891 34382 6977 34438
rect 7033 34382 7119 34438
rect 7175 34382 7261 34438
rect 7317 34382 7403 34438
rect 7459 34382 7545 34438
rect 7601 34382 7687 34438
rect 7743 34382 7829 34438
rect 7885 34382 7971 34438
rect 8027 34382 8113 34438
rect 8169 34382 8255 34438
rect 8311 34382 8397 34438
rect 8453 34382 8539 34438
rect 8595 34382 8681 34438
rect 8737 34382 8823 34438
rect 8879 34382 8965 34438
rect 9021 34382 9107 34438
rect 9163 34382 9249 34438
rect 9305 34382 9391 34438
rect 9447 34382 9533 34438
rect 9589 34382 9675 34438
rect 9731 34382 9817 34438
rect 9873 34382 9959 34438
rect 10015 34382 10101 34438
rect 10157 34382 10243 34438
rect 10299 34382 10385 34438
rect 10441 34382 10527 34438
rect 10583 34382 10669 34438
rect 10725 34382 10811 34438
rect 10867 34382 10953 34438
rect 11009 34382 11095 34438
rect 11151 34382 11237 34438
rect 11293 34382 11379 34438
rect 11435 34382 11521 34438
rect 11577 34382 11663 34438
rect 11719 34382 11805 34438
rect 11861 34382 11947 34438
rect 12003 34382 12089 34438
rect 12145 34382 12231 34438
rect 12287 34382 12373 34438
rect 12429 34382 12515 34438
rect 12571 34382 12657 34438
rect 12713 34382 12799 34438
rect 12855 34382 12941 34438
rect 12997 34382 13083 34438
rect 13139 34382 13225 34438
rect 13281 34382 13367 34438
rect 13423 34382 13509 34438
rect 13565 34382 13651 34438
rect 13707 34382 13793 34438
rect 13849 34382 13935 34438
rect 13991 34382 14077 34438
rect 14133 34382 14219 34438
rect 14275 34382 14361 34438
rect 14417 34382 14503 34438
rect 14559 34382 14645 34438
rect 14701 34382 14787 34438
rect 14843 34382 14853 34438
rect 151 34296 14853 34382
rect 151 34240 161 34296
rect 217 34240 303 34296
rect 359 34240 445 34296
rect 501 34240 587 34296
rect 643 34240 729 34296
rect 785 34240 871 34296
rect 927 34240 1013 34296
rect 1069 34240 1155 34296
rect 1211 34240 1297 34296
rect 1353 34240 1439 34296
rect 1495 34240 1581 34296
rect 1637 34240 1723 34296
rect 1779 34240 1865 34296
rect 1921 34240 2007 34296
rect 2063 34240 2149 34296
rect 2205 34240 2291 34296
rect 2347 34240 2433 34296
rect 2489 34240 2575 34296
rect 2631 34240 2717 34296
rect 2773 34240 2859 34296
rect 2915 34240 3001 34296
rect 3057 34240 3143 34296
rect 3199 34240 3285 34296
rect 3341 34240 3427 34296
rect 3483 34240 3569 34296
rect 3625 34240 3711 34296
rect 3767 34240 3853 34296
rect 3909 34240 3995 34296
rect 4051 34240 4137 34296
rect 4193 34240 4279 34296
rect 4335 34240 4421 34296
rect 4477 34240 4563 34296
rect 4619 34240 4705 34296
rect 4761 34240 4847 34296
rect 4903 34240 4989 34296
rect 5045 34240 5131 34296
rect 5187 34240 5273 34296
rect 5329 34240 5415 34296
rect 5471 34240 5557 34296
rect 5613 34240 5699 34296
rect 5755 34240 5841 34296
rect 5897 34240 5983 34296
rect 6039 34240 6125 34296
rect 6181 34240 6267 34296
rect 6323 34240 6409 34296
rect 6465 34240 6551 34296
rect 6607 34240 6693 34296
rect 6749 34240 6835 34296
rect 6891 34240 6977 34296
rect 7033 34240 7119 34296
rect 7175 34240 7261 34296
rect 7317 34240 7403 34296
rect 7459 34240 7545 34296
rect 7601 34240 7687 34296
rect 7743 34240 7829 34296
rect 7885 34240 7971 34296
rect 8027 34240 8113 34296
rect 8169 34240 8255 34296
rect 8311 34240 8397 34296
rect 8453 34240 8539 34296
rect 8595 34240 8681 34296
rect 8737 34240 8823 34296
rect 8879 34240 8965 34296
rect 9021 34240 9107 34296
rect 9163 34240 9249 34296
rect 9305 34240 9391 34296
rect 9447 34240 9533 34296
rect 9589 34240 9675 34296
rect 9731 34240 9817 34296
rect 9873 34240 9959 34296
rect 10015 34240 10101 34296
rect 10157 34240 10243 34296
rect 10299 34240 10385 34296
rect 10441 34240 10527 34296
rect 10583 34240 10669 34296
rect 10725 34240 10811 34296
rect 10867 34240 10953 34296
rect 11009 34240 11095 34296
rect 11151 34240 11237 34296
rect 11293 34240 11379 34296
rect 11435 34240 11521 34296
rect 11577 34240 11663 34296
rect 11719 34240 11805 34296
rect 11861 34240 11947 34296
rect 12003 34240 12089 34296
rect 12145 34240 12231 34296
rect 12287 34240 12373 34296
rect 12429 34240 12515 34296
rect 12571 34240 12657 34296
rect 12713 34240 12799 34296
rect 12855 34240 12941 34296
rect 12997 34240 13083 34296
rect 13139 34240 13225 34296
rect 13281 34240 13367 34296
rect 13423 34240 13509 34296
rect 13565 34240 13651 34296
rect 13707 34240 13793 34296
rect 13849 34240 13935 34296
rect 13991 34240 14077 34296
rect 14133 34240 14219 34296
rect 14275 34240 14361 34296
rect 14417 34240 14503 34296
rect 14559 34240 14645 34296
rect 14701 34240 14787 34296
rect 14843 34240 14853 34296
rect 151 34154 14853 34240
rect 151 34098 161 34154
rect 217 34098 303 34154
rect 359 34098 445 34154
rect 501 34098 587 34154
rect 643 34098 729 34154
rect 785 34098 871 34154
rect 927 34098 1013 34154
rect 1069 34098 1155 34154
rect 1211 34098 1297 34154
rect 1353 34098 1439 34154
rect 1495 34098 1581 34154
rect 1637 34098 1723 34154
rect 1779 34098 1865 34154
rect 1921 34098 2007 34154
rect 2063 34098 2149 34154
rect 2205 34098 2291 34154
rect 2347 34098 2433 34154
rect 2489 34098 2575 34154
rect 2631 34098 2717 34154
rect 2773 34098 2859 34154
rect 2915 34098 3001 34154
rect 3057 34098 3143 34154
rect 3199 34098 3285 34154
rect 3341 34098 3427 34154
rect 3483 34098 3569 34154
rect 3625 34098 3711 34154
rect 3767 34098 3853 34154
rect 3909 34098 3995 34154
rect 4051 34098 4137 34154
rect 4193 34098 4279 34154
rect 4335 34098 4421 34154
rect 4477 34098 4563 34154
rect 4619 34098 4705 34154
rect 4761 34098 4847 34154
rect 4903 34098 4989 34154
rect 5045 34098 5131 34154
rect 5187 34098 5273 34154
rect 5329 34098 5415 34154
rect 5471 34098 5557 34154
rect 5613 34098 5699 34154
rect 5755 34098 5841 34154
rect 5897 34098 5983 34154
rect 6039 34098 6125 34154
rect 6181 34098 6267 34154
rect 6323 34098 6409 34154
rect 6465 34098 6551 34154
rect 6607 34098 6693 34154
rect 6749 34098 6835 34154
rect 6891 34098 6977 34154
rect 7033 34098 7119 34154
rect 7175 34098 7261 34154
rect 7317 34098 7403 34154
rect 7459 34098 7545 34154
rect 7601 34098 7687 34154
rect 7743 34098 7829 34154
rect 7885 34098 7971 34154
rect 8027 34098 8113 34154
rect 8169 34098 8255 34154
rect 8311 34098 8397 34154
rect 8453 34098 8539 34154
rect 8595 34098 8681 34154
rect 8737 34098 8823 34154
rect 8879 34098 8965 34154
rect 9021 34098 9107 34154
rect 9163 34098 9249 34154
rect 9305 34098 9391 34154
rect 9447 34098 9533 34154
rect 9589 34098 9675 34154
rect 9731 34098 9817 34154
rect 9873 34098 9959 34154
rect 10015 34098 10101 34154
rect 10157 34098 10243 34154
rect 10299 34098 10385 34154
rect 10441 34098 10527 34154
rect 10583 34098 10669 34154
rect 10725 34098 10811 34154
rect 10867 34098 10953 34154
rect 11009 34098 11095 34154
rect 11151 34098 11237 34154
rect 11293 34098 11379 34154
rect 11435 34098 11521 34154
rect 11577 34098 11663 34154
rect 11719 34098 11805 34154
rect 11861 34098 11947 34154
rect 12003 34098 12089 34154
rect 12145 34098 12231 34154
rect 12287 34098 12373 34154
rect 12429 34098 12515 34154
rect 12571 34098 12657 34154
rect 12713 34098 12799 34154
rect 12855 34098 12941 34154
rect 12997 34098 13083 34154
rect 13139 34098 13225 34154
rect 13281 34098 13367 34154
rect 13423 34098 13509 34154
rect 13565 34098 13651 34154
rect 13707 34098 13793 34154
rect 13849 34098 13935 34154
rect 13991 34098 14077 34154
rect 14133 34098 14219 34154
rect 14275 34098 14361 34154
rect 14417 34098 14503 34154
rect 14559 34098 14645 34154
rect 14701 34098 14787 34154
rect 14843 34098 14853 34154
rect 151 34012 14853 34098
rect 151 33956 161 34012
rect 217 33956 303 34012
rect 359 33956 445 34012
rect 501 33956 587 34012
rect 643 33956 729 34012
rect 785 33956 871 34012
rect 927 33956 1013 34012
rect 1069 33956 1155 34012
rect 1211 33956 1297 34012
rect 1353 33956 1439 34012
rect 1495 33956 1581 34012
rect 1637 33956 1723 34012
rect 1779 33956 1865 34012
rect 1921 33956 2007 34012
rect 2063 33956 2149 34012
rect 2205 33956 2291 34012
rect 2347 33956 2433 34012
rect 2489 33956 2575 34012
rect 2631 33956 2717 34012
rect 2773 33956 2859 34012
rect 2915 33956 3001 34012
rect 3057 33956 3143 34012
rect 3199 33956 3285 34012
rect 3341 33956 3427 34012
rect 3483 33956 3569 34012
rect 3625 33956 3711 34012
rect 3767 33956 3853 34012
rect 3909 33956 3995 34012
rect 4051 33956 4137 34012
rect 4193 33956 4279 34012
rect 4335 33956 4421 34012
rect 4477 33956 4563 34012
rect 4619 33956 4705 34012
rect 4761 33956 4847 34012
rect 4903 33956 4989 34012
rect 5045 33956 5131 34012
rect 5187 33956 5273 34012
rect 5329 33956 5415 34012
rect 5471 33956 5557 34012
rect 5613 33956 5699 34012
rect 5755 33956 5841 34012
rect 5897 33956 5983 34012
rect 6039 33956 6125 34012
rect 6181 33956 6267 34012
rect 6323 33956 6409 34012
rect 6465 33956 6551 34012
rect 6607 33956 6693 34012
rect 6749 33956 6835 34012
rect 6891 33956 6977 34012
rect 7033 33956 7119 34012
rect 7175 33956 7261 34012
rect 7317 33956 7403 34012
rect 7459 33956 7545 34012
rect 7601 33956 7687 34012
rect 7743 33956 7829 34012
rect 7885 33956 7971 34012
rect 8027 33956 8113 34012
rect 8169 33956 8255 34012
rect 8311 33956 8397 34012
rect 8453 33956 8539 34012
rect 8595 33956 8681 34012
rect 8737 33956 8823 34012
rect 8879 33956 8965 34012
rect 9021 33956 9107 34012
rect 9163 33956 9249 34012
rect 9305 33956 9391 34012
rect 9447 33956 9533 34012
rect 9589 33956 9675 34012
rect 9731 33956 9817 34012
rect 9873 33956 9959 34012
rect 10015 33956 10101 34012
rect 10157 33956 10243 34012
rect 10299 33956 10385 34012
rect 10441 33956 10527 34012
rect 10583 33956 10669 34012
rect 10725 33956 10811 34012
rect 10867 33956 10953 34012
rect 11009 33956 11095 34012
rect 11151 33956 11237 34012
rect 11293 33956 11379 34012
rect 11435 33956 11521 34012
rect 11577 33956 11663 34012
rect 11719 33956 11805 34012
rect 11861 33956 11947 34012
rect 12003 33956 12089 34012
rect 12145 33956 12231 34012
rect 12287 33956 12373 34012
rect 12429 33956 12515 34012
rect 12571 33956 12657 34012
rect 12713 33956 12799 34012
rect 12855 33956 12941 34012
rect 12997 33956 13083 34012
rect 13139 33956 13225 34012
rect 13281 33956 13367 34012
rect 13423 33956 13509 34012
rect 13565 33956 13651 34012
rect 13707 33956 13793 34012
rect 13849 33956 13935 34012
rect 13991 33956 14077 34012
rect 14133 33956 14219 34012
rect 14275 33956 14361 34012
rect 14417 33956 14503 34012
rect 14559 33956 14645 34012
rect 14701 33956 14787 34012
rect 14843 33956 14853 34012
rect 151 33870 14853 33956
rect 151 33814 161 33870
rect 217 33814 303 33870
rect 359 33814 445 33870
rect 501 33814 587 33870
rect 643 33814 729 33870
rect 785 33814 871 33870
rect 927 33814 1013 33870
rect 1069 33814 1155 33870
rect 1211 33814 1297 33870
rect 1353 33814 1439 33870
rect 1495 33814 1581 33870
rect 1637 33814 1723 33870
rect 1779 33814 1865 33870
rect 1921 33814 2007 33870
rect 2063 33814 2149 33870
rect 2205 33814 2291 33870
rect 2347 33814 2433 33870
rect 2489 33814 2575 33870
rect 2631 33814 2717 33870
rect 2773 33814 2859 33870
rect 2915 33814 3001 33870
rect 3057 33814 3143 33870
rect 3199 33814 3285 33870
rect 3341 33814 3427 33870
rect 3483 33814 3569 33870
rect 3625 33814 3711 33870
rect 3767 33814 3853 33870
rect 3909 33814 3995 33870
rect 4051 33814 4137 33870
rect 4193 33814 4279 33870
rect 4335 33814 4421 33870
rect 4477 33814 4563 33870
rect 4619 33814 4705 33870
rect 4761 33814 4847 33870
rect 4903 33814 4989 33870
rect 5045 33814 5131 33870
rect 5187 33814 5273 33870
rect 5329 33814 5415 33870
rect 5471 33814 5557 33870
rect 5613 33814 5699 33870
rect 5755 33814 5841 33870
rect 5897 33814 5983 33870
rect 6039 33814 6125 33870
rect 6181 33814 6267 33870
rect 6323 33814 6409 33870
rect 6465 33814 6551 33870
rect 6607 33814 6693 33870
rect 6749 33814 6835 33870
rect 6891 33814 6977 33870
rect 7033 33814 7119 33870
rect 7175 33814 7261 33870
rect 7317 33814 7403 33870
rect 7459 33814 7545 33870
rect 7601 33814 7687 33870
rect 7743 33814 7829 33870
rect 7885 33814 7971 33870
rect 8027 33814 8113 33870
rect 8169 33814 8255 33870
rect 8311 33814 8397 33870
rect 8453 33814 8539 33870
rect 8595 33814 8681 33870
rect 8737 33814 8823 33870
rect 8879 33814 8965 33870
rect 9021 33814 9107 33870
rect 9163 33814 9249 33870
rect 9305 33814 9391 33870
rect 9447 33814 9533 33870
rect 9589 33814 9675 33870
rect 9731 33814 9817 33870
rect 9873 33814 9959 33870
rect 10015 33814 10101 33870
rect 10157 33814 10243 33870
rect 10299 33814 10385 33870
rect 10441 33814 10527 33870
rect 10583 33814 10669 33870
rect 10725 33814 10811 33870
rect 10867 33814 10953 33870
rect 11009 33814 11095 33870
rect 11151 33814 11237 33870
rect 11293 33814 11379 33870
rect 11435 33814 11521 33870
rect 11577 33814 11663 33870
rect 11719 33814 11805 33870
rect 11861 33814 11947 33870
rect 12003 33814 12089 33870
rect 12145 33814 12231 33870
rect 12287 33814 12373 33870
rect 12429 33814 12515 33870
rect 12571 33814 12657 33870
rect 12713 33814 12799 33870
rect 12855 33814 12941 33870
rect 12997 33814 13083 33870
rect 13139 33814 13225 33870
rect 13281 33814 13367 33870
rect 13423 33814 13509 33870
rect 13565 33814 13651 33870
rect 13707 33814 13793 33870
rect 13849 33814 13935 33870
rect 13991 33814 14077 33870
rect 14133 33814 14219 33870
rect 14275 33814 14361 33870
rect 14417 33814 14503 33870
rect 14559 33814 14645 33870
rect 14701 33814 14787 33870
rect 14843 33814 14853 33870
rect 151 33728 14853 33814
rect 151 33672 161 33728
rect 217 33672 303 33728
rect 359 33672 445 33728
rect 501 33672 587 33728
rect 643 33672 729 33728
rect 785 33672 871 33728
rect 927 33672 1013 33728
rect 1069 33672 1155 33728
rect 1211 33672 1297 33728
rect 1353 33672 1439 33728
rect 1495 33672 1581 33728
rect 1637 33672 1723 33728
rect 1779 33672 1865 33728
rect 1921 33672 2007 33728
rect 2063 33672 2149 33728
rect 2205 33672 2291 33728
rect 2347 33672 2433 33728
rect 2489 33672 2575 33728
rect 2631 33672 2717 33728
rect 2773 33672 2859 33728
rect 2915 33672 3001 33728
rect 3057 33672 3143 33728
rect 3199 33672 3285 33728
rect 3341 33672 3427 33728
rect 3483 33672 3569 33728
rect 3625 33672 3711 33728
rect 3767 33672 3853 33728
rect 3909 33672 3995 33728
rect 4051 33672 4137 33728
rect 4193 33672 4279 33728
rect 4335 33672 4421 33728
rect 4477 33672 4563 33728
rect 4619 33672 4705 33728
rect 4761 33672 4847 33728
rect 4903 33672 4989 33728
rect 5045 33672 5131 33728
rect 5187 33672 5273 33728
rect 5329 33672 5415 33728
rect 5471 33672 5557 33728
rect 5613 33672 5699 33728
rect 5755 33672 5841 33728
rect 5897 33672 5983 33728
rect 6039 33672 6125 33728
rect 6181 33672 6267 33728
rect 6323 33672 6409 33728
rect 6465 33672 6551 33728
rect 6607 33672 6693 33728
rect 6749 33672 6835 33728
rect 6891 33672 6977 33728
rect 7033 33672 7119 33728
rect 7175 33672 7261 33728
rect 7317 33672 7403 33728
rect 7459 33672 7545 33728
rect 7601 33672 7687 33728
rect 7743 33672 7829 33728
rect 7885 33672 7971 33728
rect 8027 33672 8113 33728
rect 8169 33672 8255 33728
rect 8311 33672 8397 33728
rect 8453 33672 8539 33728
rect 8595 33672 8681 33728
rect 8737 33672 8823 33728
rect 8879 33672 8965 33728
rect 9021 33672 9107 33728
rect 9163 33672 9249 33728
rect 9305 33672 9391 33728
rect 9447 33672 9533 33728
rect 9589 33672 9675 33728
rect 9731 33672 9817 33728
rect 9873 33672 9959 33728
rect 10015 33672 10101 33728
rect 10157 33672 10243 33728
rect 10299 33672 10385 33728
rect 10441 33672 10527 33728
rect 10583 33672 10669 33728
rect 10725 33672 10811 33728
rect 10867 33672 10953 33728
rect 11009 33672 11095 33728
rect 11151 33672 11237 33728
rect 11293 33672 11379 33728
rect 11435 33672 11521 33728
rect 11577 33672 11663 33728
rect 11719 33672 11805 33728
rect 11861 33672 11947 33728
rect 12003 33672 12089 33728
rect 12145 33672 12231 33728
rect 12287 33672 12373 33728
rect 12429 33672 12515 33728
rect 12571 33672 12657 33728
rect 12713 33672 12799 33728
rect 12855 33672 12941 33728
rect 12997 33672 13083 33728
rect 13139 33672 13225 33728
rect 13281 33672 13367 33728
rect 13423 33672 13509 33728
rect 13565 33672 13651 33728
rect 13707 33672 13793 33728
rect 13849 33672 13935 33728
rect 13991 33672 14077 33728
rect 14133 33672 14219 33728
rect 14275 33672 14361 33728
rect 14417 33672 14503 33728
rect 14559 33672 14645 33728
rect 14701 33672 14787 33728
rect 14843 33672 14853 33728
rect 151 33586 14853 33672
rect 151 33530 161 33586
rect 217 33530 303 33586
rect 359 33530 445 33586
rect 501 33530 587 33586
rect 643 33530 729 33586
rect 785 33530 871 33586
rect 927 33530 1013 33586
rect 1069 33530 1155 33586
rect 1211 33530 1297 33586
rect 1353 33530 1439 33586
rect 1495 33530 1581 33586
rect 1637 33530 1723 33586
rect 1779 33530 1865 33586
rect 1921 33530 2007 33586
rect 2063 33530 2149 33586
rect 2205 33530 2291 33586
rect 2347 33530 2433 33586
rect 2489 33530 2575 33586
rect 2631 33530 2717 33586
rect 2773 33530 2859 33586
rect 2915 33530 3001 33586
rect 3057 33530 3143 33586
rect 3199 33530 3285 33586
rect 3341 33530 3427 33586
rect 3483 33530 3569 33586
rect 3625 33530 3711 33586
rect 3767 33530 3853 33586
rect 3909 33530 3995 33586
rect 4051 33530 4137 33586
rect 4193 33530 4279 33586
rect 4335 33530 4421 33586
rect 4477 33530 4563 33586
rect 4619 33530 4705 33586
rect 4761 33530 4847 33586
rect 4903 33530 4989 33586
rect 5045 33530 5131 33586
rect 5187 33530 5273 33586
rect 5329 33530 5415 33586
rect 5471 33530 5557 33586
rect 5613 33530 5699 33586
rect 5755 33530 5841 33586
rect 5897 33530 5983 33586
rect 6039 33530 6125 33586
rect 6181 33530 6267 33586
rect 6323 33530 6409 33586
rect 6465 33530 6551 33586
rect 6607 33530 6693 33586
rect 6749 33530 6835 33586
rect 6891 33530 6977 33586
rect 7033 33530 7119 33586
rect 7175 33530 7261 33586
rect 7317 33530 7403 33586
rect 7459 33530 7545 33586
rect 7601 33530 7687 33586
rect 7743 33530 7829 33586
rect 7885 33530 7971 33586
rect 8027 33530 8113 33586
rect 8169 33530 8255 33586
rect 8311 33530 8397 33586
rect 8453 33530 8539 33586
rect 8595 33530 8681 33586
rect 8737 33530 8823 33586
rect 8879 33530 8965 33586
rect 9021 33530 9107 33586
rect 9163 33530 9249 33586
rect 9305 33530 9391 33586
rect 9447 33530 9533 33586
rect 9589 33530 9675 33586
rect 9731 33530 9817 33586
rect 9873 33530 9959 33586
rect 10015 33530 10101 33586
rect 10157 33530 10243 33586
rect 10299 33530 10385 33586
rect 10441 33530 10527 33586
rect 10583 33530 10669 33586
rect 10725 33530 10811 33586
rect 10867 33530 10953 33586
rect 11009 33530 11095 33586
rect 11151 33530 11237 33586
rect 11293 33530 11379 33586
rect 11435 33530 11521 33586
rect 11577 33530 11663 33586
rect 11719 33530 11805 33586
rect 11861 33530 11947 33586
rect 12003 33530 12089 33586
rect 12145 33530 12231 33586
rect 12287 33530 12373 33586
rect 12429 33530 12515 33586
rect 12571 33530 12657 33586
rect 12713 33530 12799 33586
rect 12855 33530 12941 33586
rect 12997 33530 13083 33586
rect 13139 33530 13225 33586
rect 13281 33530 13367 33586
rect 13423 33530 13509 33586
rect 13565 33530 13651 33586
rect 13707 33530 13793 33586
rect 13849 33530 13935 33586
rect 13991 33530 14077 33586
rect 14133 33530 14219 33586
rect 14275 33530 14361 33586
rect 14417 33530 14503 33586
rect 14559 33530 14645 33586
rect 14701 33530 14787 33586
rect 14843 33530 14853 33586
rect 151 33444 14853 33530
rect 151 33388 161 33444
rect 217 33388 303 33444
rect 359 33388 445 33444
rect 501 33388 587 33444
rect 643 33388 729 33444
rect 785 33388 871 33444
rect 927 33388 1013 33444
rect 1069 33388 1155 33444
rect 1211 33388 1297 33444
rect 1353 33388 1439 33444
rect 1495 33388 1581 33444
rect 1637 33388 1723 33444
rect 1779 33388 1865 33444
rect 1921 33388 2007 33444
rect 2063 33388 2149 33444
rect 2205 33388 2291 33444
rect 2347 33388 2433 33444
rect 2489 33388 2575 33444
rect 2631 33388 2717 33444
rect 2773 33388 2859 33444
rect 2915 33388 3001 33444
rect 3057 33388 3143 33444
rect 3199 33388 3285 33444
rect 3341 33388 3427 33444
rect 3483 33388 3569 33444
rect 3625 33388 3711 33444
rect 3767 33388 3853 33444
rect 3909 33388 3995 33444
rect 4051 33388 4137 33444
rect 4193 33388 4279 33444
rect 4335 33388 4421 33444
rect 4477 33388 4563 33444
rect 4619 33388 4705 33444
rect 4761 33388 4847 33444
rect 4903 33388 4989 33444
rect 5045 33388 5131 33444
rect 5187 33388 5273 33444
rect 5329 33388 5415 33444
rect 5471 33388 5557 33444
rect 5613 33388 5699 33444
rect 5755 33388 5841 33444
rect 5897 33388 5983 33444
rect 6039 33388 6125 33444
rect 6181 33388 6267 33444
rect 6323 33388 6409 33444
rect 6465 33388 6551 33444
rect 6607 33388 6693 33444
rect 6749 33388 6835 33444
rect 6891 33388 6977 33444
rect 7033 33388 7119 33444
rect 7175 33388 7261 33444
rect 7317 33388 7403 33444
rect 7459 33388 7545 33444
rect 7601 33388 7687 33444
rect 7743 33388 7829 33444
rect 7885 33388 7971 33444
rect 8027 33388 8113 33444
rect 8169 33388 8255 33444
rect 8311 33388 8397 33444
rect 8453 33388 8539 33444
rect 8595 33388 8681 33444
rect 8737 33388 8823 33444
rect 8879 33388 8965 33444
rect 9021 33388 9107 33444
rect 9163 33388 9249 33444
rect 9305 33388 9391 33444
rect 9447 33388 9533 33444
rect 9589 33388 9675 33444
rect 9731 33388 9817 33444
rect 9873 33388 9959 33444
rect 10015 33388 10101 33444
rect 10157 33388 10243 33444
rect 10299 33388 10385 33444
rect 10441 33388 10527 33444
rect 10583 33388 10669 33444
rect 10725 33388 10811 33444
rect 10867 33388 10953 33444
rect 11009 33388 11095 33444
rect 11151 33388 11237 33444
rect 11293 33388 11379 33444
rect 11435 33388 11521 33444
rect 11577 33388 11663 33444
rect 11719 33388 11805 33444
rect 11861 33388 11947 33444
rect 12003 33388 12089 33444
rect 12145 33388 12231 33444
rect 12287 33388 12373 33444
rect 12429 33388 12515 33444
rect 12571 33388 12657 33444
rect 12713 33388 12799 33444
rect 12855 33388 12941 33444
rect 12997 33388 13083 33444
rect 13139 33388 13225 33444
rect 13281 33388 13367 33444
rect 13423 33388 13509 33444
rect 13565 33388 13651 33444
rect 13707 33388 13793 33444
rect 13849 33388 13935 33444
rect 13991 33388 14077 33444
rect 14133 33388 14219 33444
rect 14275 33388 14361 33444
rect 14417 33388 14503 33444
rect 14559 33388 14645 33444
rect 14701 33388 14787 33444
rect 14843 33388 14853 33444
rect 151 33302 14853 33388
rect 151 33246 161 33302
rect 217 33246 303 33302
rect 359 33246 445 33302
rect 501 33246 587 33302
rect 643 33246 729 33302
rect 785 33246 871 33302
rect 927 33246 1013 33302
rect 1069 33246 1155 33302
rect 1211 33246 1297 33302
rect 1353 33246 1439 33302
rect 1495 33246 1581 33302
rect 1637 33246 1723 33302
rect 1779 33246 1865 33302
rect 1921 33246 2007 33302
rect 2063 33246 2149 33302
rect 2205 33246 2291 33302
rect 2347 33246 2433 33302
rect 2489 33246 2575 33302
rect 2631 33246 2717 33302
rect 2773 33246 2859 33302
rect 2915 33246 3001 33302
rect 3057 33246 3143 33302
rect 3199 33246 3285 33302
rect 3341 33246 3427 33302
rect 3483 33246 3569 33302
rect 3625 33246 3711 33302
rect 3767 33246 3853 33302
rect 3909 33246 3995 33302
rect 4051 33246 4137 33302
rect 4193 33246 4279 33302
rect 4335 33246 4421 33302
rect 4477 33246 4563 33302
rect 4619 33246 4705 33302
rect 4761 33246 4847 33302
rect 4903 33246 4989 33302
rect 5045 33246 5131 33302
rect 5187 33246 5273 33302
rect 5329 33246 5415 33302
rect 5471 33246 5557 33302
rect 5613 33246 5699 33302
rect 5755 33246 5841 33302
rect 5897 33246 5983 33302
rect 6039 33246 6125 33302
rect 6181 33246 6267 33302
rect 6323 33246 6409 33302
rect 6465 33246 6551 33302
rect 6607 33246 6693 33302
rect 6749 33246 6835 33302
rect 6891 33246 6977 33302
rect 7033 33246 7119 33302
rect 7175 33246 7261 33302
rect 7317 33246 7403 33302
rect 7459 33246 7545 33302
rect 7601 33246 7687 33302
rect 7743 33246 7829 33302
rect 7885 33246 7971 33302
rect 8027 33246 8113 33302
rect 8169 33246 8255 33302
rect 8311 33246 8397 33302
rect 8453 33246 8539 33302
rect 8595 33246 8681 33302
rect 8737 33246 8823 33302
rect 8879 33246 8965 33302
rect 9021 33246 9107 33302
rect 9163 33246 9249 33302
rect 9305 33246 9391 33302
rect 9447 33246 9533 33302
rect 9589 33246 9675 33302
rect 9731 33246 9817 33302
rect 9873 33246 9959 33302
rect 10015 33246 10101 33302
rect 10157 33246 10243 33302
rect 10299 33246 10385 33302
rect 10441 33246 10527 33302
rect 10583 33246 10669 33302
rect 10725 33246 10811 33302
rect 10867 33246 10953 33302
rect 11009 33246 11095 33302
rect 11151 33246 11237 33302
rect 11293 33246 11379 33302
rect 11435 33246 11521 33302
rect 11577 33246 11663 33302
rect 11719 33246 11805 33302
rect 11861 33246 11947 33302
rect 12003 33246 12089 33302
rect 12145 33246 12231 33302
rect 12287 33246 12373 33302
rect 12429 33246 12515 33302
rect 12571 33246 12657 33302
rect 12713 33246 12799 33302
rect 12855 33246 12941 33302
rect 12997 33246 13083 33302
rect 13139 33246 13225 33302
rect 13281 33246 13367 33302
rect 13423 33246 13509 33302
rect 13565 33246 13651 33302
rect 13707 33246 13793 33302
rect 13849 33246 13935 33302
rect 13991 33246 14077 33302
rect 14133 33246 14219 33302
rect 14275 33246 14361 33302
rect 14417 33246 14503 33302
rect 14559 33246 14645 33302
rect 14701 33246 14787 33302
rect 14843 33246 14853 33302
rect 151 33236 14853 33246
rect 151 32941 14853 32951
rect 151 32885 161 32941
rect 217 32885 303 32941
rect 359 32885 445 32941
rect 501 32885 587 32941
rect 643 32885 729 32941
rect 785 32885 871 32941
rect 927 32885 1013 32941
rect 1069 32885 1155 32941
rect 1211 32885 1297 32941
rect 1353 32885 1439 32941
rect 1495 32885 1581 32941
rect 1637 32885 1723 32941
rect 1779 32885 1865 32941
rect 1921 32885 2007 32941
rect 2063 32885 2149 32941
rect 2205 32885 2291 32941
rect 2347 32885 2433 32941
rect 2489 32885 2575 32941
rect 2631 32885 2717 32941
rect 2773 32885 2859 32941
rect 2915 32885 3001 32941
rect 3057 32885 3143 32941
rect 3199 32885 3285 32941
rect 3341 32885 3427 32941
rect 3483 32885 3569 32941
rect 3625 32885 3711 32941
rect 3767 32885 3853 32941
rect 3909 32885 3995 32941
rect 4051 32885 4137 32941
rect 4193 32885 4279 32941
rect 4335 32885 4421 32941
rect 4477 32885 4563 32941
rect 4619 32885 4705 32941
rect 4761 32885 4847 32941
rect 4903 32885 4989 32941
rect 5045 32885 5131 32941
rect 5187 32885 5273 32941
rect 5329 32885 5415 32941
rect 5471 32885 5557 32941
rect 5613 32885 5699 32941
rect 5755 32885 5841 32941
rect 5897 32885 5983 32941
rect 6039 32885 6125 32941
rect 6181 32885 6267 32941
rect 6323 32885 6409 32941
rect 6465 32885 6551 32941
rect 6607 32885 6693 32941
rect 6749 32885 6835 32941
rect 6891 32885 6977 32941
rect 7033 32885 7119 32941
rect 7175 32885 7261 32941
rect 7317 32885 7403 32941
rect 7459 32885 7545 32941
rect 7601 32885 7687 32941
rect 7743 32885 7829 32941
rect 7885 32885 7971 32941
rect 8027 32885 8113 32941
rect 8169 32885 8255 32941
rect 8311 32885 8397 32941
rect 8453 32885 8539 32941
rect 8595 32885 8681 32941
rect 8737 32885 8823 32941
rect 8879 32885 8965 32941
rect 9021 32885 9107 32941
rect 9163 32885 9249 32941
rect 9305 32885 9391 32941
rect 9447 32885 9533 32941
rect 9589 32885 9675 32941
rect 9731 32885 9817 32941
rect 9873 32885 9959 32941
rect 10015 32885 10101 32941
rect 10157 32885 10243 32941
rect 10299 32885 10385 32941
rect 10441 32885 10527 32941
rect 10583 32885 10669 32941
rect 10725 32885 10811 32941
rect 10867 32885 10953 32941
rect 11009 32885 11095 32941
rect 11151 32885 11237 32941
rect 11293 32885 11379 32941
rect 11435 32885 11521 32941
rect 11577 32885 11663 32941
rect 11719 32885 11805 32941
rect 11861 32885 11947 32941
rect 12003 32885 12089 32941
rect 12145 32885 12231 32941
rect 12287 32885 12373 32941
rect 12429 32885 12515 32941
rect 12571 32885 12657 32941
rect 12713 32885 12799 32941
rect 12855 32885 12941 32941
rect 12997 32885 13083 32941
rect 13139 32885 13225 32941
rect 13281 32885 13367 32941
rect 13423 32885 13509 32941
rect 13565 32885 13651 32941
rect 13707 32885 13793 32941
rect 13849 32885 13935 32941
rect 13991 32885 14077 32941
rect 14133 32885 14219 32941
rect 14275 32885 14361 32941
rect 14417 32885 14503 32941
rect 14559 32885 14645 32941
rect 14701 32885 14787 32941
rect 14843 32885 14853 32941
rect 151 32799 14853 32885
rect 151 32743 161 32799
rect 217 32743 303 32799
rect 359 32743 445 32799
rect 501 32743 587 32799
rect 643 32743 729 32799
rect 785 32743 871 32799
rect 927 32743 1013 32799
rect 1069 32743 1155 32799
rect 1211 32743 1297 32799
rect 1353 32743 1439 32799
rect 1495 32743 1581 32799
rect 1637 32743 1723 32799
rect 1779 32743 1865 32799
rect 1921 32743 2007 32799
rect 2063 32743 2149 32799
rect 2205 32743 2291 32799
rect 2347 32743 2433 32799
rect 2489 32743 2575 32799
rect 2631 32743 2717 32799
rect 2773 32743 2859 32799
rect 2915 32743 3001 32799
rect 3057 32743 3143 32799
rect 3199 32743 3285 32799
rect 3341 32743 3427 32799
rect 3483 32743 3569 32799
rect 3625 32743 3711 32799
rect 3767 32743 3853 32799
rect 3909 32743 3995 32799
rect 4051 32743 4137 32799
rect 4193 32743 4279 32799
rect 4335 32743 4421 32799
rect 4477 32743 4563 32799
rect 4619 32743 4705 32799
rect 4761 32743 4847 32799
rect 4903 32743 4989 32799
rect 5045 32743 5131 32799
rect 5187 32743 5273 32799
rect 5329 32743 5415 32799
rect 5471 32743 5557 32799
rect 5613 32743 5699 32799
rect 5755 32743 5841 32799
rect 5897 32743 5983 32799
rect 6039 32743 6125 32799
rect 6181 32743 6267 32799
rect 6323 32743 6409 32799
rect 6465 32743 6551 32799
rect 6607 32743 6693 32799
rect 6749 32743 6835 32799
rect 6891 32743 6977 32799
rect 7033 32743 7119 32799
rect 7175 32743 7261 32799
rect 7317 32743 7403 32799
rect 7459 32743 7545 32799
rect 7601 32743 7687 32799
rect 7743 32743 7829 32799
rect 7885 32743 7971 32799
rect 8027 32743 8113 32799
rect 8169 32743 8255 32799
rect 8311 32743 8397 32799
rect 8453 32743 8539 32799
rect 8595 32743 8681 32799
rect 8737 32743 8823 32799
rect 8879 32743 8965 32799
rect 9021 32743 9107 32799
rect 9163 32743 9249 32799
rect 9305 32743 9391 32799
rect 9447 32743 9533 32799
rect 9589 32743 9675 32799
rect 9731 32743 9817 32799
rect 9873 32743 9959 32799
rect 10015 32743 10101 32799
rect 10157 32743 10243 32799
rect 10299 32743 10385 32799
rect 10441 32743 10527 32799
rect 10583 32743 10669 32799
rect 10725 32743 10811 32799
rect 10867 32743 10953 32799
rect 11009 32743 11095 32799
rect 11151 32743 11237 32799
rect 11293 32743 11379 32799
rect 11435 32743 11521 32799
rect 11577 32743 11663 32799
rect 11719 32743 11805 32799
rect 11861 32743 11947 32799
rect 12003 32743 12089 32799
rect 12145 32743 12231 32799
rect 12287 32743 12373 32799
rect 12429 32743 12515 32799
rect 12571 32743 12657 32799
rect 12713 32743 12799 32799
rect 12855 32743 12941 32799
rect 12997 32743 13083 32799
rect 13139 32743 13225 32799
rect 13281 32743 13367 32799
rect 13423 32743 13509 32799
rect 13565 32743 13651 32799
rect 13707 32743 13793 32799
rect 13849 32743 13935 32799
rect 13991 32743 14077 32799
rect 14133 32743 14219 32799
rect 14275 32743 14361 32799
rect 14417 32743 14503 32799
rect 14559 32743 14645 32799
rect 14701 32743 14787 32799
rect 14843 32743 14853 32799
rect 151 32657 14853 32743
rect 151 32601 161 32657
rect 217 32601 303 32657
rect 359 32601 445 32657
rect 501 32601 587 32657
rect 643 32601 729 32657
rect 785 32601 871 32657
rect 927 32601 1013 32657
rect 1069 32601 1155 32657
rect 1211 32601 1297 32657
rect 1353 32601 1439 32657
rect 1495 32601 1581 32657
rect 1637 32601 1723 32657
rect 1779 32601 1865 32657
rect 1921 32601 2007 32657
rect 2063 32601 2149 32657
rect 2205 32601 2291 32657
rect 2347 32601 2433 32657
rect 2489 32601 2575 32657
rect 2631 32601 2717 32657
rect 2773 32601 2859 32657
rect 2915 32601 3001 32657
rect 3057 32601 3143 32657
rect 3199 32601 3285 32657
rect 3341 32601 3427 32657
rect 3483 32601 3569 32657
rect 3625 32601 3711 32657
rect 3767 32601 3853 32657
rect 3909 32601 3995 32657
rect 4051 32601 4137 32657
rect 4193 32601 4279 32657
rect 4335 32601 4421 32657
rect 4477 32601 4563 32657
rect 4619 32601 4705 32657
rect 4761 32601 4847 32657
rect 4903 32601 4989 32657
rect 5045 32601 5131 32657
rect 5187 32601 5273 32657
rect 5329 32601 5415 32657
rect 5471 32601 5557 32657
rect 5613 32601 5699 32657
rect 5755 32601 5841 32657
rect 5897 32601 5983 32657
rect 6039 32601 6125 32657
rect 6181 32601 6267 32657
rect 6323 32601 6409 32657
rect 6465 32601 6551 32657
rect 6607 32601 6693 32657
rect 6749 32601 6835 32657
rect 6891 32601 6977 32657
rect 7033 32601 7119 32657
rect 7175 32601 7261 32657
rect 7317 32601 7403 32657
rect 7459 32601 7545 32657
rect 7601 32601 7687 32657
rect 7743 32601 7829 32657
rect 7885 32601 7971 32657
rect 8027 32601 8113 32657
rect 8169 32601 8255 32657
rect 8311 32601 8397 32657
rect 8453 32601 8539 32657
rect 8595 32601 8681 32657
rect 8737 32601 8823 32657
rect 8879 32601 8965 32657
rect 9021 32601 9107 32657
rect 9163 32601 9249 32657
rect 9305 32601 9391 32657
rect 9447 32601 9533 32657
rect 9589 32601 9675 32657
rect 9731 32601 9817 32657
rect 9873 32601 9959 32657
rect 10015 32601 10101 32657
rect 10157 32601 10243 32657
rect 10299 32601 10385 32657
rect 10441 32601 10527 32657
rect 10583 32601 10669 32657
rect 10725 32601 10811 32657
rect 10867 32601 10953 32657
rect 11009 32601 11095 32657
rect 11151 32601 11237 32657
rect 11293 32601 11379 32657
rect 11435 32601 11521 32657
rect 11577 32601 11663 32657
rect 11719 32601 11805 32657
rect 11861 32601 11947 32657
rect 12003 32601 12089 32657
rect 12145 32601 12231 32657
rect 12287 32601 12373 32657
rect 12429 32601 12515 32657
rect 12571 32601 12657 32657
rect 12713 32601 12799 32657
rect 12855 32601 12941 32657
rect 12997 32601 13083 32657
rect 13139 32601 13225 32657
rect 13281 32601 13367 32657
rect 13423 32601 13509 32657
rect 13565 32601 13651 32657
rect 13707 32601 13793 32657
rect 13849 32601 13935 32657
rect 13991 32601 14077 32657
rect 14133 32601 14219 32657
rect 14275 32601 14361 32657
rect 14417 32601 14503 32657
rect 14559 32601 14645 32657
rect 14701 32601 14787 32657
rect 14843 32601 14853 32657
rect 151 32515 14853 32601
rect 151 32459 161 32515
rect 217 32459 303 32515
rect 359 32459 445 32515
rect 501 32459 587 32515
rect 643 32459 729 32515
rect 785 32459 871 32515
rect 927 32459 1013 32515
rect 1069 32459 1155 32515
rect 1211 32459 1297 32515
rect 1353 32459 1439 32515
rect 1495 32459 1581 32515
rect 1637 32459 1723 32515
rect 1779 32459 1865 32515
rect 1921 32459 2007 32515
rect 2063 32459 2149 32515
rect 2205 32459 2291 32515
rect 2347 32459 2433 32515
rect 2489 32459 2575 32515
rect 2631 32459 2717 32515
rect 2773 32459 2859 32515
rect 2915 32459 3001 32515
rect 3057 32459 3143 32515
rect 3199 32459 3285 32515
rect 3341 32459 3427 32515
rect 3483 32459 3569 32515
rect 3625 32459 3711 32515
rect 3767 32459 3853 32515
rect 3909 32459 3995 32515
rect 4051 32459 4137 32515
rect 4193 32459 4279 32515
rect 4335 32459 4421 32515
rect 4477 32459 4563 32515
rect 4619 32459 4705 32515
rect 4761 32459 4847 32515
rect 4903 32459 4989 32515
rect 5045 32459 5131 32515
rect 5187 32459 5273 32515
rect 5329 32459 5415 32515
rect 5471 32459 5557 32515
rect 5613 32459 5699 32515
rect 5755 32459 5841 32515
rect 5897 32459 5983 32515
rect 6039 32459 6125 32515
rect 6181 32459 6267 32515
rect 6323 32459 6409 32515
rect 6465 32459 6551 32515
rect 6607 32459 6693 32515
rect 6749 32459 6835 32515
rect 6891 32459 6977 32515
rect 7033 32459 7119 32515
rect 7175 32459 7261 32515
rect 7317 32459 7403 32515
rect 7459 32459 7545 32515
rect 7601 32459 7687 32515
rect 7743 32459 7829 32515
rect 7885 32459 7971 32515
rect 8027 32459 8113 32515
rect 8169 32459 8255 32515
rect 8311 32459 8397 32515
rect 8453 32459 8539 32515
rect 8595 32459 8681 32515
rect 8737 32459 8823 32515
rect 8879 32459 8965 32515
rect 9021 32459 9107 32515
rect 9163 32459 9249 32515
rect 9305 32459 9391 32515
rect 9447 32459 9533 32515
rect 9589 32459 9675 32515
rect 9731 32459 9817 32515
rect 9873 32459 9959 32515
rect 10015 32459 10101 32515
rect 10157 32459 10243 32515
rect 10299 32459 10385 32515
rect 10441 32459 10527 32515
rect 10583 32459 10669 32515
rect 10725 32459 10811 32515
rect 10867 32459 10953 32515
rect 11009 32459 11095 32515
rect 11151 32459 11237 32515
rect 11293 32459 11379 32515
rect 11435 32459 11521 32515
rect 11577 32459 11663 32515
rect 11719 32459 11805 32515
rect 11861 32459 11947 32515
rect 12003 32459 12089 32515
rect 12145 32459 12231 32515
rect 12287 32459 12373 32515
rect 12429 32459 12515 32515
rect 12571 32459 12657 32515
rect 12713 32459 12799 32515
rect 12855 32459 12941 32515
rect 12997 32459 13083 32515
rect 13139 32459 13225 32515
rect 13281 32459 13367 32515
rect 13423 32459 13509 32515
rect 13565 32459 13651 32515
rect 13707 32459 13793 32515
rect 13849 32459 13935 32515
rect 13991 32459 14077 32515
rect 14133 32459 14219 32515
rect 14275 32459 14361 32515
rect 14417 32459 14503 32515
rect 14559 32459 14645 32515
rect 14701 32459 14787 32515
rect 14843 32459 14853 32515
rect 151 32373 14853 32459
rect 151 32317 161 32373
rect 217 32317 303 32373
rect 359 32317 445 32373
rect 501 32317 587 32373
rect 643 32317 729 32373
rect 785 32317 871 32373
rect 927 32317 1013 32373
rect 1069 32317 1155 32373
rect 1211 32317 1297 32373
rect 1353 32317 1439 32373
rect 1495 32317 1581 32373
rect 1637 32317 1723 32373
rect 1779 32317 1865 32373
rect 1921 32317 2007 32373
rect 2063 32317 2149 32373
rect 2205 32317 2291 32373
rect 2347 32317 2433 32373
rect 2489 32317 2575 32373
rect 2631 32317 2717 32373
rect 2773 32317 2859 32373
rect 2915 32317 3001 32373
rect 3057 32317 3143 32373
rect 3199 32317 3285 32373
rect 3341 32317 3427 32373
rect 3483 32317 3569 32373
rect 3625 32317 3711 32373
rect 3767 32317 3853 32373
rect 3909 32317 3995 32373
rect 4051 32317 4137 32373
rect 4193 32317 4279 32373
rect 4335 32317 4421 32373
rect 4477 32317 4563 32373
rect 4619 32317 4705 32373
rect 4761 32317 4847 32373
rect 4903 32317 4989 32373
rect 5045 32317 5131 32373
rect 5187 32317 5273 32373
rect 5329 32317 5415 32373
rect 5471 32317 5557 32373
rect 5613 32317 5699 32373
rect 5755 32317 5841 32373
rect 5897 32317 5983 32373
rect 6039 32317 6125 32373
rect 6181 32317 6267 32373
rect 6323 32317 6409 32373
rect 6465 32317 6551 32373
rect 6607 32317 6693 32373
rect 6749 32317 6835 32373
rect 6891 32317 6977 32373
rect 7033 32317 7119 32373
rect 7175 32317 7261 32373
rect 7317 32317 7403 32373
rect 7459 32317 7545 32373
rect 7601 32317 7687 32373
rect 7743 32317 7829 32373
rect 7885 32317 7971 32373
rect 8027 32317 8113 32373
rect 8169 32317 8255 32373
rect 8311 32317 8397 32373
rect 8453 32317 8539 32373
rect 8595 32317 8681 32373
rect 8737 32317 8823 32373
rect 8879 32317 8965 32373
rect 9021 32317 9107 32373
rect 9163 32317 9249 32373
rect 9305 32317 9391 32373
rect 9447 32317 9533 32373
rect 9589 32317 9675 32373
rect 9731 32317 9817 32373
rect 9873 32317 9959 32373
rect 10015 32317 10101 32373
rect 10157 32317 10243 32373
rect 10299 32317 10385 32373
rect 10441 32317 10527 32373
rect 10583 32317 10669 32373
rect 10725 32317 10811 32373
rect 10867 32317 10953 32373
rect 11009 32317 11095 32373
rect 11151 32317 11237 32373
rect 11293 32317 11379 32373
rect 11435 32317 11521 32373
rect 11577 32317 11663 32373
rect 11719 32317 11805 32373
rect 11861 32317 11947 32373
rect 12003 32317 12089 32373
rect 12145 32317 12231 32373
rect 12287 32317 12373 32373
rect 12429 32317 12515 32373
rect 12571 32317 12657 32373
rect 12713 32317 12799 32373
rect 12855 32317 12941 32373
rect 12997 32317 13083 32373
rect 13139 32317 13225 32373
rect 13281 32317 13367 32373
rect 13423 32317 13509 32373
rect 13565 32317 13651 32373
rect 13707 32317 13793 32373
rect 13849 32317 13935 32373
rect 13991 32317 14077 32373
rect 14133 32317 14219 32373
rect 14275 32317 14361 32373
rect 14417 32317 14503 32373
rect 14559 32317 14645 32373
rect 14701 32317 14787 32373
rect 14843 32317 14853 32373
rect 151 32231 14853 32317
rect 151 32175 161 32231
rect 217 32175 303 32231
rect 359 32175 445 32231
rect 501 32175 587 32231
rect 643 32175 729 32231
rect 785 32175 871 32231
rect 927 32175 1013 32231
rect 1069 32175 1155 32231
rect 1211 32175 1297 32231
rect 1353 32175 1439 32231
rect 1495 32175 1581 32231
rect 1637 32175 1723 32231
rect 1779 32175 1865 32231
rect 1921 32175 2007 32231
rect 2063 32175 2149 32231
rect 2205 32175 2291 32231
rect 2347 32175 2433 32231
rect 2489 32175 2575 32231
rect 2631 32175 2717 32231
rect 2773 32175 2859 32231
rect 2915 32175 3001 32231
rect 3057 32175 3143 32231
rect 3199 32175 3285 32231
rect 3341 32175 3427 32231
rect 3483 32175 3569 32231
rect 3625 32175 3711 32231
rect 3767 32175 3853 32231
rect 3909 32175 3995 32231
rect 4051 32175 4137 32231
rect 4193 32175 4279 32231
rect 4335 32175 4421 32231
rect 4477 32175 4563 32231
rect 4619 32175 4705 32231
rect 4761 32175 4847 32231
rect 4903 32175 4989 32231
rect 5045 32175 5131 32231
rect 5187 32175 5273 32231
rect 5329 32175 5415 32231
rect 5471 32175 5557 32231
rect 5613 32175 5699 32231
rect 5755 32175 5841 32231
rect 5897 32175 5983 32231
rect 6039 32175 6125 32231
rect 6181 32175 6267 32231
rect 6323 32175 6409 32231
rect 6465 32175 6551 32231
rect 6607 32175 6693 32231
rect 6749 32175 6835 32231
rect 6891 32175 6977 32231
rect 7033 32175 7119 32231
rect 7175 32175 7261 32231
rect 7317 32175 7403 32231
rect 7459 32175 7545 32231
rect 7601 32175 7687 32231
rect 7743 32175 7829 32231
rect 7885 32175 7971 32231
rect 8027 32175 8113 32231
rect 8169 32175 8255 32231
rect 8311 32175 8397 32231
rect 8453 32175 8539 32231
rect 8595 32175 8681 32231
rect 8737 32175 8823 32231
rect 8879 32175 8965 32231
rect 9021 32175 9107 32231
rect 9163 32175 9249 32231
rect 9305 32175 9391 32231
rect 9447 32175 9533 32231
rect 9589 32175 9675 32231
rect 9731 32175 9817 32231
rect 9873 32175 9959 32231
rect 10015 32175 10101 32231
rect 10157 32175 10243 32231
rect 10299 32175 10385 32231
rect 10441 32175 10527 32231
rect 10583 32175 10669 32231
rect 10725 32175 10811 32231
rect 10867 32175 10953 32231
rect 11009 32175 11095 32231
rect 11151 32175 11237 32231
rect 11293 32175 11379 32231
rect 11435 32175 11521 32231
rect 11577 32175 11663 32231
rect 11719 32175 11805 32231
rect 11861 32175 11947 32231
rect 12003 32175 12089 32231
rect 12145 32175 12231 32231
rect 12287 32175 12373 32231
rect 12429 32175 12515 32231
rect 12571 32175 12657 32231
rect 12713 32175 12799 32231
rect 12855 32175 12941 32231
rect 12997 32175 13083 32231
rect 13139 32175 13225 32231
rect 13281 32175 13367 32231
rect 13423 32175 13509 32231
rect 13565 32175 13651 32231
rect 13707 32175 13793 32231
rect 13849 32175 13935 32231
rect 13991 32175 14077 32231
rect 14133 32175 14219 32231
rect 14275 32175 14361 32231
rect 14417 32175 14503 32231
rect 14559 32175 14645 32231
rect 14701 32175 14787 32231
rect 14843 32175 14853 32231
rect 151 32089 14853 32175
rect 151 32033 161 32089
rect 217 32033 303 32089
rect 359 32033 445 32089
rect 501 32033 587 32089
rect 643 32033 729 32089
rect 785 32033 871 32089
rect 927 32033 1013 32089
rect 1069 32033 1155 32089
rect 1211 32033 1297 32089
rect 1353 32033 1439 32089
rect 1495 32033 1581 32089
rect 1637 32033 1723 32089
rect 1779 32033 1865 32089
rect 1921 32033 2007 32089
rect 2063 32033 2149 32089
rect 2205 32033 2291 32089
rect 2347 32033 2433 32089
rect 2489 32033 2575 32089
rect 2631 32033 2717 32089
rect 2773 32033 2859 32089
rect 2915 32033 3001 32089
rect 3057 32033 3143 32089
rect 3199 32033 3285 32089
rect 3341 32033 3427 32089
rect 3483 32033 3569 32089
rect 3625 32033 3711 32089
rect 3767 32033 3853 32089
rect 3909 32033 3995 32089
rect 4051 32033 4137 32089
rect 4193 32033 4279 32089
rect 4335 32033 4421 32089
rect 4477 32033 4563 32089
rect 4619 32033 4705 32089
rect 4761 32033 4847 32089
rect 4903 32033 4989 32089
rect 5045 32033 5131 32089
rect 5187 32033 5273 32089
rect 5329 32033 5415 32089
rect 5471 32033 5557 32089
rect 5613 32033 5699 32089
rect 5755 32033 5841 32089
rect 5897 32033 5983 32089
rect 6039 32033 6125 32089
rect 6181 32033 6267 32089
rect 6323 32033 6409 32089
rect 6465 32033 6551 32089
rect 6607 32033 6693 32089
rect 6749 32033 6835 32089
rect 6891 32033 6977 32089
rect 7033 32033 7119 32089
rect 7175 32033 7261 32089
rect 7317 32033 7403 32089
rect 7459 32033 7545 32089
rect 7601 32033 7687 32089
rect 7743 32033 7829 32089
rect 7885 32033 7971 32089
rect 8027 32033 8113 32089
rect 8169 32033 8255 32089
rect 8311 32033 8397 32089
rect 8453 32033 8539 32089
rect 8595 32033 8681 32089
rect 8737 32033 8823 32089
rect 8879 32033 8965 32089
rect 9021 32033 9107 32089
rect 9163 32033 9249 32089
rect 9305 32033 9391 32089
rect 9447 32033 9533 32089
rect 9589 32033 9675 32089
rect 9731 32033 9817 32089
rect 9873 32033 9959 32089
rect 10015 32033 10101 32089
rect 10157 32033 10243 32089
rect 10299 32033 10385 32089
rect 10441 32033 10527 32089
rect 10583 32033 10669 32089
rect 10725 32033 10811 32089
rect 10867 32033 10953 32089
rect 11009 32033 11095 32089
rect 11151 32033 11237 32089
rect 11293 32033 11379 32089
rect 11435 32033 11521 32089
rect 11577 32033 11663 32089
rect 11719 32033 11805 32089
rect 11861 32033 11947 32089
rect 12003 32033 12089 32089
rect 12145 32033 12231 32089
rect 12287 32033 12373 32089
rect 12429 32033 12515 32089
rect 12571 32033 12657 32089
rect 12713 32033 12799 32089
rect 12855 32033 12941 32089
rect 12997 32033 13083 32089
rect 13139 32033 13225 32089
rect 13281 32033 13367 32089
rect 13423 32033 13509 32089
rect 13565 32033 13651 32089
rect 13707 32033 13793 32089
rect 13849 32033 13935 32089
rect 13991 32033 14077 32089
rect 14133 32033 14219 32089
rect 14275 32033 14361 32089
rect 14417 32033 14503 32089
rect 14559 32033 14645 32089
rect 14701 32033 14787 32089
rect 14843 32033 14853 32089
rect 151 31947 14853 32033
rect 151 31891 161 31947
rect 217 31891 303 31947
rect 359 31891 445 31947
rect 501 31891 587 31947
rect 643 31891 729 31947
rect 785 31891 871 31947
rect 927 31891 1013 31947
rect 1069 31891 1155 31947
rect 1211 31891 1297 31947
rect 1353 31891 1439 31947
rect 1495 31891 1581 31947
rect 1637 31891 1723 31947
rect 1779 31891 1865 31947
rect 1921 31891 2007 31947
rect 2063 31891 2149 31947
rect 2205 31891 2291 31947
rect 2347 31891 2433 31947
rect 2489 31891 2575 31947
rect 2631 31891 2717 31947
rect 2773 31891 2859 31947
rect 2915 31891 3001 31947
rect 3057 31891 3143 31947
rect 3199 31891 3285 31947
rect 3341 31891 3427 31947
rect 3483 31891 3569 31947
rect 3625 31891 3711 31947
rect 3767 31891 3853 31947
rect 3909 31891 3995 31947
rect 4051 31891 4137 31947
rect 4193 31891 4279 31947
rect 4335 31891 4421 31947
rect 4477 31891 4563 31947
rect 4619 31891 4705 31947
rect 4761 31891 4847 31947
rect 4903 31891 4989 31947
rect 5045 31891 5131 31947
rect 5187 31891 5273 31947
rect 5329 31891 5415 31947
rect 5471 31891 5557 31947
rect 5613 31891 5699 31947
rect 5755 31891 5841 31947
rect 5897 31891 5983 31947
rect 6039 31891 6125 31947
rect 6181 31891 6267 31947
rect 6323 31891 6409 31947
rect 6465 31891 6551 31947
rect 6607 31891 6693 31947
rect 6749 31891 6835 31947
rect 6891 31891 6977 31947
rect 7033 31891 7119 31947
rect 7175 31891 7261 31947
rect 7317 31891 7403 31947
rect 7459 31891 7545 31947
rect 7601 31891 7687 31947
rect 7743 31891 7829 31947
rect 7885 31891 7971 31947
rect 8027 31891 8113 31947
rect 8169 31891 8255 31947
rect 8311 31891 8397 31947
rect 8453 31891 8539 31947
rect 8595 31891 8681 31947
rect 8737 31891 8823 31947
rect 8879 31891 8965 31947
rect 9021 31891 9107 31947
rect 9163 31891 9249 31947
rect 9305 31891 9391 31947
rect 9447 31891 9533 31947
rect 9589 31891 9675 31947
rect 9731 31891 9817 31947
rect 9873 31891 9959 31947
rect 10015 31891 10101 31947
rect 10157 31891 10243 31947
rect 10299 31891 10385 31947
rect 10441 31891 10527 31947
rect 10583 31891 10669 31947
rect 10725 31891 10811 31947
rect 10867 31891 10953 31947
rect 11009 31891 11095 31947
rect 11151 31891 11237 31947
rect 11293 31891 11379 31947
rect 11435 31891 11521 31947
rect 11577 31891 11663 31947
rect 11719 31891 11805 31947
rect 11861 31891 11947 31947
rect 12003 31891 12089 31947
rect 12145 31891 12231 31947
rect 12287 31891 12373 31947
rect 12429 31891 12515 31947
rect 12571 31891 12657 31947
rect 12713 31891 12799 31947
rect 12855 31891 12941 31947
rect 12997 31891 13083 31947
rect 13139 31891 13225 31947
rect 13281 31891 13367 31947
rect 13423 31891 13509 31947
rect 13565 31891 13651 31947
rect 13707 31891 13793 31947
rect 13849 31891 13935 31947
rect 13991 31891 14077 31947
rect 14133 31891 14219 31947
rect 14275 31891 14361 31947
rect 14417 31891 14503 31947
rect 14559 31891 14645 31947
rect 14701 31891 14787 31947
rect 14843 31891 14853 31947
rect 151 31805 14853 31891
rect 151 31749 161 31805
rect 217 31749 303 31805
rect 359 31749 445 31805
rect 501 31749 587 31805
rect 643 31749 729 31805
rect 785 31749 871 31805
rect 927 31749 1013 31805
rect 1069 31749 1155 31805
rect 1211 31749 1297 31805
rect 1353 31749 1439 31805
rect 1495 31749 1581 31805
rect 1637 31749 1723 31805
rect 1779 31749 1865 31805
rect 1921 31749 2007 31805
rect 2063 31749 2149 31805
rect 2205 31749 2291 31805
rect 2347 31749 2433 31805
rect 2489 31749 2575 31805
rect 2631 31749 2717 31805
rect 2773 31749 2859 31805
rect 2915 31749 3001 31805
rect 3057 31749 3143 31805
rect 3199 31749 3285 31805
rect 3341 31749 3427 31805
rect 3483 31749 3569 31805
rect 3625 31749 3711 31805
rect 3767 31749 3853 31805
rect 3909 31749 3995 31805
rect 4051 31749 4137 31805
rect 4193 31749 4279 31805
rect 4335 31749 4421 31805
rect 4477 31749 4563 31805
rect 4619 31749 4705 31805
rect 4761 31749 4847 31805
rect 4903 31749 4989 31805
rect 5045 31749 5131 31805
rect 5187 31749 5273 31805
rect 5329 31749 5415 31805
rect 5471 31749 5557 31805
rect 5613 31749 5699 31805
rect 5755 31749 5841 31805
rect 5897 31749 5983 31805
rect 6039 31749 6125 31805
rect 6181 31749 6267 31805
rect 6323 31749 6409 31805
rect 6465 31749 6551 31805
rect 6607 31749 6693 31805
rect 6749 31749 6835 31805
rect 6891 31749 6977 31805
rect 7033 31749 7119 31805
rect 7175 31749 7261 31805
rect 7317 31749 7403 31805
rect 7459 31749 7545 31805
rect 7601 31749 7687 31805
rect 7743 31749 7829 31805
rect 7885 31749 7971 31805
rect 8027 31749 8113 31805
rect 8169 31749 8255 31805
rect 8311 31749 8397 31805
rect 8453 31749 8539 31805
rect 8595 31749 8681 31805
rect 8737 31749 8823 31805
rect 8879 31749 8965 31805
rect 9021 31749 9107 31805
rect 9163 31749 9249 31805
rect 9305 31749 9391 31805
rect 9447 31749 9533 31805
rect 9589 31749 9675 31805
rect 9731 31749 9817 31805
rect 9873 31749 9959 31805
rect 10015 31749 10101 31805
rect 10157 31749 10243 31805
rect 10299 31749 10385 31805
rect 10441 31749 10527 31805
rect 10583 31749 10669 31805
rect 10725 31749 10811 31805
rect 10867 31749 10953 31805
rect 11009 31749 11095 31805
rect 11151 31749 11237 31805
rect 11293 31749 11379 31805
rect 11435 31749 11521 31805
rect 11577 31749 11663 31805
rect 11719 31749 11805 31805
rect 11861 31749 11947 31805
rect 12003 31749 12089 31805
rect 12145 31749 12231 31805
rect 12287 31749 12373 31805
rect 12429 31749 12515 31805
rect 12571 31749 12657 31805
rect 12713 31749 12799 31805
rect 12855 31749 12941 31805
rect 12997 31749 13083 31805
rect 13139 31749 13225 31805
rect 13281 31749 13367 31805
rect 13423 31749 13509 31805
rect 13565 31749 13651 31805
rect 13707 31749 13793 31805
rect 13849 31749 13935 31805
rect 13991 31749 14077 31805
rect 14133 31749 14219 31805
rect 14275 31749 14361 31805
rect 14417 31749 14503 31805
rect 14559 31749 14645 31805
rect 14701 31749 14787 31805
rect 14843 31749 14853 31805
rect 151 31663 14853 31749
rect 151 31607 161 31663
rect 217 31607 303 31663
rect 359 31607 445 31663
rect 501 31607 587 31663
rect 643 31607 729 31663
rect 785 31607 871 31663
rect 927 31607 1013 31663
rect 1069 31607 1155 31663
rect 1211 31607 1297 31663
rect 1353 31607 1439 31663
rect 1495 31607 1581 31663
rect 1637 31607 1723 31663
rect 1779 31607 1865 31663
rect 1921 31607 2007 31663
rect 2063 31607 2149 31663
rect 2205 31607 2291 31663
rect 2347 31607 2433 31663
rect 2489 31607 2575 31663
rect 2631 31607 2717 31663
rect 2773 31607 2859 31663
rect 2915 31607 3001 31663
rect 3057 31607 3143 31663
rect 3199 31607 3285 31663
rect 3341 31607 3427 31663
rect 3483 31607 3569 31663
rect 3625 31607 3711 31663
rect 3767 31607 3853 31663
rect 3909 31607 3995 31663
rect 4051 31607 4137 31663
rect 4193 31607 4279 31663
rect 4335 31607 4421 31663
rect 4477 31607 4563 31663
rect 4619 31607 4705 31663
rect 4761 31607 4847 31663
rect 4903 31607 4989 31663
rect 5045 31607 5131 31663
rect 5187 31607 5273 31663
rect 5329 31607 5415 31663
rect 5471 31607 5557 31663
rect 5613 31607 5699 31663
rect 5755 31607 5841 31663
rect 5897 31607 5983 31663
rect 6039 31607 6125 31663
rect 6181 31607 6267 31663
rect 6323 31607 6409 31663
rect 6465 31607 6551 31663
rect 6607 31607 6693 31663
rect 6749 31607 6835 31663
rect 6891 31607 6977 31663
rect 7033 31607 7119 31663
rect 7175 31607 7261 31663
rect 7317 31607 7403 31663
rect 7459 31607 7545 31663
rect 7601 31607 7687 31663
rect 7743 31607 7829 31663
rect 7885 31607 7971 31663
rect 8027 31607 8113 31663
rect 8169 31607 8255 31663
rect 8311 31607 8397 31663
rect 8453 31607 8539 31663
rect 8595 31607 8681 31663
rect 8737 31607 8823 31663
rect 8879 31607 8965 31663
rect 9021 31607 9107 31663
rect 9163 31607 9249 31663
rect 9305 31607 9391 31663
rect 9447 31607 9533 31663
rect 9589 31607 9675 31663
rect 9731 31607 9817 31663
rect 9873 31607 9959 31663
rect 10015 31607 10101 31663
rect 10157 31607 10243 31663
rect 10299 31607 10385 31663
rect 10441 31607 10527 31663
rect 10583 31607 10669 31663
rect 10725 31607 10811 31663
rect 10867 31607 10953 31663
rect 11009 31607 11095 31663
rect 11151 31607 11237 31663
rect 11293 31607 11379 31663
rect 11435 31607 11521 31663
rect 11577 31607 11663 31663
rect 11719 31607 11805 31663
rect 11861 31607 11947 31663
rect 12003 31607 12089 31663
rect 12145 31607 12231 31663
rect 12287 31607 12373 31663
rect 12429 31607 12515 31663
rect 12571 31607 12657 31663
rect 12713 31607 12799 31663
rect 12855 31607 12941 31663
rect 12997 31607 13083 31663
rect 13139 31607 13225 31663
rect 13281 31607 13367 31663
rect 13423 31607 13509 31663
rect 13565 31607 13651 31663
rect 13707 31607 13793 31663
rect 13849 31607 13935 31663
rect 13991 31607 14077 31663
rect 14133 31607 14219 31663
rect 14275 31607 14361 31663
rect 14417 31607 14503 31663
rect 14559 31607 14645 31663
rect 14701 31607 14787 31663
rect 14843 31607 14853 31663
rect 151 31521 14853 31607
rect 151 31465 161 31521
rect 217 31465 303 31521
rect 359 31465 445 31521
rect 501 31465 587 31521
rect 643 31465 729 31521
rect 785 31465 871 31521
rect 927 31465 1013 31521
rect 1069 31465 1155 31521
rect 1211 31465 1297 31521
rect 1353 31465 1439 31521
rect 1495 31465 1581 31521
rect 1637 31465 1723 31521
rect 1779 31465 1865 31521
rect 1921 31465 2007 31521
rect 2063 31465 2149 31521
rect 2205 31465 2291 31521
rect 2347 31465 2433 31521
rect 2489 31465 2575 31521
rect 2631 31465 2717 31521
rect 2773 31465 2859 31521
rect 2915 31465 3001 31521
rect 3057 31465 3143 31521
rect 3199 31465 3285 31521
rect 3341 31465 3427 31521
rect 3483 31465 3569 31521
rect 3625 31465 3711 31521
rect 3767 31465 3853 31521
rect 3909 31465 3995 31521
rect 4051 31465 4137 31521
rect 4193 31465 4279 31521
rect 4335 31465 4421 31521
rect 4477 31465 4563 31521
rect 4619 31465 4705 31521
rect 4761 31465 4847 31521
rect 4903 31465 4989 31521
rect 5045 31465 5131 31521
rect 5187 31465 5273 31521
rect 5329 31465 5415 31521
rect 5471 31465 5557 31521
rect 5613 31465 5699 31521
rect 5755 31465 5841 31521
rect 5897 31465 5983 31521
rect 6039 31465 6125 31521
rect 6181 31465 6267 31521
rect 6323 31465 6409 31521
rect 6465 31465 6551 31521
rect 6607 31465 6693 31521
rect 6749 31465 6835 31521
rect 6891 31465 6977 31521
rect 7033 31465 7119 31521
rect 7175 31465 7261 31521
rect 7317 31465 7403 31521
rect 7459 31465 7545 31521
rect 7601 31465 7687 31521
rect 7743 31465 7829 31521
rect 7885 31465 7971 31521
rect 8027 31465 8113 31521
rect 8169 31465 8255 31521
rect 8311 31465 8397 31521
rect 8453 31465 8539 31521
rect 8595 31465 8681 31521
rect 8737 31465 8823 31521
rect 8879 31465 8965 31521
rect 9021 31465 9107 31521
rect 9163 31465 9249 31521
rect 9305 31465 9391 31521
rect 9447 31465 9533 31521
rect 9589 31465 9675 31521
rect 9731 31465 9817 31521
rect 9873 31465 9959 31521
rect 10015 31465 10101 31521
rect 10157 31465 10243 31521
rect 10299 31465 10385 31521
rect 10441 31465 10527 31521
rect 10583 31465 10669 31521
rect 10725 31465 10811 31521
rect 10867 31465 10953 31521
rect 11009 31465 11095 31521
rect 11151 31465 11237 31521
rect 11293 31465 11379 31521
rect 11435 31465 11521 31521
rect 11577 31465 11663 31521
rect 11719 31465 11805 31521
rect 11861 31465 11947 31521
rect 12003 31465 12089 31521
rect 12145 31465 12231 31521
rect 12287 31465 12373 31521
rect 12429 31465 12515 31521
rect 12571 31465 12657 31521
rect 12713 31465 12799 31521
rect 12855 31465 12941 31521
rect 12997 31465 13083 31521
rect 13139 31465 13225 31521
rect 13281 31465 13367 31521
rect 13423 31465 13509 31521
rect 13565 31465 13651 31521
rect 13707 31465 13793 31521
rect 13849 31465 13935 31521
rect 13991 31465 14077 31521
rect 14133 31465 14219 31521
rect 14275 31465 14361 31521
rect 14417 31465 14503 31521
rect 14559 31465 14645 31521
rect 14701 31465 14787 31521
rect 14843 31465 14853 31521
rect 151 31379 14853 31465
rect 151 31323 161 31379
rect 217 31323 303 31379
rect 359 31323 445 31379
rect 501 31323 587 31379
rect 643 31323 729 31379
rect 785 31323 871 31379
rect 927 31323 1013 31379
rect 1069 31323 1155 31379
rect 1211 31323 1297 31379
rect 1353 31323 1439 31379
rect 1495 31323 1581 31379
rect 1637 31323 1723 31379
rect 1779 31323 1865 31379
rect 1921 31323 2007 31379
rect 2063 31323 2149 31379
rect 2205 31323 2291 31379
rect 2347 31323 2433 31379
rect 2489 31323 2575 31379
rect 2631 31323 2717 31379
rect 2773 31323 2859 31379
rect 2915 31323 3001 31379
rect 3057 31323 3143 31379
rect 3199 31323 3285 31379
rect 3341 31323 3427 31379
rect 3483 31323 3569 31379
rect 3625 31323 3711 31379
rect 3767 31323 3853 31379
rect 3909 31323 3995 31379
rect 4051 31323 4137 31379
rect 4193 31323 4279 31379
rect 4335 31323 4421 31379
rect 4477 31323 4563 31379
rect 4619 31323 4705 31379
rect 4761 31323 4847 31379
rect 4903 31323 4989 31379
rect 5045 31323 5131 31379
rect 5187 31323 5273 31379
rect 5329 31323 5415 31379
rect 5471 31323 5557 31379
rect 5613 31323 5699 31379
rect 5755 31323 5841 31379
rect 5897 31323 5983 31379
rect 6039 31323 6125 31379
rect 6181 31323 6267 31379
rect 6323 31323 6409 31379
rect 6465 31323 6551 31379
rect 6607 31323 6693 31379
rect 6749 31323 6835 31379
rect 6891 31323 6977 31379
rect 7033 31323 7119 31379
rect 7175 31323 7261 31379
rect 7317 31323 7403 31379
rect 7459 31323 7545 31379
rect 7601 31323 7687 31379
rect 7743 31323 7829 31379
rect 7885 31323 7971 31379
rect 8027 31323 8113 31379
rect 8169 31323 8255 31379
rect 8311 31323 8397 31379
rect 8453 31323 8539 31379
rect 8595 31323 8681 31379
rect 8737 31323 8823 31379
rect 8879 31323 8965 31379
rect 9021 31323 9107 31379
rect 9163 31323 9249 31379
rect 9305 31323 9391 31379
rect 9447 31323 9533 31379
rect 9589 31323 9675 31379
rect 9731 31323 9817 31379
rect 9873 31323 9959 31379
rect 10015 31323 10101 31379
rect 10157 31323 10243 31379
rect 10299 31323 10385 31379
rect 10441 31323 10527 31379
rect 10583 31323 10669 31379
rect 10725 31323 10811 31379
rect 10867 31323 10953 31379
rect 11009 31323 11095 31379
rect 11151 31323 11237 31379
rect 11293 31323 11379 31379
rect 11435 31323 11521 31379
rect 11577 31323 11663 31379
rect 11719 31323 11805 31379
rect 11861 31323 11947 31379
rect 12003 31323 12089 31379
rect 12145 31323 12231 31379
rect 12287 31323 12373 31379
rect 12429 31323 12515 31379
rect 12571 31323 12657 31379
rect 12713 31323 12799 31379
rect 12855 31323 12941 31379
rect 12997 31323 13083 31379
rect 13139 31323 13225 31379
rect 13281 31323 13367 31379
rect 13423 31323 13509 31379
rect 13565 31323 13651 31379
rect 13707 31323 13793 31379
rect 13849 31323 13935 31379
rect 13991 31323 14077 31379
rect 14133 31323 14219 31379
rect 14275 31323 14361 31379
rect 14417 31323 14503 31379
rect 14559 31323 14645 31379
rect 14701 31323 14787 31379
rect 14843 31323 14853 31379
rect 151 31237 14853 31323
rect 151 31181 161 31237
rect 217 31181 303 31237
rect 359 31181 445 31237
rect 501 31181 587 31237
rect 643 31181 729 31237
rect 785 31181 871 31237
rect 927 31181 1013 31237
rect 1069 31181 1155 31237
rect 1211 31181 1297 31237
rect 1353 31181 1439 31237
rect 1495 31181 1581 31237
rect 1637 31181 1723 31237
rect 1779 31181 1865 31237
rect 1921 31181 2007 31237
rect 2063 31181 2149 31237
rect 2205 31181 2291 31237
rect 2347 31181 2433 31237
rect 2489 31181 2575 31237
rect 2631 31181 2717 31237
rect 2773 31181 2859 31237
rect 2915 31181 3001 31237
rect 3057 31181 3143 31237
rect 3199 31181 3285 31237
rect 3341 31181 3427 31237
rect 3483 31181 3569 31237
rect 3625 31181 3711 31237
rect 3767 31181 3853 31237
rect 3909 31181 3995 31237
rect 4051 31181 4137 31237
rect 4193 31181 4279 31237
rect 4335 31181 4421 31237
rect 4477 31181 4563 31237
rect 4619 31181 4705 31237
rect 4761 31181 4847 31237
rect 4903 31181 4989 31237
rect 5045 31181 5131 31237
rect 5187 31181 5273 31237
rect 5329 31181 5415 31237
rect 5471 31181 5557 31237
rect 5613 31181 5699 31237
rect 5755 31181 5841 31237
rect 5897 31181 5983 31237
rect 6039 31181 6125 31237
rect 6181 31181 6267 31237
rect 6323 31181 6409 31237
rect 6465 31181 6551 31237
rect 6607 31181 6693 31237
rect 6749 31181 6835 31237
rect 6891 31181 6977 31237
rect 7033 31181 7119 31237
rect 7175 31181 7261 31237
rect 7317 31181 7403 31237
rect 7459 31181 7545 31237
rect 7601 31181 7687 31237
rect 7743 31181 7829 31237
rect 7885 31181 7971 31237
rect 8027 31181 8113 31237
rect 8169 31181 8255 31237
rect 8311 31181 8397 31237
rect 8453 31181 8539 31237
rect 8595 31181 8681 31237
rect 8737 31181 8823 31237
rect 8879 31181 8965 31237
rect 9021 31181 9107 31237
rect 9163 31181 9249 31237
rect 9305 31181 9391 31237
rect 9447 31181 9533 31237
rect 9589 31181 9675 31237
rect 9731 31181 9817 31237
rect 9873 31181 9959 31237
rect 10015 31181 10101 31237
rect 10157 31181 10243 31237
rect 10299 31181 10385 31237
rect 10441 31181 10527 31237
rect 10583 31181 10669 31237
rect 10725 31181 10811 31237
rect 10867 31181 10953 31237
rect 11009 31181 11095 31237
rect 11151 31181 11237 31237
rect 11293 31181 11379 31237
rect 11435 31181 11521 31237
rect 11577 31181 11663 31237
rect 11719 31181 11805 31237
rect 11861 31181 11947 31237
rect 12003 31181 12089 31237
rect 12145 31181 12231 31237
rect 12287 31181 12373 31237
rect 12429 31181 12515 31237
rect 12571 31181 12657 31237
rect 12713 31181 12799 31237
rect 12855 31181 12941 31237
rect 12997 31181 13083 31237
rect 13139 31181 13225 31237
rect 13281 31181 13367 31237
rect 13423 31181 13509 31237
rect 13565 31181 13651 31237
rect 13707 31181 13793 31237
rect 13849 31181 13935 31237
rect 13991 31181 14077 31237
rect 14133 31181 14219 31237
rect 14275 31181 14361 31237
rect 14417 31181 14503 31237
rect 14559 31181 14645 31237
rect 14701 31181 14787 31237
rect 14843 31181 14853 31237
rect 151 31095 14853 31181
rect 151 31039 161 31095
rect 217 31039 303 31095
rect 359 31039 445 31095
rect 501 31039 587 31095
rect 643 31039 729 31095
rect 785 31039 871 31095
rect 927 31039 1013 31095
rect 1069 31039 1155 31095
rect 1211 31039 1297 31095
rect 1353 31039 1439 31095
rect 1495 31039 1581 31095
rect 1637 31039 1723 31095
rect 1779 31039 1865 31095
rect 1921 31039 2007 31095
rect 2063 31039 2149 31095
rect 2205 31039 2291 31095
rect 2347 31039 2433 31095
rect 2489 31039 2575 31095
rect 2631 31039 2717 31095
rect 2773 31039 2859 31095
rect 2915 31039 3001 31095
rect 3057 31039 3143 31095
rect 3199 31039 3285 31095
rect 3341 31039 3427 31095
rect 3483 31039 3569 31095
rect 3625 31039 3711 31095
rect 3767 31039 3853 31095
rect 3909 31039 3995 31095
rect 4051 31039 4137 31095
rect 4193 31039 4279 31095
rect 4335 31039 4421 31095
rect 4477 31039 4563 31095
rect 4619 31039 4705 31095
rect 4761 31039 4847 31095
rect 4903 31039 4989 31095
rect 5045 31039 5131 31095
rect 5187 31039 5273 31095
rect 5329 31039 5415 31095
rect 5471 31039 5557 31095
rect 5613 31039 5699 31095
rect 5755 31039 5841 31095
rect 5897 31039 5983 31095
rect 6039 31039 6125 31095
rect 6181 31039 6267 31095
rect 6323 31039 6409 31095
rect 6465 31039 6551 31095
rect 6607 31039 6693 31095
rect 6749 31039 6835 31095
rect 6891 31039 6977 31095
rect 7033 31039 7119 31095
rect 7175 31039 7261 31095
rect 7317 31039 7403 31095
rect 7459 31039 7545 31095
rect 7601 31039 7687 31095
rect 7743 31039 7829 31095
rect 7885 31039 7971 31095
rect 8027 31039 8113 31095
rect 8169 31039 8255 31095
rect 8311 31039 8397 31095
rect 8453 31039 8539 31095
rect 8595 31039 8681 31095
rect 8737 31039 8823 31095
rect 8879 31039 8965 31095
rect 9021 31039 9107 31095
rect 9163 31039 9249 31095
rect 9305 31039 9391 31095
rect 9447 31039 9533 31095
rect 9589 31039 9675 31095
rect 9731 31039 9817 31095
rect 9873 31039 9959 31095
rect 10015 31039 10101 31095
rect 10157 31039 10243 31095
rect 10299 31039 10385 31095
rect 10441 31039 10527 31095
rect 10583 31039 10669 31095
rect 10725 31039 10811 31095
rect 10867 31039 10953 31095
rect 11009 31039 11095 31095
rect 11151 31039 11237 31095
rect 11293 31039 11379 31095
rect 11435 31039 11521 31095
rect 11577 31039 11663 31095
rect 11719 31039 11805 31095
rect 11861 31039 11947 31095
rect 12003 31039 12089 31095
rect 12145 31039 12231 31095
rect 12287 31039 12373 31095
rect 12429 31039 12515 31095
rect 12571 31039 12657 31095
rect 12713 31039 12799 31095
rect 12855 31039 12941 31095
rect 12997 31039 13083 31095
rect 13139 31039 13225 31095
rect 13281 31039 13367 31095
rect 13423 31039 13509 31095
rect 13565 31039 13651 31095
rect 13707 31039 13793 31095
rect 13849 31039 13935 31095
rect 13991 31039 14077 31095
rect 14133 31039 14219 31095
rect 14275 31039 14361 31095
rect 14417 31039 14503 31095
rect 14559 31039 14645 31095
rect 14701 31039 14787 31095
rect 14843 31039 14853 31095
rect 151 30953 14853 31039
rect 151 30897 161 30953
rect 217 30897 303 30953
rect 359 30897 445 30953
rect 501 30897 587 30953
rect 643 30897 729 30953
rect 785 30897 871 30953
rect 927 30897 1013 30953
rect 1069 30897 1155 30953
rect 1211 30897 1297 30953
rect 1353 30897 1439 30953
rect 1495 30897 1581 30953
rect 1637 30897 1723 30953
rect 1779 30897 1865 30953
rect 1921 30897 2007 30953
rect 2063 30897 2149 30953
rect 2205 30897 2291 30953
rect 2347 30897 2433 30953
rect 2489 30897 2575 30953
rect 2631 30897 2717 30953
rect 2773 30897 2859 30953
rect 2915 30897 3001 30953
rect 3057 30897 3143 30953
rect 3199 30897 3285 30953
rect 3341 30897 3427 30953
rect 3483 30897 3569 30953
rect 3625 30897 3711 30953
rect 3767 30897 3853 30953
rect 3909 30897 3995 30953
rect 4051 30897 4137 30953
rect 4193 30897 4279 30953
rect 4335 30897 4421 30953
rect 4477 30897 4563 30953
rect 4619 30897 4705 30953
rect 4761 30897 4847 30953
rect 4903 30897 4989 30953
rect 5045 30897 5131 30953
rect 5187 30897 5273 30953
rect 5329 30897 5415 30953
rect 5471 30897 5557 30953
rect 5613 30897 5699 30953
rect 5755 30897 5841 30953
rect 5897 30897 5983 30953
rect 6039 30897 6125 30953
rect 6181 30897 6267 30953
rect 6323 30897 6409 30953
rect 6465 30897 6551 30953
rect 6607 30897 6693 30953
rect 6749 30897 6835 30953
rect 6891 30897 6977 30953
rect 7033 30897 7119 30953
rect 7175 30897 7261 30953
rect 7317 30897 7403 30953
rect 7459 30897 7545 30953
rect 7601 30897 7687 30953
rect 7743 30897 7829 30953
rect 7885 30897 7971 30953
rect 8027 30897 8113 30953
rect 8169 30897 8255 30953
rect 8311 30897 8397 30953
rect 8453 30897 8539 30953
rect 8595 30897 8681 30953
rect 8737 30897 8823 30953
rect 8879 30897 8965 30953
rect 9021 30897 9107 30953
rect 9163 30897 9249 30953
rect 9305 30897 9391 30953
rect 9447 30897 9533 30953
rect 9589 30897 9675 30953
rect 9731 30897 9817 30953
rect 9873 30897 9959 30953
rect 10015 30897 10101 30953
rect 10157 30897 10243 30953
rect 10299 30897 10385 30953
rect 10441 30897 10527 30953
rect 10583 30897 10669 30953
rect 10725 30897 10811 30953
rect 10867 30897 10953 30953
rect 11009 30897 11095 30953
rect 11151 30897 11237 30953
rect 11293 30897 11379 30953
rect 11435 30897 11521 30953
rect 11577 30897 11663 30953
rect 11719 30897 11805 30953
rect 11861 30897 11947 30953
rect 12003 30897 12089 30953
rect 12145 30897 12231 30953
rect 12287 30897 12373 30953
rect 12429 30897 12515 30953
rect 12571 30897 12657 30953
rect 12713 30897 12799 30953
rect 12855 30897 12941 30953
rect 12997 30897 13083 30953
rect 13139 30897 13225 30953
rect 13281 30897 13367 30953
rect 13423 30897 13509 30953
rect 13565 30897 13651 30953
rect 13707 30897 13793 30953
rect 13849 30897 13935 30953
rect 13991 30897 14077 30953
rect 14133 30897 14219 30953
rect 14275 30897 14361 30953
rect 14417 30897 14503 30953
rect 14559 30897 14645 30953
rect 14701 30897 14787 30953
rect 14843 30897 14853 30953
rect 151 30811 14853 30897
rect 151 30755 161 30811
rect 217 30755 303 30811
rect 359 30755 445 30811
rect 501 30755 587 30811
rect 643 30755 729 30811
rect 785 30755 871 30811
rect 927 30755 1013 30811
rect 1069 30755 1155 30811
rect 1211 30755 1297 30811
rect 1353 30755 1439 30811
rect 1495 30755 1581 30811
rect 1637 30755 1723 30811
rect 1779 30755 1865 30811
rect 1921 30755 2007 30811
rect 2063 30755 2149 30811
rect 2205 30755 2291 30811
rect 2347 30755 2433 30811
rect 2489 30755 2575 30811
rect 2631 30755 2717 30811
rect 2773 30755 2859 30811
rect 2915 30755 3001 30811
rect 3057 30755 3143 30811
rect 3199 30755 3285 30811
rect 3341 30755 3427 30811
rect 3483 30755 3569 30811
rect 3625 30755 3711 30811
rect 3767 30755 3853 30811
rect 3909 30755 3995 30811
rect 4051 30755 4137 30811
rect 4193 30755 4279 30811
rect 4335 30755 4421 30811
rect 4477 30755 4563 30811
rect 4619 30755 4705 30811
rect 4761 30755 4847 30811
rect 4903 30755 4989 30811
rect 5045 30755 5131 30811
rect 5187 30755 5273 30811
rect 5329 30755 5415 30811
rect 5471 30755 5557 30811
rect 5613 30755 5699 30811
rect 5755 30755 5841 30811
rect 5897 30755 5983 30811
rect 6039 30755 6125 30811
rect 6181 30755 6267 30811
rect 6323 30755 6409 30811
rect 6465 30755 6551 30811
rect 6607 30755 6693 30811
rect 6749 30755 6835 30811
rect 6891 30755 6977 30811
rect 7033 30755 7119 30811
rect 7175 30755 7261 30811
rect 7317 30755 7403 30811
rect 7459 30755 7545 30811
rect 7601 30755 7687 30811
rect 7743 30755 7829 30811
rect 7885 30755 7971 30811
rect 8027 30755 8113 30811
rect 8169 30755 8255 30811
rect 8311 30755 8397 30811
rect 8453 30755 8539 30811
rect 8595 30755 8681 30811
rect 8737 30755 8823 30811
rect 8879 30755 8965 30811
rect 9021 30755 9107 30811
rect 9163 30755 9249 30811
rect 9305 30755 9391 30811
rect 9447 30755 9533 30811
rect 9589 30755 9675 30811
rect 9731 30755 9817 30811
rect 9873 30755 9959 30811
rect 10015 30755 10101 30811
rect 10157 30755 10243 30811
rect 10299 30755 10385 30811
rect 10441 30755 10527 30811
rect 10583 30755 10669 30811
rect 10725 30755 10811 30811
rect 10867 30755 10953 30811
rect 11009 30755 11095 30811
rect 11151 30755 11237 30811
rect 11293 30755 11379 30811
rect 11435 30755 11521 30811
rect 11577 30755 11663 30811
rect 11719 30755 11805 30811
rect 11861 30755 11947 30811
rect 12003 30755 12089 30811
rect 12145 30755 12231 30811
rect 12287 30755 12373 30811
rect 12429 30755 12515 30811
rect 12571 30755 12657 30811
rect 12713 30755 12799 30811
rect 12855 30755 12941 30811
rect 12997 30755 13083 30811
rect 13139 30755 13225 30811
rect 13281 30755 13367 30811
rect 13423 30755 13509 30811
rect 13565 30755 13651 30811
rect 13707 30755 13793 30811
rect 13849 30755 13935 30811
rect 13991 30755 14077 30811
rect 14133 30755 14219 30811
rect 14275 30755 14361 30811
rect 14417 30755 14503 30811
rect 14559 30755 14645 30811
rect 14701 30755 14787 30811
rect 14843 30755 14853 30811
rect 151 30669 14853 30755
rect 151 30613 161 30669
rect 217 30613 303 30669
rect 359 30613 445 30669
rect 501 30613 587 30669
rect 643 30613 729 30669
rect 785 30613 871 30669
rect 927 30613 1013 30669
rect 1069 30613 1155 30669
rect 1211 30613 1297 30669
rect 1353 30613 1439 30669
rect 1495 30613 1581 30669
rect 1637 30613 1723 30669
rect 1779 30613 1865 30669
rect 1921 30613 2007 30669
rect 2063 30613 2149 30669
rect 2205 30613 2291 30669
rect 2347 30613 2433 30669
rect 2489 30613 2575 30669
rect 2631 30613 2717 30669
rect 2773 30613 2859 30669
rect 2915 30613 3001 30669
rect 3057 30613 3143 30669
rect 3199 30613 3285 30669
rect 3341 30613 3427 30669
rect 3483 30613 3569 30669
rect 3625 30613 3711 30669
rect 3767 30613 3853 30669
rect 3909 30613 3995 30669
rect 4051 30613 4137 30669
rect 4193 30613 4279 30669
rect 4335 30613 4421 30669
rect 4477 30613 4563 30669
rect 4619 30613 4705 30669
rect 4761 30613 4847 30669
rect 4903 30613 4989 30669
rect 5045 30613 5131 30669
rect 5187 30613 5273 30669
rect 5329 30613 5415 30669
rect 5471 30613 5557 30669
rect 5613 30613 5699 30669
rect 5755 30613 5841 30669
rect 5897 30613 5983 30669
rect 6039 30613 6125 30669
rect 6181 30613 6267 30669
rect 6323 30613 6409 30669
rect 6465 30613 6551 30669
rect 6607 30613 6693 30669
rect 6749 30613 6835 30669
rect 6891 30613 6977 30669
rect 7033 30613 7119 30669
rect 7175 30613 7261 30669
rect 7317 30613 7403 30669
rect 7459 30613 7545 30669
rect 7601 30613 7687 30669
rect 7743 30613 7829 30669
rect 7885 30613 7971 30669
rect 8027 30613 8113 30669
rect 8169 30613 8255 30669
rect 8311 30613 8397 30669
rect 8453 30613 8539 30669
rect 8595 30613 8681 30669
rect 8737 30613 8823 30669
rect 8879 30613 8965 30669
rect 9021 30613 9107 30669
rect 9163 30613 9249 30669
rect 9305 30613 9391 30669
rect 9447 30613 9533 30669
rect 9589 30613 9675 30669
rect 9731 30613 9817 30669
rect 9873 30613 9959 30669
rect 10015 30613 10101 30669
rect 10157 30613 10243 30669
rect 10299 30613 10385 30669
rect 10441 30613 10527 30669
rect 10583 30613 10669 30669
rect 10725 30613 10811 30669
rect 10867 30613 10953 30669
rect 11009 30613 11095 30669
rect 11151 30613 11237 30669
rect 11293 30613 11379 30669
rect 11435 30613 11521 30669
rect 11577 30613 11663 30669
rect 11719 30613 11805 30669
rect 11861 30613 11947 30669
rect 12003 30613 12089 30669
rect 12145 30613 12231 30669
rect 12287 30613 12373 30669
rect 12429 30613 12515 30669
rect 12571 30613 12657 30669
rect 12713 30613 12799 30669
rect 12855 30613 12941 30669
rect 12997 30613 13083 30669
rect 13139 30613 13225 30669
rect 13281 30613 13367 30669
rect 13423 30613 13509 30669
rect 13565 30613 13651 30669
rect 13707 30613 13793 30669
rect 13849 30613 13935 30669
rect 13991 30613 14077 30669
rect 14133 30613 14219 30669
rect 14275 30613 14361 30669
rect 14417 30613 14503 30669
rect 14559 30613 14645 30669
rect 14701 30613 14787 30669
rect 14843 30613 14853 30669
rect 151 30527 14853 30613
rect 151 30471 161 30527
rect 217 30471 303 30527
rect 359 30471 445 30527
rect 501 30471 587 30527
rect 643 30471 729 30527
rect 785 30471 871 30527
rect 927 30471 1013 30527
rect 1069 30471 1155 30527
rect 1211 30471 1297 30527
rect 1353 30471 1439 30527
rect 1495 30471 1581 30527
rect 1637 30471 1723 30527
rect 1779 30471 1865 30527
rect 1921 30471 2007 30527
rect 2063 30471 2149 30527
rect 2205 30471 2291 30527
rect 2347 30471 2433 30527
rect 2489 30471 2575 30527
rect 2631 30471 2717 30527
rect 2773 30471 2859 30527
rect 2915 30471 3001 30527
rect 3057 30471 3143 30527
rect 3199 30471 3285 30527
rect 3341 30471 3427 30527
rect 3483 30471 3569 30527
rect 3625 30471 3711 30527
rect 3767 30471 3853 30527
rect 3909 30471 3995 30527
rect 4051 30471 4137 30527
rect 4193 30471 4279 30527
rect 4335 30471 4421 30527
rect 4477 30471 4563 30527
rect 4619 30471 4705 30527
rect 4761 30471 4847 30527
rect 4903 30471 4989 30527
rect 5045 30471 5131 30527
rect 5187 30471 5273 30527
rect 5329 30471 5415 30527
rect 5471 30471 5557 30527
rect 5613 30471 5699 30527
rect 5755 30471 5841 30527
rect 5897 30471 5983 30527
rect 6039 30471 6125 30527
rect 6181 30471 6267 30527
rect 6323 30471 6409 30527
rect 6465 30471 6551 30527
rect 6607 30471 6693 30527
rect 6749 30471 6835 30527
rect 6891 30471 6977 30527
rect 7033 30471 7119 30527
rect 7175 30471 7261 30527
rect 7317 30471 7403 30527
rect 7459 30471 7545 30527
rect 7601 30471 7687 30527
rect 7743 30471 7829 30527
rect 7885 30471 7971 30527
rect 8027 30471 8113 30527
rect 8169 30471 8255 30527
rect 8311 30471 8397 30527
rect 8453 30471 8539 30527
rect 8595 30471 8681 30527
rect 8737 30471 8823 30527
rect 8879 30471 8965 30527
rect 9021 30471 9107 30527
rect 9163 30471 9249 30527
rect 9305 30471 9391 30527
rect 9447 30471 9533 30527
rect 9589 30471 9675 30527
rect 9731 30471 9817 30527
rect 9873 30471 9959 30527
rect 10015 30471 10101 30527
rect 10157 30471 10243 30527
rect 10299 30471 10385 30527
rect 10441 30471 10527 30527
rect 10583 30471 10669 30527
rect 10725 30471 10811 30527
rect 10867 30471 10953 30527
rect 11009 30471 11095 30527
rect 11151 30471 11237 30527
rect 11293 30471 11379 30527
rect 11435 30471 11521 30527
rect 11577 30471 11663 30527
rect 11719 30471 11805 30527
rect 11861 30471 11947 30527
rect 12003 30471 12089 30527
rect 12145 30471 12231 30527
rect 12287 30471 12373 30527
rect 12429 30471 12515 30527
rect 12571 30471 12657 30527
rect 12713 30471 12799 30527
rect 12855 30471 12941 30527
rect 12997 30471 13083 30527
rect 13139 30471 13225 30527
rect 13281 30471 13367 30527
rect 13423 30471 13509 30527
rect 13565 30471 13651 30527
rect 13707 30471 13793 30527
rect 13849 30471 13935 30527
rect 13991 30471 14077 30527
rect 14133 30471 14219 30527
rect 14275 30471 14361 30527
rect 14417 30471 14503 30527
rect 14559 30471 14645 30527
rect 14701 30471 14787 30527
rect 14843 30471 14853 30527
rect 151 30385 14853 30471
rect 151 30329 161 30385
rect 217 30329 303 30385
rect 359 30329 445 30385
rect 501 30329 587 30385
rect 643 30329 729 30385
rect 785 30329 871 30385
rect 927 30329 1013 30385
rect 1069 30329 1155 30385
rect 1211 30329 1297 30385
rect 1353 30329 1439 30385
rect 1495 30329 1581 30385
rect 1637 30329 1723 30385
rect 1779 30329 1865 30385
rect 1921 30329 2007 30385
rect 2063 30329 2149 30385
rect 2205 30329 2291 30385
rect 2347 30329 2433 30385
rect 2489 30329 2575 30385
rect 2631 30329 2717 30385
rect 2773 30329 2859 30385
rect 2915 30329 3001 30385
rect 3057 30329 3143 30385
rect 3199 30329 3285 30385
rect 3341 30329 3427 30385
rect 3483 30329 3569 30385
rect 3625 30329 3711 30385
rect 3767 30329 3853 30385
rect 3909 30329 3995 30385
rect 4051 30329 4137 30385
rect 4193 30329 4279 30385
rect 4335 30329 4421 30385
rect 4477 30329 4563 30385
rect 4619 30329 4705 30385
rect 4761 30329 4847 30385
rect 4903 30329 4989 30385
rect 5045 30329 5131 30385
rect 5187 30329 5273 30385
rect 5329 30329 5415 30385
rect 5471 30329 5557 30385
rect 5613 30329 5699 30385
rect 5755 30329 5841 30385
rect 5897 30329 5983 30385
rect 6039 30329 6125 30385
rect 6181 30329 6267 30385
rect 6323 30329 6409 30385
rect 6465 30329 6551 30385
rect 6607 30329 6693 30385
rect 6749 30329 6835 30385
rect 6891 30329 6977 30385
rect 7033 30329 7119 30385
rect 7175 30329 7261 30385
rect 7317 30329 7403 30385
rect 7459 30329 7545 30385
rect 7601 30329 7687 30385
rect 7743 30329 7829 30385
rect 7885 30329 7971 30385
rect 8027 30329 8113 30385
rect 8169 30329 8255 30385
rect 8311 30329 8397 30385
rect 8453 30329 8539 30385
rect 8595 30329 8681 30385
rect 8737 30329 8823 30385
rect 8879 30329 8965 30385
rect 9021 30329 9107 30385
rect 9163 30329 9249 30385
rect 9305 30329 9391 30385
rect 9447 30329 9533 30385
rect 9589 30329 9675 30385
rect 9731 30329 9817 30385
rect 9873 30329 9959 30385
rect 10015 30329 10101 30385
rect 10157 30329 10243 30385
rect 10299 30329 10385 30385
rect 10441 30329 10527 30385
rect 10583 30329 10669 30385
rect 10725 30329 10811 30385
rect 10867 30329 10953 30385
rect 11009 30329 11095 30385
rect 11151 30329 11237 30385
rect 11293 30329 11379 30385
rect 11435 30329 11521 30385
rect 11577 30329 11663 30385
rect 11719 30329 11805 30385
rect 11861 30329 11947 30385
rect 12003 30329 12089 30385
rect 12145 30329 12231 30385
rect 12287 30329 12373 30385
rect 12429 30329 12515 30385
rect 12571 30329 12657 30385
rect 12713 30329 12799 30385
rect 12855 30329 12941 30385
rect 12997 30329 13083 30385
rect 13139 30329 13225 30385
rect 13281 30329 13367 30385
rect 13423 30329 13509 30385
rect 13565 30329 13651 30385
rect 13707 30329 13793 30385
rect 13849 30329 13935 30385
rect 13991 30329 14077 30385
rect 14133 30329 14219 30385
rect 14275 30329 14361 30385
rect 14417 30329 14503 30385
rect 14559 30329 14645 30385
rect 14701 30329 14787 30385
rect 14843 30329 14853 30385
rect 151 30243 14853 30329
rect 151 30187 161 30243
rect 217 30187 303 30243
rect 359 30187 445 30243
rect 501 30187 587 30243
rect 643 30187 729 30243
rect 785 30187 871 30243
rect 927 30187 1013 30243
rect 1069 30187 1155 30243
rect 1211 30187 1297 30243
rect 1353 30187 1439 30243
rect 1495 30187 1581 30243
rect 1637 30187 1723 30243
rect 1779 30187 1865 30243
rect 1921 30187 2007 30243
rect 2063 30187 2149 30243
rect 2205 30187 2291 30243
rect 2347 30187 2433 30243
rect 2489 30187 2575 30243
rect 2631 30187 2717 30243
rect 2773 30187 2859 30243
rect 2915 30187 3001 30243
rect 3057 30187 3143 30243
rect 3199 30187 3285 30243
rect 3341 30187 3427 30243
rect 3483 30187 3569 30243
rect 3625 30187 3711 30243
rect 3767 30187 3853 30243
rect 3909 30187 3995 30243
rect 4051 30187 4137 30243
rect 4193 30187 4279 30243
rect 4335 30187 4421 30243
rect 4477 30187 4563 30243
rect 4619 30187 4705 30243
rect 4761 30187 4847 30243
rect 4903 30187 4989 30243
rect 5045 30187 5131 30243
rect 5187 30187 5273 30243
rect 5329 30187 5415 30243
rect 5471 30187 5557 30243
rect 5613 30187 5699 30243
rect 5755 30187 5841 30243
rect 5897 30187 5983 30243
rect 6039 30187 6125 30243
rect 6181 30187 6267 30243
rect 6323 30187 6409 30243
rect 6465 30187 6551 30243
rect 6607 30187 6693 30243
rect 6749 30187 6835 30243
rect 6891 30187 6977 30243
rect 7033 30187 7119 30243
rect 7175 30187 7261 30243
rect 7317 30187 7403 30243
rect 7459 30187 7545 30243
rect 7601 30187 7687 30243
rect 7743 30187 7829 30243
rect 7885 30187 7971 30243
rect 8027 30187 8113 30243
rect 8169 30187 8255 30243
rect 8311 30187 8397 30243
rect 8453 30187 8539 30243
rect 8595 30187 8681 30243
rect 8737 30187 8823 30243
rect 8879 30187 8965 30243
rect 9021 30187 9107 30243
rect 9163 30187 9249 30243
rect 9305 30187 9391 30243
rect 9447 30187 9533 30243
rect 9589 30187 9675 30243
rect 9731 30187 9817 30243
rect 9873 30187 9959 30243
rect 10015 30187 10101 30243
rect 10157 30187 10243 30243
rect 10299 30187 10385 30243
rect 10441 30187 10527 30243
rect 10583 30187 10669 30243
rect 10725 30187 10811 30243
rect 10867 30187 10953 30243
rect 11009 30187 11095 30243
rect 11151 30187 11237 30243
rect 11293 30187 11379 30243
rect 11435 30187 11521 30243
rect 11577 30187 11663 30243
rect 11719 30187 11805 30243
rect 11861 30187 11947 30243
rect 12003 30187 12089 30243
rect 12145 30187 12231 30243
rect 12287 30187 12373 30243
rect 12429 30187 12515 30243
rect 12571 30187 12657 30243
rect 12713 30187 12799 30243
rect 12855 30187 12941 30243
rect 12997 30187 13083 30243
rect 13139 30187 13225 30243
rect 13281 30187 13367 30243
rect 13423 30187 13509 30243
rect 13565 30187 13651 30243
rect 13707 30187 13793 30243
rect 13849 30187 13935 30243
rect 13991 30187 14077 30243
rect 14133 30187 14219 30243
rect 14275 30187 14361 30243
rect 14417 30187 14503 30243
rect 14559 30187 14645 30243
rect 14701 30187 14787 30243
rect 14843 30187 14853 30243
rect 151 30101 14853 30187
rect 151 30045 161 30101
rect 217 30045 303 30101
rect 359 30045 445 30101
rect 501 30045 587 30101
rect 643 30045 729 30101
rect 785 30045 871 30101
rect 927 30045 1013 30101
rect 1069 30045 1155 30101
rect 1211 30045 1297 30101
rect 1353 30045 1439 30101
rect 1495 30045 1581 30101
rect 1637 30045 1723 30101
rect 1779 30045 1865 30101
rect 1921 30045 2007 30101
rect 2063 30045 2149 30101
rect 2205 30045 2291 30101
rect 2347 30045 2433 30101
rect 2489 30045 2575 30101
rect 2631 30045 2717 30101
rect 2773 30045 2859 30101
rect 2915 30045 3001 30101
rect 3057 30045 3143 30101
rect 3199 30045 3285 30101
rect 3341 30045 3427 30101
rect 3483 30045 3569 30101
rect 3625 30045 3711 30101
rect 3767 30045 3853 30101
rect 3909 30045 3995 30101
rect 4051 30045 4137 30101
rect 4193 30045 4279 30101
rect 4335 30045 4421 30101
rect 4477 30045 4563 30101
rect 4619 30045 4705 30101
rect 4761 30045 4847 30101
rect 4903 30045 4989 30101
rect 5045 30045 5131 30101
rect 5187 30045 5273 30101
rect 5329 30045 5415 30101
rect 5471 30045 5557 30101
rect 5613 30045 5699 30101
rect 5755 30045 5841 30101
rect 5897 30045 5983 30101
rect 6039 30045 6125 30101
rect 6181 30045 6267 30101
rect 6323 30045 6409 30101
rect 6465 30045 6551 30101
rect 6607 30045 6693 30101
rect 6749 30045 6835 30101
rect 6891 30045 6977 30101
rect 7033 30045 7119 30101
rect 7175 30045 7261 30101
rect 7317 30045 7403 30101
rect 7459 30045 7545 30101
rect 7601 30045 7687 30101
rect 7743 30045 7829 30101
rect 7885 30045 7971 30101
rect 8027 30045 8113 30101
rect 8169 30045 8255 30101
rect 8311 30045 8397 30101
rect 8453 30045 8539 30101
rect 8595 30045 8681 30101
rect 8737 30045 8823 30101
rect 8879 30045 8965 30101
rect 9021 30045 9107 30101
rect 9163 30045 9249 30101
rect 9305 30045 9391 30101
rect 9447 30045 9533 30101
rect 9589 30045 9675 30101
rect 9731 30045 9817 30101
rect 9873 30045 9959 30101
rect 10015 30045 10101 30101
rect 10157 30045 10243 30101
rect 10299 30045 10385 30101
rect 10441 30045 10527 30101
rect 10583 30045 10669 30101
rect 10725 30045 10811 30101
rect 10867 30045 10953 30101
rect 11009 30045 11095 30101
rect 11151 30045 11237 30101
rect 11293 30045 11379 30101
rect 11435 30045 11521 30101
rect 11577 30045 11663 30101
rect 11719 30045 11805 30101
rect 11861 30045 11947 30101
rect 12003 30045 12089 30101
rect 12145 30045 12231 30101
rect 12287 30045 12373 30101
rect 12429 30045 12515 30101
rect 12571 30045 12657 30101
rect 12713 30045 12799 30101
rect 12855 30045 12941 30101
rect 12997 30045 13083 30101
rect 13139 30045 13225 30101
rect 13281 30045 13367 30101
rect 13423 30045 13509 30101
rect 13565 30045 13651 30101
rect 13707 30045 13793 30101
rect 13849 30045 13935 30101
rect 13991 30045 14077 30101
rect 14133 30045 14219 30101
rect 14275 30045 14361 30101
rect 14417 30045 14503 30101
rect 14559 30045 14645 30101
rect 14701 30045 14787 30101
rect 14843 30045 14853 30101
rect 151 30035 14853 30045
rect 151 29741 14853 29751
rect 151 29685 161 29741
rect 217 29685 303 29741
rect 359 29685 445 29741
rect 501 29685 587 29741
rect 643 29685 729 29741
rect 785 29685 871 29741
rect 927 29685 1013 29741
rect 1069 29685 1155 29741
rect 1211 29685 1297 29741
rect 1353 29685 1439 29741
rect 1495 29685 1581 29741
rect 1637 29685 1723 29741
rect 1779 29685 1865 29741
rect 1921 29685 2007 29741
rect 2063 29685 2149 29741
rect 2205 29685 2291 29741
rect 2347 29685 2433 29741
rect 2489 29685 2575 29741
rect 2631 29685 2717 29741
rect 2773 29685 2859 29741
rect 2915 29685 3001 29741
rect 3057 29685 3143 29741
rect 3199 29685 3285 29741
rect 3341 29685 3427 29741
rect 3483 29685 3569 29741
rect 3625 29685 3711 29741
rect 3767 29685 3853 29741
rect 3909 29685 3995 29741
rect 4051 29685 4137 29741
rect 4193 29685 4279 29741
rect 4335 29685 4421 29741
rect 4477 29685 4563 29741
rect 4619 29685 4705 29741
rect 4761 29685 4847 29741
rect 4903 29685 4989 29741
rect 5045 29685 5131 29741
rect 5187 29685 5273 29741
rect 5329 29685 5415 29741
rect 5471 29685 5557 29741
rect 5613 29685 5699 29741
rect 5755 29685 5841 29741
rect 5897 29685 5983 29741
rect 6039 29685 6125 29741
rect 6181 29685 6267 29741
rect 6323 29685 6409 29741
rect 6465 29685 6551 29741
rect 6607 29685 6693 29741
rect 6749 29685 6835 29741
rect 6891 29685 6977 29741
rect 7033 29685 7119 29741
rect 7175 29685 7261 29741
rect 7317 29685 7403 29741
rect 7459 29685 7545 29741
rect 7601 29685 7687 29741
rect 7743 29685 7829 29741
rect 7885 29685 7971 29741
rect 8027 29685 8113 29741
rect 8169 29685 8255 29741
rect 8311 29685 8397 29741
rect 8453 29685 8539 29741
rect 8595 29685 8681 29741
rect 8737 29685 8823 29741
rect 8879 29685 8965 29741
rect 9021 29685 9107 29741
rect 9163 29685 9249 29741
rect 9305 29685 9391 29741
rect 9447 29685 9533 29741
rect 9589 29685 9675 29741
rect 9731 29685 9817 29741
rect 9873 29685 9959 29741
rect 10015 29685 10101 29741
rect 10157 29685 10243 29741
rect 10299 29685 10385 29741
rect 10441 29685 10527 29741
rect 10583 29685 10669 29741
rect 10725 29685 10811 29741
rect 10867 29685 10953 29741
rect 11009 29685 11095 29741
rect 11151 29685 11237 29741
rect 11293 29685 11379 29741
rect 11435 29685 11521 29741
rect 11577 29685 11663 29741
rect 11719 29685 11805 29741
rect 11861 29685 11947 29741
rect 12003 29685 12089 29741
rect 12145 29685 12231 29741
rect 12287 29685 12373 29741
rect 12429 29685 12515 29741
rect 12571 29685 12657 29741
rect 12713 29685 12799 29741
rect 12855 29685 12941 29741
rect 12997 29685 13083 29741
rect 13139 29685 13225 29741
rect 13281 29685 13367 29741
rect 13423 29685 13509 29741
rect 13565 29685 13651 29741
rect 13707 29685 13793 29741
rect 13849 29685 13935 29741
rect 13991 29685 14077 29741
rect 14133 29685 14219 29741
rect 14275 29685 14361 29741
rect 14417 29685 14503 29741
rect 14559 29685 14645 29741
rect 14701 29685 14787 29741
rect 14843 29685 14853 29741
rect 151 29599 14853 29685
rect 151 29543 161 29599
rect 217 29543 303 29599
rect 359 29543 445 29599
rect 501 29543 587 29599
rect 643 29543 729 29599
rect 785 29543 871 29599
rect 927 29543 1013 29599
rect 1069 29543 1155 29599
rect 1211 29543 1297 29599
rect 1353 29543 1439 29599
rect 1495 29543 1581 29599
rect 1637 29543 1723 29599
rect 1779 29543 1865 29599
rect 1921 29543 2007 29599
rect 2063 29543 2149 29599
rect 2205 29543 2291 29599
rect 2347 29543 2433 29599
rect 2489 29543 2575 29599
rect 2631 29543 2717 29599
rect 2773 29543 2859 29599
rect 2915 29543 3001 29599
rect 3057 29543 3143 29599
rect 3199 29543 3285 29599
rect 3341 29543 3427 29599
rect 3483 29543 3569 29599
rect 3625 29543 3711 29599
rect 3767 29543 3853 29599
rect 3909 29543 3995 29599
rect 4051 29543 4137 29599
rect 4193 29543 4279 29599
rect 4335 29543 4421 29599
rect 4477 29543 4563 29599
rect 4619 29543 4705 29599
rect 4761 29543 4847 29599
rect 4903 29543 4989 29599
rect 5045 29543 5131 29599
rect 5187 29543 5273 29599
rect 5329 29543 5415 29599
rect 5471 29543 5557 29599
rect 5613 29543 5699 29599
rect 5755 29543 5841 29599
rect 5897 29543 5983 29599
rect 6039 29543 6125 29599
rect 6181 29543 6267 29599
rect 6323 29543 6409 29599
rect 6465 29543 6551 29599
rect 6607 29543 6693 29599
rect 6749 29543 6835 29599
rect 6891 29543 6977 29599
rect 7033 29543 7119 29599
rect 7175 29543 7261 29599
rect 7317 29543 7403 29599
rect 7459 29543 7545 29599
rect 7601 29543 7687 29599
rect 7743 29543 7829 29599
rect 7885 29543 7971 29599
rect 8027 29543 8113 29599
rect 8169 29543 8255 29599
rect 8311 29543 8397 29599
rect 8453 29543 8539 29599
rect 8595 29543 8681 29599
rect 8737 29543 8823 29599
rect 8879 29543 8965 29599
rect 9021 29543 9107 29599
rect 9163 29543 9249 29599
rect 9305 29543 9391 29599
rect 9447 29543 9533 29599
rect 9589 29543 9675 29599
rect 9731 29543 9817 29599
rect 9873 29543 9959 29599
rect 10015 29543 10101 29599
rect 10157 29543 10243 29599
rect 10299 29543 10385 29599
rect 10441 29543 10527 29599
rect 10583 29543 10669 29599
rect 10725 29543 10811 29599
rect 10867 29543 10953 29599
rect 11009 29543 11095 29599
rect 11151 29543 11237 29599
rect 11293 29543 11379 29599
rect 11435 29543 11521 29599
rect 11577 29543 11663 29599
rect 11719 29543 11805 29599
rect 11861 29543 11947 29599
rect 12003 29543 12089 29599
rect 12145 29543 12231 29599
rect 12287 29543 12373 29599
rect 12429 29543 12515 29599
rect 12571 29543 12657 29599
rect 12713 29543 12799 29599
rect 12855 29543 12941 29599
rect 12997 29543 13083 29599
rect 13139 29543 13225 29599
rect 13281 29543 13367 29599
rect 13423 29543 13509 29599
rect 13565 29543 13651 29599
rect 13707 29543 13793 29599
rect 13849 29543 13935 29599
rect 13991 29543 14077 29599
rect 14133 29543 14219 29599
rect 14275 29543 14361 29599
rect 14417 29543 14503 29599
rect 14559 29543 14645 29599
rect 14701 29543 14787 29599
rect 14843 29543 14853 29599
rect 151 29457 14853 29543
rect 151 29401 161 29457
rect 217 29401 303 29457
rect 359 29401 445 29457
rect 501 29401 587 29457
rect 643 29401 729 29457
rect 785 29401 871 29457
rect 927 29401 1013 29457
rect 1069 29401 1155 29457
rect 1211 29401 1297 29457
rect 1353 29401 1439 29457
rect 1495 29401 1581 29457
rect 1637 29401 1723 29457
rect 1779 29401 1865 29457
rect 1921 29401 2007 29457
rect 2063 29401 2149 29457
rect 2205 29401 2291 29457
rect 2347 29401 2433 29457
rect 2489 29401 2575 29457
rect 2631 29401 2717 29457
rect 2773 29401 2859 29457
rect 2915 29401 3001 29457
rect 3057 29401 3143 29457
rect 3199 29401 3285 29457
rect 3341 29401 3427 29457
rect 3483 29401 3569 29457
rect 3625 29401 3711 29457
rect 3767 29401 3853 29457
rect 3909 29401 3995 29457
rect 4051 29401 4137 29457
rect 4193 29401 4279 29457
rect 4335 29401 4421 29457
rect 4477 29401 4563 29457
rect 4619 29401 4705 29457
rect 4761 29401 4847 29457
rect 4903 29401 4989 29457
rect 5045 29401 5131 29457
rect 5187 29401 5273 29457
rect 5329 29401 5415 29457
rect 5471 29401 5557 29457
rect 5613 29401 5699 29457
rect 5755 29401 5841 29457
rect 5897 29401 5983 29457
rect 6039 29401 6125 29457
rect 6181 29401 6267 29457
rect 6323 29401 6409 29457
rect 6465 29401 6551 29457
rect 6607 29401 6693 29457
rect 6749 29401 6835 29457
rect 6891 29401 6977 29457
rect 7033 29401 7119 29457
rect 7175 29401 7261 29457
rect 7317 29401 7403 29457
rect 7459 29401 7545 29457
rect 7601 29401 7687 29457
rect 7743 29401 7829 29457
rect 7885 29401 7971 29457
rect 8027 29401 8113 29457
rect 8169 29401 8255 29457
rect 8311 29401 8397 29457
rect 8453 29401 8539 29457
rect 8595 29401 8681 29457
rect 8737 29401 8823 29457
rect 8879 29401 8965 29457
rect 9021 29401 9107 29457
rect 9163 29401 9249 29457
rect 9305 29401 9391 29457
rect 9447 29401 9533 29457
rect 9589 29401 9675 29457
rect 9731 29401 9817 29457
rect 9873 29401 9959 29457
rect 10015 29401 10101 29457
rect 10157 29401 10243 29457
rect 10299 29401 10385 29457
rect 10441 29401 10527 29457
rect 10583 29401 10669 29457
rect 10725 29401 10811 29457
rect 10867 29401 10953 29457
rect 11009 29401 11095 29457
rect 11151 29401 11237 29457
rect 11293 29401 11379 29457
rect 11435 29401 11521 29457
rect 11577 29401 11663 29457
rect 11719 29401 11805 29457
rect 11861 29401 11947 29457
rect 12003 29401 12089 29457
rect 12145 29401 12231 29457
rect 12287 29401 12373 29457
rect 12429 29401 12515 29457
rect 12571 29401 12657 29457
rect 12713 29401 12799 29457
rect 12855 29401 12941 29457
rect 12997 29401 13083 29457
rect 13139 29401 13225 29457
rect 13281 29401 13367 29457
rect 13423 29401 13509 29457
rect 13565 29401 13651 29457
rect 13707 29401 13793 29457
rect 13849 29401 13935 29457
rect 13991 29401 14077 29457
rect 14133 29401 14219 29457
rect 14275 29401 14361 29457
rect 14417 29401 14503 29457
rect 14559 29401 14645 29457
rect 14701 29401 14787 29457
rect 14843 29401 14853 29457
rect 151 29315 14853 29401
rect 151 29259 161 29315
rect 217 29259 303 29315
rect 359 29259 445 29315
rect 501 29259 587 29315
rect 643 29259 729 29315
rect 785 29259 871 29315
rect 927 29259 1013 29315
rect 1069 29259 1155 29315
rect 1211 29259 1297 29315
rect 1353 29259 1439 29315
rect 1495 29259 1581 29315
rect 1637 29259 1723 29315
rect 1779 29259 1865 29315
rect 1921 29259 2007 29315
rect 2063 29259 2149 29315
rect 2205 29259 2291 29315
rect 2347 29259 2433 29315
rect 2489 29259 2575 29315
rect 2631 29259 2717 29315
rect 2773 29259 2859 29315
rect 2915 29259 3001 29315
rect 3057 29259 3143 29315
rect 3199 29259 3285 29315
rect 3341 29259 3427 29315
rect 3483 29259 3569 29315
rect 3625 29259 3711 29315
rect 3767 29259 3853 29315
rect 3909 29259 3995 29315
rect 4051 29259 4137 29315
rect 4193 29259 4279 29315
rect 4335 29259 4421 29315
rect 4477 29259 4563 29315
rect 4619 29259 4705 29315
rect 4761 29259 4847 29315
rect 4903 29259 4989 29315
rect 5045 29259 5131 29315
rect 5187 29259 5273 29315
rect 5329 29259 5415 29315
rect 5471 29259 5557 29315
rect 5613 29259 5699 29315
rect 5755 29259 5841 29315
rect 5897 29259 5983 29315
rect 6039 29259 6125 29315
rect 6181 29259 6267 29315
rect 6323 29259 6409 29315
rect 6465 29259 6551 29315
rect 6607 29259 6693 29315
rect 6749 29259 6835 29315
rect 6891 29259 6977 29315
rect 7033 29259 7119 29315
rect 7175 29259 7261 29315
rect 7317 29259 7403 29315
rect 7459 29259 7545 29315
rect 7601 29259 7687 29315
rect 7743 29259 7829 29315
rect 7885 29259 7971 29315
rect 8027 29259 8113 29315
rect 8169 29259 8255 29315
rect 8311 29259 8397 29315
rect 8453 29259 8539 29315
rect 8595 29259 8681 29315
rect 8737 29259 8823 29315
rect 8879 29259 8965 29315
rect 9021 29259 9107 29315
rect 9163 29259 9249 29315
rect 9305 29259 9391 29315
rect 9447 29259 9533 29315
rect 9589 29259 9675 29315
rect 9731 29259 9817 29315
rect 9873 29259 9959 29315
rect 10015 29259 10101 29315
rect 10157 29259 10243 29315
rect 10299 29259 10385 29315
rect 10441 29259 10527 29315
rect 10583 29259 10669 29315
rect 10725 29259 10811 29315
rect 10867 29259 10953 29315
rect 11009 29259 11095 29315
rect 11151 29259 11237 29315
rect 11293 29259 11379 29315
rect 11435 29259 11521 29315
rect 11577 29259 11663 29315
rect 11719 29259 11805 29315
rect 11861 29259 11947 29315
rect 12003 29259 12089 29315
rect 12145 29259 12231 29315
rect 12287 29259 12373 29315
rect 12429 29259 12515 29315
rect 12571 29259 12657 29315
rect 12713 29259 12799 29315
rect 12855 29259 12941 29315
rect 12997 29259 13083 29315
rect 13139 29259 13225 29315
rect 13281 29259 13367 29315
rect 13423 29259 13509 29315
rect 13565 29259 13651 29315
rect 13707 29259 13793 29315
rect 13849 29259 13935 29315
rect 13991 29259 14077 29315
rect 14133 29259 14219 29315
rect 14275 29259 14361 29315
rect 14417 29259 14503 29315
rect 14559 29259 14645 29315
rect 14701 29259 14787 29315
rect 14843 29259 14853 29315
rect 151 29173 14853 29259
rect 151 29117 161 29173
rect 217 29117 303 29173
rect 359 29117 445 29173
rect 501 29117 587 29173
rect 643 29117 729 29173
rect 785 29117 871 29173
rect 927 29117 1013 29173
rect 1069 29117 1155 29173
rect 1211 29117 1297 29173
rect 1353 29117 1439 29173
rect 1495 29117 1581 29173
rect 1637 29117 1723 29173
rect 1779 29117 1865 29173
rect 1921 29117 2007 29173
rect 2063 29117 2149 29173
rect 2205 29117 2291 29173
rect 2347 29117 2433 29173
rect 2489 29117 2575 29173
rect 2631 29117 2717 29173
rect 2773 29117 2859 29173
rect 2915 29117 3001 29173
rect 3057 29117 3143 29173
rect 3199 29117 3285 29173
rect 3341 29117 3427 29173
rect 3483 29117 3569 29173
rect 3625 29117 3711 29173
rect 3767 29117 3853 29173
rect 3909 29117 3995 29173
rect 4051 29117 4137 29173
rect 4193 29117 4279 29173
rect 4335 29117 4421 29173
rect 4477 29117 4563 29173
rect 4619 29117 4705 29173
rect 4761 29117 4847 29173
rect 4903 29117 4989 29173
rect 5045 29117 5131 29173
rect 5187 29117 5273 29173
rect 5329 29117 5415 29173
rect 5471 29117 5557 29173
rect 5613 29117 5699 29173
rect 5755 29117 5841 29173
rect 5897 29117 5983 29173
rect 6039 29117 6125 29173
rect 6181 29117 6267 29173
rect 6323 29117 6409 29173
rect 6465 29117 6551 29173
rect 6607 29117 6693 29173
rect 6749 29117 6835 29173
rect 6891 29117 6977 29173
rect 7033 29117 7119 29173
rect 7175 29117 7261 29173
rect 7317 29117 7403 29173
rect 7459 29117 7545 29173
rect 7601 29117 7687 29173
rect 7743 29117 7829 29173
rect 7885 29117 7971 29173
rect 8027 29117 8113 29173
rect 8169 29117 8255 29173
rect 8311 29117 8397 29173
rect 8453 29117 8539 29173
rect 8595 29117 8681 29173
rect 8737 29117 8823 29173
rect 8879 29117 8965 29173
rect 9021 29117 9107 29173
rect 9163 29117 9249 29173
rect 9305 29117 9391 29173
rect 9447 29117 9533 29173
rect 9589 29117 9675 29173
rect 9731 29117 9817 29173
rect 9873 29117 9959 29173
rect 10015 29117 10101 29173
rect 10157 29117 10243 29173
rect 10299 29117 10385 29173
rect 10441 29117 10527 29173
rect 10583 29117 10669 29173
rect 10725 29117 10811 29173
rect 10867 29117 10953 29173
rect 11009 29117 11095 29173
rect 11151 29117 11237 29173
rect 11293 29117 11379 29173
rect 11435 29117 11521 29173
rect 11577 29117 11663 29173
rect 11719 29117 11805 29173
rect 11861 29117 11947 29173
rect 12003 29117 12089 29173
rect 12145 29117 12231 29173
rect 12287 29117 12373 29173
rect 12429 29117 12515 29173
rect 12571 29117 12657 29173
rect 12713 29117 12799 29173
rect 12855 29117 12941 29173
rect 12997 29117 13083 29173
rect 13139 29117 13225 29173
rect 13281 29117 13367 29173
rect 13423 29117 13509 29173
rect 13565 29117 13651 29173
rect 13707 29117 13793 29173
rect 13849 29117 13935 29173
rect 13991 29117 14077 29173
rect 14133 29117 14219 29173
rect 14275 29117 14361 29173
rect 14417 29117 14503 29173
rect 14559 29117 14645 29173
rect 14701 29117 14787 29173
rect 14843 29117 14853 29173
rect 151 29031 14853 29117
rect 151 28975 161 29031
rect 217 28975 303 29031
rect 359 28975 445 29031
rect 501 28975 587 29031
rect 643 28975 729 29031
rect 785 28975 871 29031
rect 927 28975 1013 29031
rect 1069 28975 1155 29031
rect 1211 28975 1297 29031
rect 1353 28975 1439 29031
rect 1495 28975 1581 29031
rect 1637 28975 1723 29031
rect 1779 28975 1865 29031
rect 1921 28975 2007 29031
rect 2063 28975 2149 29031
rect 2205 28975 2291 29031
rect 2347 28975 2433 29031
rect 2489 28975 2575 29031
rect 2631 28975 2717 29031
rect 2773 28975 2859 29031
rect 2915 28975 3001 29031
rect 3057 28975 3143 29031
rect 3199 28975 3285 29031
rect 3341 28975 3427 29031
rect 3483 28975 3569 29031
rect 3625 28975 3711 29031
rect 3767 28975 3853 29031
rect 3909 28975 3995 29031
rect 4051 28975 4137 29031
rect 4193 28975 4279 29031
rect 4335 28975 4421 29031
rect 4477 28975 4563 29031
rect 4619 28975 4705 29031
rect 4761 28975 4847 29031
rect 4903 28975 4989 29031
rect 5045 28975 5131 29031
rect 5187 28975 5273 29031
rect 5329 28975 5415 29031
rect 5471 28975 5557 29031
rect 5613 28975 5699 29031
rect 5755 28975 5841 29031
rect 5897 28975 5983 29031
rect 6039 28975 6125 29031
rect 6181 28975 6267 29031
rect 6323 28975 6409 29031
rect 6465 28975 6551 29031
rect 6607 28975 6693 29031
rect 6749 28975 6835 29031
rect 6891 28975 6977 29031
rect 7033 28975 7119 29031
rect 7175 28975 7261 29031
rect 7317 28975 7403 29031
rect 7459 28975 7545 29031
rect 7601 28975 7687 29031
rect 7743 28975 7829 29031
rect 7885 28975 7971 29031
rect 8027 28975 8113 29031
rect 8169 28975 8255 29031
rect 8311 28975 8397 29031
rect 8453 28975 8539 29031
rect 8595 28975 8681 29031
rect 8737 28975 8823 29031
rect 8879 28975 8965 29031
rect 9021 28975 9107 29031
rect 9163 28975 9249 29031
rect 9305 28975 9391 29031
rect 9447 28975 9533 29031
rect 9589 28975 9675 29031
rect 9731 28975 9817 29031
rect 9873 28975 9959 29031
rect 10015 28975 10101 29031
rect 10157 28975 10243 29031
rect 10299 28975 10385 29031
rect 10441 28975 10527 29031
rect 10583 28975 10669 29031
rect 10725 28975 10811 29031
rect 10867 28975 10953 29031
rect 11009 28975 11095 29031
rect 11151 28975 11237 29031
rect 11293 28975 11379 29031
rect 11435 28975 11521 29031
rect 11577 28975 11663 29031
rect 11719 28975 11805 29031
rect 11861 28975 11947 29031
rect 12003 28975 12089 29031
rect 12145 28975 12231 29031
rect 12287 28975 12373 29031
rect 12429 28975 12515 29031
rect 12571 28975 12657 29031
rect 12713 28975 12799 29031
rect 12855 28975 12941 29031
rect 12997 28975 13083 29031
rect 13139 28975 13225 29031
rect 13281 28975 13367 29031
rect 13423 28975 13509 29031
rect 13565 28975 13651 29031
rect 13707 28975 13793 29031
rect 13849 28975 13935 29031
rect 13991 28975 14077 29031
rect 14133 28975 14219 29031
rect 14275 28975 14361 29031
rect 14417 28975 14503 29031
rect 14559 28975 14645 29031
rect 14701 28975 14787 29031
rect 14843 28975 14853 29031
rect 151 28889 14853 28975
rect 151 28833 161 28889
rect 217 28833 303 28889
rect 359 28833 445 28889
rect 501 28833 587 28889
rect 643 28833 729 28889
rect 785 28833 871 28889
rect 927 28833 1013 28889
rect 1069 28833 1155 28889
rect 1211 28833 1297 28889
rect 1353 28833 1439 28889
rect 1495 28833 1581 28889
rect 1637 28833 1723 28889
rect 1779 28833 1865 28889
rect 1921 28833 2007 28889
rect 2063 28833 2149 28889
rect 2205 28833 2291 28889
rect 2347 28833 2433 28889
rect 2489 28833 2575 28889
rect 2631 28833 2717 28889
rect 2773 28833 2859 28889
rect 2915 28833 3001 28889
rect 3057 28833 3143 28889
rect 3199 28833 3285 28889
rect 3341 28833 3427 28889
rect 3483 28833 3569 28889
rect 3625 28833 3711 28889
rect 3767 28833 3853 28889
rect 3909 28833 3995 28889
rect 4051 28833 4137 28889
rect 4193 28833 4279 28889
rect 4335 28833 4421 28889
rect 4477 28833 4563 28889
rect 4619 28833 4705 28889
rect 4761 28833 4847 28889
rect 4903 28833 4989 28889
rect 5045 28833 5131 28889
rect 5187 28833 5273 28889
rect 5329 28833 5415 28889
rect 5471 28833 5557 28889
rect 5613 28833 5699 28889
rect 5755 28833 5841 28889
rect 5897 28833 5983 28889
rect 6039 28833 6125 28889
rect 6181 28833 6267 28889
rect 6323 28833 6409 28889
rect 6465 28833 6551 28889
rect 6607 28833 6693 28889
rect 6749 28833 6835 28889
rect 6891 28833 6977 28889
rect 7033 28833 7119 28889
rect 7175 28833 7261 28889
rect 7317 28833 7403 28889
rect 7459 28833 7545 28889
rect 7601 28833 7687 28889
rect 7743 28833 7829 28889
rect 7885 28833 7971 28889
rect 8027 28833 8113 28889
rect 8169 28833 8255 28889
rect 8311 28833 8397 28889
rect 8453 28833 8539 28889
rect 8595 28833 8681 28889
rect 8737 28833 8823 28889
rect 8879 28833 8965 28889
rect 9021 28833 9107 28889
rect 9163 28833 9249 28889
rect 9305 28833 9391 28889
rect 9447 28833 9533 28889
rect 9589 28833 9675 28889
rect 9731 28833 9817 28889
rect 9873 28833 9959 28889
rect 10015 28833 10101 28889
rect 10157 28833 10243 28889
rect 10299 28833 10385 28889
rect 10441 28833 10527 28889
rect 10583 28833 10669 28889
rect 10725 28833 10811 28889
rect 10867 28833 10953 28889
rect 11009 28833 11095 28889
rect 11151 28833 11237 28889
rect 11293 28833 11379 28889
rect 11435 28833 11521 28889
rect 11577 28833 11663 28889
rect 11719 28833 11805 28889
rect 11861 28833 11947 28889
rect 12003 28833 12089 28889
rect 12145 28833 12231 28889
rect 12287 28833 12373 28889
rect 12429 28833 12515 28889
rect 12571 28833 12657 28889
rect 12713 28833 12799 28889
rect 12855 28833 12941 28889
rect 12997 28833 13083 28889
rect 13139 28833 13225 28889
rect 13281 28833 13367 28889
rect 13423 28833 13509 28889
rect 13565 28833 13651 28889
rect 13707 28833 13793 28889
rect 13849 28833 13935 28889
rect 13991 28833 14077 28889
rect 14133 28833 14219 28889
rect 14275 28833 14361 28889
rect 14417 28833 14503 28889
rect 14559 28833 14645 28889
rect 14701 28833 14787 28889
rect 14843 28833 14853 28889
rect 151 28747 14853 28833
rect 151 28691 161 28747
rect 217 28691 303 28747
rect 359 28691 445 28747
rect 501 28691 587 28747
rect 643 28691 729 28747
rect 785 28691 871 28747
rect 927 28691 1013 28747
rect 1069 28691 1155 28747
rect 1211 28691 1297 28747
rect 1353 28691 1439 28747
rect 1495 28691 1581 28747
rect 1637 28691 1723 28747
rect 1779 28691 1865 28747
rect 1921 28691 2007 28747
rect 2063 28691 2149 28747
rect 2205 28691 2291 28747
rect 2347 28691 2433 28747
rect 2489 28691 2575 28747
rect 2631 28691 2717 28747
rect 2773 28691 2859 28747
rect 2915 28691 3001 28747
rect 3057 28691 3143 28747
rect 3199 28691 3285 28747
rect 3341 28691 3427 28747
rect 3483 28691 3569 28747
rect 3625 28691 3711 28747
rect 3767 28691 3853 28747
rect 3909 28691 3995 28747
rect 4051 28691 4137 28747
rect 4193 28691 4279 28747
rect 4335 28691 4421 28747
rect 4477 28691 4563 28747
rect 4619 28691 4705 28747
rect 4761 28691 4847 28747
rect 4903 28691 4989 28747
rect 5045 28691 5131 28747
rect 5187 28691 5273 28747
rect 5329 28691 5415 28747
rect 5471 28691 5557 28747
rect 5613 28691 5699 28747
rect 5755 28691 5841 28747
rect 5897 28691 5983 28747
rect 6039 28691 6125 28747
rect 6181 28691 6267 28747
rect 6323 28691 6409 28747
rect 6465 28691 6551 28747
rect 6607 28691 6693 28747
rect 6749 28691 6835 28747
rect 6891 28691 6977 28747
rect 7033 28691 7119 28747
rect 7175 28691 7261 28747
rect 7317 28691 7403 28747
rect 7459 28691 7545 28747
rect 7601 28691 7687 28747
rect 7743 28691 7829 28747
rect 7885 28691 7971 28747
rect 8027 28691 8113 28747
rect 8169 28691 8255 28747
rect 8311 28691 8397 28747
rect 8453 28691 8539 28747
rect 8595 28691 8681 28747
rect 8737 28691 8823 28747
rect 8879 28691 8965 28747
rect 9021 28691 9107 28747
rect 9163 28691 9249 28747
rect 9305 28691 9391 28747
rect 9447 28691 9533 28747
rect 9589 28691 9675 28747
rect 9731 28691 9817 28747
rect 9873 28691 9959 28747
rect 10015 28691 10101 28747
rect 10157 28691 10243 28747
rect 10299 28691 10385 28747
rect 10441 28691 10527 28747
rect 10583 28691 10669 28747
rect 10725 28691 10811 28747
rect 10867 28691 10953 28747
rect 11009 28691 11095 28747
rect 11151 28691 11237 28747
rect 11293 28691 11379 28747
rect 11435 28691 11521 28747
rect 11577 28691 11663 28747
rect 11719 28691 11805 28747
rect 11861 28691 11947 28747
rect 12003 28691 12089 28747
rect 12145 28691 12231 28747
rect 12287 28691 12373 28747
rect 12429 28691 12515 28747
rect 12571 28691 12657 28747
rect 12713 28691 12799 28747
rect 12855 28691 12941 28747
rect 12997 28691 13083 28747
rect 13139 28691 13225 28747
rect 13281 28691 13367 28747
rect 13423 28691 13509 28747
rect 13565 28691 13651 28747
rect 13707 28691 13793 28747
rect 13849 28691 13935 28747
rect 13991 28691 14077 28747
rect 14133 28691 14219 28747
rect 14275 28691 14361 28747
rect 14417 28691 14503 28747
rect 14559 28691 14645 28747
rect 14701 28691 14787 28747
rect 14843 28691 14853 28747
rect 151 28605 14853 28691
rect 151 28549 161 28605
rect 217 28549 303 28605
rect 359 28549 445 28605
rect 501 28549 587 28605
rect 643 28549 729 28605
rect 785 28549 871 28605
rect 927 28549 1013 28605
rect 1069 28549 1155 28605
rect 1211 28549 1297 28605
rect 1353 28549 1439 28605
rect 1495 28549 1581 28605
rect 1637 28549 1723 28605
rect 1779 28549 1865 28605
rect 1921 28549 2007 28605
rect 2063 28549 2149 28605
rect 2205 28549 2291 28605
rect 2347 28549 2433 28605
rect 2489 28549 2575 28605
rect 2631 28549 2717 28605
rect 2773 28549 2859 28605
rect 2915 28549 3001 28605
rect 3057 28549 3143 28605
rect 3199 28549 3285 28605
rect 3341 28549 3427 28605
rect 3483 28549 3569 28605
rect 3625 28549 3711 28605
rect 3767 28549 3853 28605
rect 3909 28549 3995 28605
rect 4051 28549 4137 28605
rect 4193 28549 4279 28605
rect 4335 28549 4421 28605
rect 4477 28549 4563 28605
rect 4619 28549 4705 28605
rect 4761 28549 4847 28605
rect 4903 28549 4989 28605
rect 5045 28549 5131 28605
rect 5187 28549 5273 28605
rect 5329 28549 5415 28605
rect 5471 28549 5557 28605
rect 5613 28549 5699 28605
rect 5755 28549 5841 28605
rect 5897 28549 5983 28605
rect 6039 28549 6125 28605
rect 6181 28549 6267 28605
rect 6323 28549 6409 28605
rect 6465 28549 6551 28605
rect 6607 28549 6693 28605
rect 6749 28549 6835 28605
rect 6891 28549 6977 28605
rect 7033 28549 7119 28605
rect 7175 28549 7261 28605
rect 7317 28549 7403 28605
rect 7459 28549 7545 28605
rect 7601 28549 7687 28605
rect 7743 28549 7829 28605
rect 7885 28549 7971 28605
rect 8027 28549 8113 28605
rect 8169 28549 8255 28605
rect 8311 28549 8397 28605
rect 8453 28549 8539 28605
rect 8595 28549 8681 28605
rect 8737 28549 8823 28605
rect 8879 28549 8965 28605
rect 9021 28549 9107 28605
rect 9163 28549 9249 28605
rect 9305 28549 9391 28605
rect 9447 28549 9533 28605
rect 9589 28549 9675 28605
rect 9731 28549 9817 28605
rect 9873 28549 9959 28605
rect 10015 28549 10101 28605
rect 10157 28549 10243 28605
rect 10299 28549 10385 28605
rect 10441 28549 10527 28605
rect 10583 28549 10669 28605
rect 10725 28549 10811 28605
rect 10867 28549 10953 28605
rect 11009 28549 11095 28605
rect 11151 28549 11237 28605
rect 11293 28549 11379 28605
rect 11435 28549 11521 28605
rect 11577 28549 11663 28605
rect 11719 28549 11805 28605
rect 11861 28549 11947 28605
rect 12003 28549 12089 28605
rect 12145 28549 12231 28605
rect 12287 28549 12373 28605
rect 12429 28549 12515 28605
rect 12571 28549 12657 28605
rect 12713 28549 12799 28605
rect 12855 28549 12941 28605
rect 12997 28549 13083 28605
rect 13139 28549 13225 28605
rect 13281 28549 13367 28605
rect 13423 28549 13509 28605
rect 13565 28549 13651 28605
rect 13707 28549 13793 28605
rect 13849 28549 13935 28605
rect 13991 28549 14077 28605
rect 14133 28549 14219 28605
rect 14275 28549 14361 28605
rect 14417 28549 14503 28605
rect 14559 28549 14645 28605
rect 14701 28549 14787 28605
rect 14843 28549 14853 28605
rect 151 28463 14853 28549
rect 151 28407 161 28463
rect 217 28407 303 28463
rect 359 28407 445 28463
rect 501 28407 587 28463
rect 643 28407 729 28463
rect 785 28407 871 28463
rect 927 28407 1013 28463
rect 1069 28407 1155 28463
rect 1211 28407 1297 28463
rect 1353 28407 1439 28463
rect 1495 28407 1581 28463
rect 1637 28407 1723 28463
rect 1779 28407 1865 28463
rect 1921 28407 2007 28463
rect 2063 28407 2149 28463
rect 2205 28407 2291 28463
rect 2347 28407 2433 28463
rect 2489 28407 2575 28463
rect 2631 28407 2717 28463
rect 2773 28407 2859 28463
rect 2915 28407 3001 28463
rect 3057 28407 3143 28463
rect 3199 28407 3285 28463
rect 3341 28407 3427 28463
rect 3483 28407 3569 28463
rect 3625 28407 3711 28463
rect 3767 28407 3853 28463
rect 3909 28407 3995 28463
rect 4051 28407 4137 28463
rect 4193 28407 4279 28463
rect 4335 28407 4421 28463
rect 4477 28407 4563 28463
rect 4619 28407 4705 28463
rect 4761 28407 4847 28463
rect 4903 28407 4989 28463
rect 5045 28407 5131 28463
rect 5187 28407 5273 28463
rect 5329 28407 5415 28463
rect 5471 28407 5557 28463
rect 5613 28407 5699 28463
rect 5755 28407 5841 28463
rect 5897 28407 5983 28463
rect 6039 28407 6125 28463
rect 6181 28407 6267 28463
rect 6323 28407 6409 28463
rect 6465 28407 6551 28463
rect 6607 28407 6693 28463
rect 6749 28407 6835 28463
rect 6891 28407 6977 28463
rect 7033 28407 7119 28463
rect 7175 28407 7261 28463
rect 7317 28407 7403 28463
rect 7459 28407 7545 28463
rect 7601 28407 7687 28463
rect 7743 28407 7829 28463
rect 7885 28407 7971 28463
rect 8027 28407 8113 28463
rect 8169 28407 8255 28463
rect 8311 28407 8397 28463
rect 8453 28407 8539 28463
rect 8595 28407 8681 28463
rect 8737 28407 8823 28463
rect 8879 28407 8965 28463
rect 9021 28407 9107 28463
rect 9163 28407 9249 28463
rect 9305 28407 9391 28463
rect 9447 28407 9533 28463
rect 9589 28407 9675 28463
rect 9731 28407 9817 28463
rect 9873 28407 9959 28463
rect 10015 28407 10101 28463
rect 10157 28407 10243 28463
rect 10299 28407 10385 28463
rect 10441 28407 10527 28463
rect 10583 28407 10669 28463
rect 10725 28407 10811 28463
rect 10867 28407 10953 28463
rect 11009 28407 11095 28463
rect 11151 28407 11237 28463
rect 11293 28407 11379 28463
rect 11435 28407 11521 28463
rect 11577 28407 11663 28463
rect 11719 28407 11805 28463
rect 11861 28407 11947 28463
rect 12003 28407 12089 28463
rect 12145 28407 12231 28463
rect 12287 28407 12373 28463
rect 12429 28407 12515 28463
rect 12571 28407 12657 28463
rect 12713 28407 12799 28463
rect 12855 28407 12941 28463
rect 12997 28407 13083 28463
rect 13139 28407 13225 28463
rect 13281 28407 13367 28463
rect 13423 28407 13509 28463
rect 13565 28407 13651 28463
rect 13707 28407 13793 28463
rect 13849 28407 13935 28463
rect 13991 28407 14077 28463
rect 14133 28407 14219 28463
rect 14275 28407 14361 28463
rect 14417 28407 14503 28463
rect 14559 28407 14645 28463
rect 14701 28407 14787 28463
rect 14843 28407 14853 28463
rect 151 28321 14853 28407
rect 151 28265 161 28321
rect 217 28265 303 28321
rect 359 28265 445 28321
rect 501 28265 587 28321
rect 643 28265 729 28321
rect 785 28265 871 28321
rect 927 28265 1013 28321
rect 1069 28265 1155 28321
rect 1211 28265 1297 28321
rect 1353 28265 1439 28321
rect 1495 28265 1581 28321
rect 1637 28265 1723 28321
rect 1779 28265 1865 28321
rect 1921 28265 2007 28321
rect 2063 28265 2149 28321
rect 2205 28265 2291 28321
rect 2347 28265 2433 28321
rect 2489 28265 2575 28321
rect 2631 28265 2717 28321
rect 2773 28265 2859 28321
rect 2915 28265 3001 28321
rect 3057 28265 3143 28321
rect 3199 28265 3285 28321
rect 3341 28265 3427 28321
rect 3483 28265 3569 28321
rect 3625 28265 3711 28321
rect 3767 28265 3853 28321
rect 3909 28265 3995 28321
rect 4051 28265 4137 28321
rect 4193 28265 4279 28321
rect 4335 28265 4421 28321
rect 4477 28265 4563 28321
rect 4619 28265 4705 28321
rect 4761 28265 4847 28321
rect 4903 28265 4989 28321
rect 5045 28265 5131 28321
rect 5187 28265 5273 28321
rect 5329 28265 5415 28321
rect 5471 28265 5557 28321
rect 5613 28265 5699 28321
rect 5755 28265 5841 28321
rect 5897 28265 5983 28321
rect 6039 28265 6125 28321
rect 6181 28265 6267 28321
rect 6323 28265 6409 28321
rect 6465 28265 6551 28321
rect 6607 28265 6693 28321
rect 6749 28265 6835 28321
rect 6891 28265 6977 28321
rect 7033 28265 7119 28321
rect 7175 28265 7261 28321
rect 7317 28265 7403 28321
rect 7459 28265 7545 28321
rect 7601 28265 7687 28321
rect 7743 28265 7829 28321
rect 7885 28265 7971 28321
rect 8027 28265 8113 28321
rect 8169 28265 8255 28321
rect 8311 28265 8397 28321
rect 8453 28265 8539 28321
rect 8595 28265 8681 28321
rect 8737 28265 8823 28321
rect 8879 28265 8965 28321
rect 9021 28265 9107 28321
rect 9163 28265 9249 28321
rect 9305 28265 9391 28321
rect 9447 28265 9533 28321
rect 9589 28265 9675 28321
rect 9731 28265 9817 28321
rect 9873 28265 9959 28321
rect 10015 28265 10101 28321
rect 10157 28265 10243 28321
rect 10299 28265 10385 28321
rect 10441 28265 10527 28321
rect 10583 28265 10669 28321
rect 10725 28265 10811 28321
rect 10867 28265 10953 28321
rect 11009 28265 11095 28321
rect 11151 28265 11237 28321
rect 11293 28265 11379 28321
rect 11435 28265 11521 28321
rect 11577 28265 11663 28321
rect 11719 28265 11805 28321
rect 11861 28265 11947 28321
rect 12003 28265 12089 28321
rect 12145 28265 12231 28321
rect 12287 28265 12373 28321
rect 12429 28265 12515 28321
rect 12571 28265 12657 28321
rect 12713 28265 12799 28321
rect 12855 28265 12941 28321
rect 12997 28265 13083 28321
rect 13139 28265 13225 28321
rect 13281 28265 13367 28321
rect 13423 28265 13509 28321
rect 13565 28265 13651 28321
rect 13707 28265 13793 28321
rect 13849 28265 13935 28321
rect 13991 28265 14077 28321
rect 14133 28265 14219 28321
rect 14275 28265 14361 28321
rect 14417 28265 14503 28321
rect 14559 28265 14645 28321
rect 14701 28265 14787 28321
rect 14843 28265 14853 28321
rect 151 28179 14853 28265
rect 151 28123 161 28179
rect 217 28123 303 28179
rect 359 28123 445 28179
rect 501 28123 587 28179
rect 643 28123 729 28179
rect 785 28123 871 28179
rect 927 28123 1013 28179
rect 1069 28123 1155 28179
rect 1211 28123 1297 28179
rect 1353 28123 1439 28179
rect 1495 28123 1581 28179
rect 1637 28123 1723 28179
rect 1779 28123 1865 28179
rect 1921 28123 2007 28179
rect 2063 28123 2149 28179
rect 2205 28123 2291 28179
rect 2347 28123 2433 28179
rect 2489 28123 2575 28179
rect 2631 28123 2717 28179
rect 2773 28123 2859 28179
rect 2915 28123 3001 28179
rect 3057 28123 3143 28179
rect 3199 28123 3285 28179
rect 3341 28123 3427 28179
rect 3483 28123 3569 28179
rect 3625 28123 3711 28179
rect 3767 28123 3853 28179
rect 3909 28123 3995 28179
rect 4051 28123 4137 28179
rect 4193 28123 4279 28179
rect 4335 28123 4421 28179
rect 4477 28123 4563 28179
rect 4619 28123 4705 28179
rect 4761 28123 4847 28179
rect 4903 28123 4989 28179
rect 5045 28123 5131 28179
rect 5187 28123 5273 28179
rect 5329 28123 5415 28179
rect 5471 28123 5557 28179
rect 5613 28123 5699 28179
rect 5755 28123 5841 28179
rect 5897 28123 5983 28179
rect 6039 28123 6125 28179
rect 6181 28123 6267 28179
rect 6323 28123 6409 28179
rect 6465 28123 6551 28179
rect 6607 28123 6693 28179
rect 6749 28123 6835 28179
rect 6891 28123 6977 28179
rect 7033 28123 7119 28179
rect 7175 28123 7261 28179
rect 7317 28123 7403 28179
rect 7459 28123 7545 28179
rect 7601 28123 7687 28179
rect 7743 28123 7829 28179
rect 7885 28123 7971 28179
rect 8027 28123 8113 28179
rect 8169 28123 8255 28179
rect 8311 28123 8397 28179
rect 8453 28123 8539 28179
rect 8595 28123 8681 28179
rect 8737 28123 8823 28179
rect 8879 28123 8965 28179
rect 9021 28123 9107 28179
rect 9163 28123 9249 28179
rect 9305 28123 9391 28179
rect 9447 28123 9533 28179
rect 9589 28123 9675 28179
rect 9731 28123 9817 28179
rect 9873 28123 9959 28179
rect 10015 28123 10101 28179
rect 10157 28123 10243 28179
rect 10299 28123 10385 28179
rect 10441 28123 10527 28179
rect 10583 28123 10669 28179
rect 10725 28123 10811 28179
rect 10867 28123 10953 28179
rect 11009 28123 11095 28179
rect 11151 28123 11237 28179
rect 11293 28123 11379 28179
rect 11435 28123 11521 28179
rect 11577 28123 11663 28179
rect 11719 28123 11805 28179
rect 11861 28123 11947 28179
rect 12003 28123 12089 28179
rect 12145 28123 12231 28179
rect 12287 28123 12373 28179
rect 12429 28123 12515 28179
rect 12571 28123 12657 28179
rect 12713 28123 12799 28179
rect 12855 28123 12941 28179
rect 12997 28123 13083 28179
rect 13139 28123 13225 28179
rect 13281 28123 13367 28179
rect 13423 28123 13509 28179
rect 13565 28123 13651 28179
rect 13707 28123 13793 28179
rect 13849 28123 13935 28179
rect 13991 28123 14077 28179
rect 14133 28123 14219 28179
rect 14275 28123 14361 28179
rect 14417 28123 14503 28179
rect 14559 28123 14645 28179
rect 14701 28123 14787 28179
rect 14843 28123 14853 28179
rect 151 28037 14853 28123
rect 151 27981 161 28037
rect 217 27981 303 28037
rect 359 27981 445 28037
rect 501 27981 587 28037
rect 643 27981 729 28037
rect 785 27981 871 28037
rect 927 27981 1013 28037
rect 1069 27981 1155 28037
rect 1211 27981 1297 28037
rect 1353 27981 1439 28037
rect 1495 27981 1581 28037
rect 1637 27981 1723 28037
rect 1779 27981 1865 28037
rect 1921 27981 2007 28037
rect 2063 27981 2149 28037
rect 2205 27981 2291 28037
rect 2347 27981 2433 28037
rect 2489 27981 2575 28037
rect 2631 27981 2717 28037
rect 2773 27981 2859 28037
rect 2915 27981 3001 28037
rect 3057 27981 3143 28037
rect 3199 27981 3285 28037
rect 3341 27981 3427 28037
rect 3483 27981 3569 28037
rect 3625 27981 3711 28037
rect 3767 27981 3853 28037
rect 3909 27981 3995 28037
rect 4051 27981 4137 28037
rect 4193 27981 4279 28037
rect 4335 27981 4421 28037
rect 4477 27981 4563 28037
rect 4619 27981 4705 28037
rect 4761 27981 4847 28037
rect 4903 27981 4989 28037
rect 5045 27981 5131 28037
rect 5187 27981 5273 28037
rect 5329 27981 5415 28037
rect 5471 27981 5557 28037
rect 5613 27981 5699 28037
rect 5755 27981 5841 28037
rect 5897 27981 5983 28037
rect 6039 27981 6125 28037
rect 6181 27981 6267 28037
rect 6323 27981 6409 28037
rect 6465 27981 6551 28037
rect 6607 27981 6693 28037
rect 6749 27981 6835 28037
rect 6891 27981 6977 28037
rect 7033 27981 7119 28037
rect 7175 27981 7261 28037
rect 7317 27981 7403 28037
rect 7459 27981 7545 28037
rect 7601 27981 7687 28037
rect 7743 27981 7829 28037
rect 7885 27981 7971 28037
rect 8027 27981 8113 28037
rect 8169 27981 8255 28037
rect 8311 27981 8397 28037
rect 8453 27981 8539 28037
rect 8595 27981 8681 28037
rect 8737 27981 8823 28037
rect 8879 27981 8965 28037
rect 9021 27981 9107 28037
rect 9163 27981 9249 28037
rect 9305 27981 9391 28037
rect 9447 27981 9533 28037
rect 9589 27981 9675 28037
rect 9731 27981 9817 28037
rect 9873 27981 9959 28037
rect 10015 27981 10101 28037
rect 10157 27981 10243 28037
rect 10299 27981 10385 28037
rect 10441 27981 10527 28037
rect 10583 27981 10669 28037
rect 10725 27981 10811 28037
rect 10867 27981 10953 28037
rect 11009 27981 11095 28037
rect 11151 27981 11237 28037
rect 11293 27981 11379 28037
rect 11435 27981 11521 28037
rect 11577 27981 11663 28037
rect 11719 27981 11805 28037
rect 11861 27981 11947 28037
rect 12003 27981 12089 28037
rect 12145 27981 12231 28037
rect 12287 27981 12373 28037
rect 12429 27981 12515 28037
rect 12571 27981 12657 28037
rect 12713 27981 12799 28037
rect 12855 27981 12941 28037
rect 12997 27981 13083 28037
rect 13139 27981 13225 28037
rect 13281 27981 13367 28037
rect 13423 27981 13509 28037
rect 13565 27981 13651 28037
rect 13707 27981 13793 28037
rect 13849 27981 13935 28037
rect 13991 27981 14077 28037
rect 14133 27981 14219 28037
rect 14275 27981 14361 28037
rect 14417 27981 14503 28037
rect 14559 27981 14645 28037
rect 14701 27981 14787 28037
rect 14843 27981 14853 28037
rect 151 27895 14853 27981
rect 151 27839 161 27895
rect 217 27839 303 27895
rect 359 27839 445 27895
rect 501 27839 587 27895
rect 643 27839 729 27895
rect 785 27839 871 27895
rect 927 27839 1013 27895
rect 1069 27839 1155 27895
rect 1211 27839 1297 27895
rect 1353 27839 1439 27895
rect 1495 27839 1581 27895
rect 1637 27839 1723 27895
rect 1779 27839 1865 27895
rect 1921 27839 2007 27895
rect 2063 27839 2149 27895
rect 2205 27839 2291 27895
rect 2347 27839 2433 27895
rect 2489 27839 2575 27895
rect 2631 27839 2717 27895
rect 2773 27839 2859 27895
rect 2915 27839 3001 27895
rect 3057 27839 3143 27895
rect 3199 27839 3285 27895
rect 3341 27839 3427 27895
rect 3483 27839 3569 27895
rect 3625 27839 3711 27895
rect 3767 27839 3853 27895
rect 3909 27839 3995 27895
rect 4051 27839 4137 27895
rect 4193 27839 4279 27895
rect 4335 27839 4421 27895
rect 4477 27839 4563 27895
rect 4619 27839 4705 27895
rect 4761 27839 4847 27895
rect 4903 27839 4989 27895
rect 5045 27839 5131 27895
rect 5187 27839 5273 27895
rect 5329 27839 5415 27895
rect 5471 27839 5557 27895
rect 5613 27839 5699 27895
rect 5755 27839 5841 27895
rect 5897 27839 5983 27895
rect 6039 27839 6125 27895
rect 6181 27839 6267 27895
rect 6323 27839 6409 27895
rect 6465 27839 6551 27895
rect 6607 27839 6693 27895
rect 6749 27839 6835 27895
rect 6891 27839 6977 27895
rect 7033 27839 7119 27895
rect 7175 27839 7261 27895
rect 7317 27839 7403 27895
rect 7459 27839 7545 27895
rect 7601 27839 7687 27895
rect 7743 27839 7829 27895
rect 7885 27839 7971 27895
rect 8027 27839 8113 27895
rect 8169 27839 8255 27895
rect 8311 27839 8397 27895
rect 8453 27839 8539 27895
rect 8595 27839 8681 27895
rect 8737 27839 8823 27895
rect 8879 27839 8965 27895
rect 9021 27839 9107 27895
rect 9163 27839 9249 27895
rect 9305 27839 9391 27895
rect 9447 27839 9533 27895
rect 9589 27839 9675 27895
rect 9731 27839 9817 27895
rect 9873 27839 9959 27895
rect 10015 27839 10101 27895
rect 10157 27839 10243 27895
rect 10299 27839 10385 27895
rect 10441 27839 10527 27895
rect 10583 27839 10669 27895
rect 10725 27839 10811 27895
rect 10867 27839 10953 27895
rect 11009 27839 11095 27895
rect 11151 27839 11237 27895
rect 11293 27839 11379 27895
rect 11435 27839 11521 27895
rect 11577 27839 11663 27895
rect 11719 27839 11805 27895
rect 11861 27839 11947 27895
rect 12003 27839 12089 27895
rect 12145 27839 12231 27895
rect 12287 27839 12373 27895
rect 12429 27839 12515 27895
rect 12571 27839 12657 27895
rect 12713 27839 12799 27895
rect 12855 27839 12941 27895
rect 12997 27839 13083 27895
rect 13139 27839 13225 27895
rect 13281 27839 13367 27895
rect 13423 27839 13509 27895
rect 13565 27839 13651 27895
rect 13707 27839 13793 27895
rect 13849 27839 13935 27895
rect 13991 27839 14077 27895
rect 14133 27839 14219 27895
rect 14275 27839 14361 27895
rect 14417 27839 14503 27895
rect 14559 27839 14645 27895
rect 14701 27839 14787 27895
rect 14843 27839 14853 27895
rect 151 27753 14853 27839
rect 151 27697 161 27753
rect 217 27697 303 27753
rect 359 27697 445 27753
rect 501 27697 587 27753
rect 643 27697 729 27753
rect 785 27697 871 27753
rect 927 27697 1013 27753
rect 1069 27697 1155 27753
rect 1211 27697 1297 27753
rect 1353 27697 1439 27753
rect 1495 27697 1581 27753
rect 1637 27697 1723 27753
rect 1779 27697 1865 27753
rect 1921 27697 2007 27753
rect 2063 27697 2149 27753
rect 2205 27697 2291 27753
rect 2347 27697 2433 27753
rect 2489 27697 2575 27753
rect 2631 27697 2717 27753
rect 2773 27697 2859 27753
rect 2915 27697 3001 27753
rect 3057 27697 3143 27753
rect 3199 27697 3285 27753
rect 3341 27697 3427 27753
rect 3483 27697 3569 27753
rect 3625 27697 3711 27753
rect 3767 27697 3853 27753
rect 3909 27697 3995 27753
rect 4051 27697 4137 27753
rect 4193 27697 4279 27753
rect 4335 27697 4421 27753
rect 4477 27697 4563 27753
rect 4619 27697 4705 27753
rect 4761 27697 4847 27753
rect 4903 27697 4989 27753
rect 5045 27697 5131 27753
rect 5187 27697 5273 27753
rect 5329 27697 5415 27753
rect 5471 27697 5557 27753
rect 5613 27697 5699 27753
rect 5755 27697 5841 27753
rect 5897 27697 5983 27753
rect 6039 27697 6125 27753
rect 6181 27697 6267 27753
rect 6323 27697 6409 27753
rect 6465 27697 6551 27753
rect 6607 27697 6693 27753
rect 6749 27697 6835 27753
rect 6891 27697 6977 27753
rect 7033 27697 7119 27753
rect 7175 27697 7261 27753
rect 7317 27697 7403 27753
rect 7459 27697 7545 27753
rect 7601 27697 7687 27753
rect 7743 27697 7829 27753
rect 7885 27697 7971 27753
rect 8027 27697 8113 27753
rect 8169 27697 8255 27753
rect 8311 27697 8397 27753
rect 8453 27697 8539 27753
rect 8595 27697 8681 27753
rect 8737 27697 8823 27753
rect 8879 27697 8965 27753
rect 9021 27697 9107 27753
rect 9163 27697 9249 27753
rect 9305 27697 9391 27753
rect 9447 27697 9533 27753
rect 9589 27697 9675 27753
rect 9731 27697 9817 27753
rect 9873 27697 9959 27753
rect 10015 27697 10101 27753
rect 10157 27697 10243 27753
rect 10299 27697 10385 27753
rect 10441 27697 10527 27753
rect 10583 27697 10669 27753
rect 10725 27697 10811 27753
rect 10867 27697 10953 27753
rect 11009 27697 11095 27753
rect 11151 27697 11237 27753
rect 11293 27697 11379 27753
rect 11435 27697 11521 27753
rect 11577 27697 11663 27753
rect 11719 27697 11805 27753
rect 11861 27697 11947 27753
rect 12003 27697 12089 27753
rect 12145 27697 12231 27753
rect 12287 27697 12373 27753
rect 12429 27697 12515 27753
rect 12571 27697 12657 27753
rect 12713 27697 12799 27753
rect 12855 27697 12941 27753
rect 12997 27697 13083 27753
rect 13139 27697 13225 27753
rect 13281 27697 13367 27753
rect 13423 27697 13509 27753
rect 13565 27697 13651 27753
rect 13707 27697 13793 27753
rect 13849 27697 13935 27753
rect 13991 27697 14077 27753
rect 14133 27697 14219 27753
rect 14275 27697 14361 27753
rect 14417 27697 14503 27753
rect 14559 27697 14645 27753
rect 14701 27697 14787 27753
rect 14843 27697 14853 27753
rect 151 27611 14853 27697
rect 151 27555 161 27611
rect 217 27555 303 27611
rect 359 27555 445 27611
rect 501 27555 587 27611
rect 643 27555 729 27611
rect 785 27555 871 27611
rect 927 27555 1013 27611
rect 1069 27555 1155 27611
rect 1211 27555 1297 27611
rect 1353 27555 1439 27611
rect 1495 27555 1581 27611
rect 1637 27555 1723 27611
rect 1779 27555 1865 27611
rect 1921 27555 2007 27611
rect 2063 27555 2149 27611
rect 2205 27555 2291 27611
rect 2347 27555 2433 27611
rect 2489 27555 2575 27611
rect 2631 27555 2717 27611
rect 2773 27555 2859 27611
rect 2915 27555 3001 27611
rect 3057 27555 3143 27611
rect 3199 27555 3285 27611
rect 3341 27555 3427 27611
rect 3483 27555 3569 27611
rect 3625 27555 3711 27611
rect 3767 27555 3853 27611
rect 3909 27555 3995 27611
rect 4051 27555 4137 27611
rect 4193 27555 4279 27611
rect 4335 27555 4421 27611
rect 4477 27555 4563 27611
rect 4619 27555 4705 27611
rect 4761 27555 4847 27611
rect 4903 27555 4989 27611
rect 5045 27555 5131 27611
rect 5187 27555 5273 27611
rect 5329 27555 5415 27611
rect 5471 27555 5557 27611
rect 5613 27555 5699 27611
rect 5755 27555 5841 27611
rect 5897 27555 5983 27611
rect 6039 27555 6125 27611
rect 6181 27555 6267 27611
rect 6323 27555 6409 27611
rect 6465 27555 6551 27611
rect 6607 27555 6693 27611
rect 6749 27555 6835 27611
rect 6891 27555 6977 27611
rect 7033 27555 7119 27611
rect 7175 27555 7261 27611
rect 7317 27555 7403 27611
rect 7459 27555 7545 27611
rect 7601 27555 7687 27611
rect 7743 27555 7829 27611
rect 7885 27555 7971 27611
rect 8027 27555 8113 27611
rect 8169 27555 8255 27611
rect 8311 27555 8397 27611
rect 8453 27555 8539 27611
rect 8595 27555 8681 27611
rect 8737 27555 8823 27611
rect 8879 27555 8965 27611
rect 9021 27555 9107 27611
rect 9163 27555 9249 27611
rect 9305 27555 9391 27611
rect 9447 27555 9533 27611
rect 9589 27555 9675 27611
rect 9731 27555 9817 27611
rect 9873 27555 9959 27611
rect 10015 27555 10101 27611
rect 10157 27555 10243 27611
rect 10299 27555 10385 27611
rect 10441 27555 10527 27611
rect 10583 27555 10669 27611
rect 10725 27555 10811 27611
rect 10867 27555 10953 27611
rect 11009 27555 11095 27611
rect 11151 27555 11237 27611
rect 11293 27555 11379 27611
rect 11435 27555 11521 27611
rect 11577 27555 11663 27611
rect 11719 27555 11805 27611
rect 11861 27555 11947 27611
rect 12003 27555 12089 27611
rect 12145 27555 12231 27611
rect 12287 27555 12373 27611
rect 12429 27555 12515 27611
rect 12571 27555 12657 27611
rect 12713 27555 12799 27611
rect 12855 27555 12941 27611
rect 12997 27555 13083 27611
rect 13139 27555 13225 27611
rect 13281 27555 13367 27611
rect 13423 27555 13509 27611
rect 13565 27555 13651 27611
rect 13707 27555 13793 27611
rect 13849 27555 13935 27611
rect 13991 27555 14077 27611
rect 14133 27555 14219 27611
rect 14275 27555 14361 27611
rect 14417 27555 14503 27611
rect 14559 27555 14645 27611
rect 14701 27555 14787 27611
rect 14843 27555 14853 27611
rect 151 27469 14853 27555
rect 151 27413 161 27469
rect 217 27413 303 27469
rect 359 27413 445 27469
rect 501 27413 587 27469
rect 643 27413 729 27469
rect 785 27413 871 27469
rect 927 27413 1013 27469
rect 1069 27413 1155 27469
rect 1211 27413 1297 27469
rect 1353 27413 1439 27469
rect 1495 27413 1581 27469
rect 1637 27413 1723 27469
rect 1779 27413 1865 27469
rect 1921 27413 2007 27469
rect 2063 27413 2149 27469
rect 2205 27413 2291 27469
rect 2347 27413 2433 27469
rect 2489 27413 2575 27469
rect 2631 27413 2717 27469
rect 2773 27413 2859 27469
rect 2915 27413 3001 27469
rect 3057 27413 3143 27469
rect 3199 27413 3285 27469
rect 3341 27413 3427 27469
rect 3483 27413 3569 27469
rect 3625 27413 3711 27469
rect 3767 27413 3853 27469
rect 3909 27413 3995 27469
rect 4051 27413 4137 27469
rect 4193 27413 4279 27469
rect 4335 27413 4421 27469
rect 4477 27413 4563 27469
rect 4619 27413 4705 27469
rect 4761 27413 4847 27469
rect 4903 27413 4989 27469
rect 5045 27413 5131 27469
rect 5187 27413 5273 27469
rect 5329 27413 5415 27469
rect 5471 27413 5557 27469
rect 5613 27413 5699 27469
rect 5755 27413 5841 27469
rect 5897 27413 5983 27469
rect 6039 27413 6125 27469
rect 6181 27413 6267 27469
rect 6323 27413 6409 27469
rect 6465 27413 6551 27469
rect 6607 27413 6693 27469
rect 6749 27413 6835 27469
rect 6891 27413 6977 27469
rect 7033 27413 7119 27469
rect 7175 27413 7261 27469
rect 7317 27413 7403 27469
rect 7459 27413 7545 27469
rect 7601 27413 7687 27469
rect 7743 27413 7829 27469
rect 7885 27413 7971 27469
rect 8027 27413 8113 27469
rect 8169 27413 8255 27469
rect 8311 27413 8397 27469
rect 8453 27413 8539 27469
rect 8595 27413 8681 27469
rect 8737 27413 8823 27469
rect 8879 27413 8965 27469
rect 9021 27413 9107 27469
rect 9163 27413 9249 27469
rect 9305 27413 9391 27469
rect 9447 27413 9533 27469
rect 9589 27413 9675 27469
rect 9731 27413 9817 27469
rect 9873 27413 9959 27469
rect 10015 27413 10101 27469
rect 10157 27413 10243 27469
rect 10299 27413 10385 27469
rect 10441 27413 10527 27469
rect 10583 27413 10669 27469
rect 10725 27413 10811 27469
rect 10867 27413 10953 27469
rect 11009 27413 11095 27469
rect 11151 27413 11237 27469
rect 11293 27413 11379 27469
rect 11435 27413 11521 27469
rect 11577 27413 11663 27469
rect 11719 27413 11805 27469
rect 11861 27413 11947 27469
rect 12003 27413 12089 27469
rect 12145 27413 12231 27469
rect 12287 27413 12373 27469
rect 12429 27413 12515 27469
rect 12571 27413 12657 27469
rect 12713 27413 12799 27469
rect 12855 27413 12941 27469
rect 12997 27413 13083 27469
rect 13139 27413 13225 27469
rect 13281 27413 13367 27469
rect 13423 27413 13509 27469
rect 13565 27413 13651 27469
rect 13707 27413 13793 27469
rect 13849 27413 13935 27469
rect 13991 27413 14077 27469
rect 14133 27413 14219 27469
rect 14275 27413 14361 27469
rect 14417 27413 14503 27469
rect 14559 27413 14645 27469
rect 14701 27413 14787 27469
rect 14843 27413 14853 27469
rect 151 27327 14853 27413
rect 151 27271 161 27327
rect 217 27271 303 27327
rect 359 27271 445 27327
rect 501 27271 587 27327
rect 643 27271 729 27327
rect 785 27271 871 27327
rect 927 27271 1013 27327
rect 1069 27271 1155 27327
rect 1211 27271 1297 27327
rect 1353 27271 1439 27327
rect 1495 27271 1581 27327
rect 1637 27271 1723 27327
rect 1779 27271 1865 27327
rect 1921 27271 2007 27327
rect 2063 27271 2149 27327
rect 2205 27271 2291 27327
rect 2347 27271 2433 27327
rect 2489 27271 2575 27327
rect 2631 27271 2717 27327
rect 2773 27271 2859 27327
rect 2915 27271 3001 27327
rect 3057 27271 3143 27327
rect 3199 27271 3285 27327
rect 3341 27271 3427 27327
rect 3483 27271 3569 27327
rect 3625 27271 3711 27327
rect 3767 27271 3853 27327
rect 3909 27271 3995 27327
rect 4051 27271 4137 27327
rect 4193 27271 4279 27327
rect 4335 27271 4421 27327
rect 4477 27271 4563 27327
rect 4619 27271 4705 27327
rect 4761 27271 4847 27327
rect 4903 27271 4989 27327
rect 5045 27271 5131 27327
rect 5187 27271 5273 27327
rect 5329 27271 5415 27327
rect 5471 27271 5557 27327
rect 5613 27271 5699 27327
rect 5755 27271 5841 27327
rect 5897 27271 5983 27327
rect 6039 27271 6125 27327
rect 6181 27271 6267 27327
rect 6323 27271 6409 27327
rect 6465 27271 6551 27327
rect 6607 27271 6693 27327
rect 6749 27271 6835 27327
rect 6891 27271 6977 27327
rect 7033 27271 7119 27327
rect 7175 27271 7261 27327
rect 7317 27271 7403 27327
rect 7459 27271 7545 27327
rect 7601 27271 7687 27327
rect 7743 27271 7829 27327
rect 7885 27271 7971 27327
rect 8027 27271 8113 27327
rect 8169 27271 8255 27327
rect 8311 27271 8397 27327
rect 8453 27271 8539 27327
rect 8595 27271 8681 27327
rect 8737 27271 8823 27327
rect 8879 27271 8965 27327
rect 9021 27271 9107 27327
rect 9163 27271 9249 27327
rect 9305 27271 9391 27327
rect 9447 27271 9533 27327
rect 9589 27271 9675 27327
rect 9731 27271 9817 27327
rect 9873 27271 9959 27327
rect 10015 27271 10101 27327
rect 10157 27271 10243 27327
rect 10299 27271 10385 27327
rect 10441 27271 10527 27327
rect 10583 27271 10669 27327
rect 10725 27271 10811 27327
rect 10867 27271 10953 27327
rect 11009 27271 11095 27327
rect 11151 27271 11237 27327
rect 11293 27271 11379 27327
rect 11435 27271 11521 27327
rect 11577 27271 11663 27327
rect 11719 27271 11805 27327
rect 11861 27271 11947 27327
rect 12003 27271 12089 27327
rect 12145 27271 12231 27327
rect 12287 27271 12373 27327
rect 12429 27271 12515 27327
rect 12571 27271 12657 27327
rect 12713 27271 12799 27327
rect 12855 27271 12941 27327
rect 12997 27271 13083 27327
rect 13139 27271 13225 27327
rect 13281 27271 13367 27327
rect 13423 27271 13509 27327
rect 13565 27271 13651 27327
rect 13707 27271 13793 27327
rect 13849 27271 13935 27327
rect 13991 27271 14077 27327
rect 14133 27271 14219 27327
rect 14275 27271 14361 27327
rect 14417 27271 14503 27327
rect 14559 27271 14645 27327
rect 14701 27271 14787 27327
rect 14843 27271 14853 27327
rect 151 27185 14853 27271
rect 151 27129 161 27185
rect 217 27129 303 27185
rect 359 27129 445 27185
rect 501 27129 587 27185
rect 643 27129 729 27185
rect 785 27129 871 27185
rect 927 27129 1013 27185
rect 1069 27129 1155 27185
rect 1211 27129 1297 27185
rect 1353 27129 1439 27185
rect 1495 27129 1581 27185
rect 1637 27129 1723 27185
rect 1779 27129 1865 27185
rect 1921 27129 2007 27185
rect 2063 27129 2149 27185
rect 2205 27129 2291 27185
rect 2347 27129 2433 27185
rect 2489 27129 2575 27185
rect 2631 27129 2717 27185
rect 2773 27129 2859 27185
rect 2915 27129 3001 27185
rect 3057 27129 3143 27185
rect 3199 27129 3285 27185
rect 3341 27129 3427 27185
rect 3483 27129 3569 27185
rect 3625 27129 3711 27185
rect 3767 27129 3853 27185
rect 3909 27129 3995 27185
rect 4051 27129 4137 27185
rect 4193 27129 4279 27185
rect 4335 27129 4421 27185
rect 4477 27129 4563 27185
rect 4619 27129 4705 27185
rect 4761 27129 4847 27185
rect 4903 27129 4989 27185
rect 5045 27129 5131 27185
rect 5187 27129 5273 27185
rect 5329 27129 5415 27185
rect 5471 27129 5557 27185
rect 5613 27129 5699 27185
rect 5755 27129 5841 27185
rect 5897 27129 5983 27185
rect 6039 27129 6125 27185
rect 6181 27129 6267 27185
rect 6323 27129 6409 27185
rect 6465 27129 6551 27185
rect 6607 27129 6693 27185
rect 6749 27129 6835 27185
rect 6891 27129 6977 27185
rect 7033 27129 7119 27185
rect 7175 27129 7261 27185
rect 7317 27129 7403 27185
rect 7459 27129 7545 27185
rect 7601 27129 7687 27185
rect 7743 27129 7829 27185
rect 7885 27129 7971 27185
rect 8027 27129 8113 27185
rect 8169 27129 8255 27185
rect 8311 27129 8397 27185
rect 8453 27129 8539 27185
rect 8595 27129 8681 27185
rect 8737 27129 8823 27185
rect 8879 27129 8965 27185
rect 9021 27129 9107 27185
rect 9163 27129 9249 27185
rect 9305 27129 9391 27185
rect 9447 27129 9533 27185
rect 9589 27129 9675 27185
rect 9731 27129 9817 27185
rect 9873 27129 9959 27185
rect 10015 27129 10101 27185
rect 10157 27129 10243 27185
rect 10299 27129 10385 27185
rect 10441 27129 10527 27185
rect 10583 27129 10669 27185
rect 10725 27129 10811 27185
rect 10867 27129 10953 27185
rect 11009 27129 11095 27185
rect 11151 27129 11237 27185
rect 11293 27129 11379 27185
rect 11435 27129 11521 27185
rect 11577 27129 11663 27185
rect 11719 27129 11805 27185
rect 11861 27129 11947 27185
rect 12003 27129 12089 27185
rect 12145 27129 12231 27185
rect 12287 27129 12373 27185
rect 12429 27129 12515 27185
rect 12571 27129 12657 27185
rect 12713 27129 12799 27185
rect 12855 27129 12941 27185
rect 12997 27129 13083 27185
rect 13139 27129 13225 27185
rect 13281 27129 13367 27185
rect 13423 27129 13509 27185
rect 13565 27129 13651 27185
rect 13707 27129 13793 27185
rect 13849 27129 13935 27185
rect 13991 27129 14077 27185
rect 14133 27129 14219 27185
rect 14275 27129 14361 27185
rect 14417 27129 14503 27185
rect 14559 27129 14645 27185
rect 14701 27129 14787 27185
rect 14843 27129 14853 27185
rect 151 27043 14853 27129
rect 151 26987 161 27043
rect 217 26987 303 27043
rect 359 26987 445 27043
rect 501 26987 587 27043
rect 643 26987 729 27043
rect 785 26987 871 27043
rect 927 26987 1013 27043
rect 1069 26987 1155 27043
rect 1211 26987 1297 27043
rect 1353 26987 1439 27043
rect 1495 26987 1581 27043
rect 1637 26987 1723 27043
rect 1779 26987 1865 27043
rect 1921 26987 2007 27043
rect 2063 26987 2149 27043
rect 2205 26987 2291 27043
rect 2347 26987 2433 27043
rect 2489 26987 2575 27043
rect 2631 26987 2717 27043
rect 2773 26987 2859 27043
rect 2915 26987 3001 27043
rect 3057 26987 3143 27043
rect 3199 26987 3285 27043
rect 3341 26987 3427 27043
rect 3483 26987 3569 27043
rect 3625 26987 3711 27043
rect 3767 26987 3853 27043
rect 3909 26987 3995 27043
rect 4051 26987 4137 27043
rect 4193 26987 4279 27043
rect 4335 26987 4421 27043
rect 4477 26987 4563 27043
rect 4619 26987 4705 27043
rect 4761 26987 4847 27043
rect 4903 26987 4989 27043
rect 5045 26987 5131 27043
rect 5187 26987 5273 27043
rect 5329 26987 5415 27043
rect 5471 26987 5557 27043
rect 5613 26987 5699 27043
rect 5755 26987 5841 27043
rect 5897 26987 5983 27043
rect 6039 26987 6125 27043
rect 6181 26987 6267 27043
rect 6323 26987 6409 27043
rect 6465 26987 6551 27043
rect 6607 26987 6693 27043
rect 6749 26987 6835 27043
rect 6891 26987 6977 27043
rect 7033 26987 7119 27043
rect 7175 26987 7261 27043
rect 7317 26987 7403 27043
rect 7459 26987 7545 27043
rect 7601 26987 7687 27043
rect 7743 26987 7829 27043
rect 7885 26987 7971 27043
rect 8027 26987 8113 27043
rect 8169 26987 8255 27043
rect 8311 26987 8397 27043
rect 8453 26987 8539 27043
rect 8595 26987 8681 27043
rect 8737 26987 8823 27043
rect 8879 26987 8965 27043
rect 9021 26987 9107 27043
rect 9163 26987 9249 27043
rect 9305 26987 9391 27043
rect 9447 26987 9533 27043
rect 9589 26987 9675 27043
rect 9731 26987 9817 27043
rect 9873 26987 9959 27043
rect 10015 26987 10101 27043
rect 10157 26987 10243 27043
rect 10299 26987 10385 27043
rect 10441 26987 10527 27043
rect 10583 26987 10669 27043
rect 10725 26987 10811 27043
rect 10867 26987 10953 27043
rect 11009 26987 11095 27043
rect 11151 26987 11237 27043
rect 11293 26987 11379 27043
rect 11435 26987 11521 27043
rect 11577 26987 11663 27043
rect 11719 26987 11805 27043
rect 11861 26987 11947 27043
rect 12003 26987 12089 27043
rect 12145 26987 12231 27043
rect 12287 26987 12373 27043
rect 12429 26987 12515 27043
rect 12571 26987 12657 27043
rect 12713 26987 12799 27043
rect 12855 26987 12941 27043
rect 12997 26987 13083 27043
rect 13139 26987 13225 27043
rect 13281 26987 13367 27043
rect 13423 26987 13509 27043
rect 13565 26987 13651 27043
rect 13707 26987 13793 27043
rect 13849 26987 13935 27043
rect 13991 26987 14077 27043
rect 14133 26987 14219 27043
rect 14275 26987 14361 27043
rect 14417 26987 14503 27043
rect 14559 26987 14645 27043
rect 14701 26987 14787 27043
rect 14843 26987 14853 27043
rect 151 26901 14853 26987
rect 151 26845 161 26901
rect 217 26845 303 26901
rect 359 26845 445 26901
rect 501 26845 587 26901
rect 643 26845 729 26901
rect 785 26845 871 26901
rect 927 26845 1013 26901
rect 1069 26845 1155 26901
rect 1211 26845 1297 26901
rect 1353 26845 1439 26901
rect 1495 26845 1581 26901
rect 1637 26845 1723 26901
rect 1779 26845 1865 26901
rect 1921 26845 2007 26901
rect 2063 26845 2149 26901
rect 2205 26845 2291 26901
rect 2347 26845 2433 26901
rect 2489 26845 2575 26901
rect 2631 26845 2717 26901
rect 2773 26845 2859 26901
rect 2915 26845 3001 26901
rect 3057 26845 3143 26901
rect 3199 26845 3285 26901
rect 3341 26845 3427 26901
rect 3483 26845 3569 26901
rect 3625 26845 3711 26901
rect 3767 26845 3853 26901
rect 3909 26845 3995 26901
rect 4051 26845 4137 26901
rect 4193 26845 4279 26901
rect 4335 26845 4421 26901
rect 4477 26845 4563 26901
rect 4619 26845 4705 26901
rect 4761 26845 4847 26901
rect 4903 26845 4989 26901
rect 5045 26845 5131 26901
rect 5187 26845 5273 26901
rect 5329 26845 5415 26901
rect 5471 26845 5557 26901
rect 5613 26845 5699 26901
rect 5755 26845 5841 26901
rect 5897 26845 5983 26901
rect 6039 26845 6125 26901
rect 6181 26845 6267 26901
rect 6323 26845 6409 26901
rect 6465 26845 6551 26901
rect 6607 26845 6693 26901
rect 6749 26845 6835 26901
rect 6891 26845 6977 26901
rect 7033 26845 7119 26901
rect 7175 26845 7261 26901
rect 7317 26845 7403 26901
rect 7459 26845 7545 26901
rect 7601 26845 7687 26901
rect 7743 26845 7829 26901
rect 7885 26845 7971 26901
rect 8027 26845 8113 26901
rect 8169 26845 8255 26901
rect 8311 26845 8397 26901
rect 8453 26845 8539 26901
rect 8595 26845 8681 26901
rect 8737 26845 8823 26901
rect 8879 26845 8965 26901
rect 9021 26845 9107 26901
rect 9163 26845 9249 26901
rect 9305 26845 9391 26901
rect 9447 26845 9533 26901
rect 9589 26845 9675 26901
rect 9731 26845 9817 26901
rect 9873 26845 9959 26901
rect 10015 26845 10101 26901
rect 10157 26845 10243 26901
rect 10299 26845 10385 26901
rect 10441 26845 10527 26901
rect 10583 26845 10669 26901
rect 10725 26845 10811 26901
rect 10867 26845 10953 26901
rect 11009 26845 11095 26901
rect 11151 26845 11237 26901
rect 11293 26845 11379 26901
rect 11435 26845 11521 26901
rect 11577 26845 11663 26901
rect 11719 26845 11805 26901
rect 11861 26845 11947 26901
rect 12003 26845 12089 26901
rect 12145 26845 12231 26901
rect 12287 26845 12373 26901
rect 12429 26845 12515 26901
rect 12571 26845 12657 26901
rect 12713 26845 12799 26901
rect 12855 26845 12941 26901
rect 12997 26845 13083 26901
rect 13139 26845 13225 26901
rect 13281 26845 13367 26901
rect 13423 26845 13509 26901
rect 13565 26845 13651 26901
rect 13707 26845 13793 26901
rect 13849 26845 13935 26901
rect 13991 26845 14077 26901
rect 14133 26845 14219 26901
rect 14275 26845 14361 26901
rect 14417 26845 14503 26901
rect 14559 26845 14645 26901
rect 14701 26845 14787 26901
rect 14843 26845 14853 26901
rect 151 26835 14853 26845
rect 151 26563 14853 26573
rect 151 26507 161 26563
rect 217 26507 303 26563
rect 359 26507 445 26563
rect 501 26507 587 26563
rect 643 26507 729 26563
rect 785 26507 871 26563
rect 927 26507 1013 26563
rect 1069 26507 1155 26563
rect 1211 26507 1297 26563
rect 1353 26507 1439 26563
rect 1495 26507 1581 26563
rect 1637 26507 1723 26563
rect 1779 26507 1865 26563
rect 1921 26507 2007 26563
rect 2063 26507 2149 26563
rect 2205 26507 2291 26563
rect 2347 26507 2433 26563
rect 2489 26507 2575 26563
rect 2631 26507 2717 26563
rect 2773 26507 2859 26563
rect 2915 26507 3001 26563
rect 3057 26507 3143 26563
rect 3199 26507 3285 26563
rect 3341 26507 3427 26563
rect 3483 26507 3569 26563
rect 3625 26507 3711 26563
rect 3767 26507 3853 26563
rect 3909 26507 3995 26563
rect 4051 26507 4137 26563
rect 4193 26507 4279 26563
rect 4335 26507 4421 26563
rect 4477 26507 4563 26563
rect 4619 26507 4705 26563
rect 4761 26507 4847 26563
rect 4903 26507 4989 26563
rect 5045 26507 5131 26563
rect 5187 26507 5273 26563
rect 5329 26507 5415 26563
rect 5471 26507 5557 26563
rect 5613 26507 5699 26563
rect 5755 26507 5841 26563
rect 5897 26507 5983 26563
rect 6039 26507 6125 26563
rect 6181 26507 6267 26563
rect 6323 26507 6409 26563
rect 6465 26507 6551 26563
rect 6607 26507 6693 26563
rect 6749 26507 6835 26563
rect 6891 26507 6977 26563
rect 7033 26507 7119 26563
rect 7175 26507 7261 26563
rect 7317 26507 7403 26563
rect 7459 26507 7545 26563
rect 7601 26507 7687 26563
rect 7743 26507 7829 26563
rect 7885 26507 7971 26563
rect 8027 26507 8113 26563
rect 8169 26507 8255 26563
rect 8311 26507 8397 26563
rect 8453 26507 8539 26563
rect 8595 26507 8681 26563
rect 8737 26507 8823 26563
rect 8879 26507 8965 26563
rect 9021 26507 9107 26563
rect 9163 26507 9249 26563
rect 9305 26507 9391 26563
rect 9447 26507 9533 26563
rect 9589 26507 9675 26563
rect 9731 26507 9817 26563
rect 9873 26507 9959 26563
rect 10015 26507 10101 26563
rect 10157 26507 10243 26563
rect 10299 26507 10385 26563
rect 10441 26507 10527 26563
rect 10583 26507 10669 26563
rect 10725 26507 10811 26563
rect 10867 26507 10953 26563
rect 11009 26507 11095 26563
rect 11151 26507 11237 26563
rect 11293 26507 11379 26563
rect 11435 26507 11521 26563
rect 11577 26507 11663 26563
rect 11719 26507 11805 26563
rect 11861 26507 11947 26563
rect 12003 26507 12089 26563
rect 12145 26507 12231 26563
rect 12287 26507 12373 26563
rect 12429 26507 12515 26563
rect 12571 26507 12657 26563
rect 12713 26507 12799 26563
rect 12855 26507 12941 26563
rect 12997 26507 13083 26563
rect 13139 26507 13225 26563
rect 13281 26507 13367 26563
rect 13423 26507 13509 26563
rect 13565 26507 13651 26563
rect 13707 26507 13793 26563
rect 13849 26507 13935 26563
rect 13991 26507 14077 26563
rect 14133 26507 14219 26563
rect 14275 26507 14361 26563
rect 14417 26507 14503 26563
rect 14559 26507 14645 26563
rect 14701 26507 14787 26563
rect 14843 26507 14853 26563
rect 151 26421 14853 26507
rect 151 26365 161 26421
rect 217 26365 303 26421
rect 359 26365 445 26421
rect 501 26365 587 26421
rect 643 26365 729 26421
rect 785 26365 871 26421
rect 927 26365 1013 26421
rect 1069 26365 1155 26421
rect 1211 26365 1297 26421
rect 1353 26365 1439 26421
rect 1495 26365 1581 26421
rect 1637 26365 1723 26421
rect 1779 26365 1865 26421
rect 1921 26365 2007 26421
rect 2063 26365 2149 26421
rect 2205 26365 2291 26421
rect 2347 26365 2433 26421
rect 2489 26365 2575 26421
rect 2631 26365 2717 26421
rect 2773 26365 2859 26421
rect 2915 26365 3001 26421
rect 3057 26365 3143 26421
rect 3199 26365 3285 26421
rect 3341 26365 3427 26421
rect 3483 26365 3569 26421
rect 3625 26365 3711 26421
rect 3767 26365 3853 26421
rect 3909 26365 3995 26421
rect 4051 26365 4137 26421
rect 4193 26365 4279 26421
rect 4335 26365 4421 26421
rect 4477 26365 4563 26421
rect 4619 26365 4705 26421
rect 4761 26365 4847 26421
rect 4903 26365 4989 26421
rect 5045 26365 5131 26421
rect 5187 26365 5273 26421
rect 5329 26365 5415 26421
rect 5471 26365 5557 26421
rect 5613 26365 5699 26421
rect 5755 26365 5841 26421
rect 5897 26365 5983 26421
rect 6039 26365 6125 26421
rect 6181 26365 6267 26421
rect 6323 26365 6409 26421
rect 6465 26365 6551 26421
rect 6607 26365 6693 26421
rect 6749 26365 6835 26421
rect 6891 26365 6977 26421
rect 7033 26365 7119 26421
rect 7175 26365 7261 26421
rect 7317 26365 7403 26421
rect 7459 26365 7545 26421
rect 7601 26365 7687 26421
rect 7743 26365 7829 26421
rect 7885 26365 7971 26421
rect 8027 26365 8113 26421
rect 8169 26365 8255 26421
rect 8311 26365 8397 26421
rect 8453 26365 8539 26421
rect 8595 26365 8681 26421
rect 8737 26365 8823 26421
rect 8879 26365 8965 26421
rect 9021 26365 9107 26421
rect 9163 26365 9249 26421
rect 9305 26365 9391 26421
rect 9447 26365 9533 26421
rect 9589 26365 9675 26421
rect 9731 26365 9817 26421
rect 9873 26365 9959 26421
rect 10015 26365 10101 26421
rect 10157 26365 10243 26421
rect 10299 26365 10385 26421
rect 10441 26365 10527 26421
rect 10583 26365 10669 26421
rect 10725 26365 10811 26421
rect 10867 26365 10953 26421
rect 11009 26365 11095 26421
rect 11151 26365 11237 26421
rect 11293 26365 11379 26421
rect 11435 26365 11521 26421
rect 11577 26365 11663 26421
rect 11719 26365 11805 26421
rect 11861 26365 11947 26421
rect 12003 26365 12089 26421
rect 12145 26365 12231 26421
rect 12287 26365 12373 26421
rect 12429 26365 12515 26421
rect 12571 26365 12657 26421
rect 12713 26365 12799 26421
rect 12855 26365 12941 26421
rect 12997 26365 13083 26421
rect 13139 26365 13225 26421
rect 13281 26365 13367 26421
rect 13423 26365 13509 26421
rect 13565 26365 13651 26421
rect 13707 26365 13793 26421
rect 13849 26365 13935 26421
rect 13991 26365 14077 26421
rect 14133 26365 14219 26421
rect 14275 26365 14361 26421
rect 14417 26365 14503 26421
rect 14559 26365 14645 26421
rect 14701 26365 14787 26421
rect 14843 26365 14853 26421
rect 151 26279 14853 26365
rect 151 26223 161 26279
rect 217 26223 303 26279
rect 359 26223 445 26279
rect 501 26223 587 26279
rect 643 26223 729 26279
rect 785 26223 871 26279
rect 927 26223 1013 26279
rect 1069 26223 1155 26279
rect 1211 26223 1297 26279
rect 1353 26223 1439 26279
rect 1495 26223 1581 26279
rect 1637 26223 1723 26279
rect 1779 26223 1865 26279
rect 1921 26223 2007 26279
rect 2063 26223 2149 26279
rect 2205 26223 2291 26279
rect 2347 26223 2433 26279
rect 2489 26223 2575 26279
rect 2631 26223 2717 26279
rect 2773 26223 2859 26279
rect 2915 26223 3001 26279
rect 3057 26223 3143 26279
rect 3199 26223 3285 26279
rect 3341 26223 3427 26279
rect 3483 26223 3569 26279
rect 3625 26223 3711 26279
rect 3767 26223 3853 26279
rect 3909 26223 3995 26279
rect 4051 26223 4137 26279
rect 4193 26223 4279 26279
rect 4335 26223 4421 26279
rect 4477 26223 4563 26279
rect 4619 26223 4705 26279
rect 4761 26223 4847 26279
rect 4903 26223 4989 26279
rect 5045 26223 5131 26279
rect 5187 26223 5273 26279
rect 5329 26223 5415 26279
rect 5471 26223 5557 26279
rect 5613 26223 5699 26279
rect 5755 26223 5841 26279
rect 5897 26223 5983 26279
rect 6039 26223 6125 26279
rect 6181 26223 6267 26279
rect 6323 26223 6409 26279
rect 6465 26223 6551 26279
rect 6607 26223 6693 26279
rect 6749 26223 6835 26279
rect 6891 26223 6977 26279
rect 7033 26223 7119 26279
rect 7175 26223 7261 26279
rect 7317 26223 7403 26279
rect 7459 26223 7545 26279
rect 7601 26223 7687 26279
rect 7743 26223 7829 26279
rect 7885 26223 7971 26279
rect 8027 26223 8113 26279
rect 8169 26223 8255 26279
rect 8311 26223 8397 26279
rect 8453 26223 8539 26279
rect 8595 26223 8681 26279
rect 8737 26223 8823 26279
rect 8879 26223 8965 26279
rect 9021 26223 9107 26279
rect 9163 26223 9249 26279
rect 9305 26223 9391 26279
rect 9447 26223 9533 26279
rect 9589 26223 9675 26279
rect 9731 26223 9817 26279
rect 9873 26223 9959 26279
rect 10015 26223 10101 26279
rect 10157 26223 10243 26279
rect 10299 26223 10385 26279
rect 10441 26223 10527 26279
rect 10583 26223 10669 26279
rect 10725 26223 10811 26279
rect 10867 26223 10953 26279
rect 11009 26223 11095 26279
rect 11151 26223 11237 26279
rect 11293 26223 11379 26279
rect 11435 26223 11521 26279
rect 11577 26223 11663 26279
rect 11719 26223 11805 26279
rect 11861 26223 11947 26279
rect 12003 26223 12089 26279
rect 12145 26223 12231 26279
rect 12287 26223 12373 26279
rect 12429 26223 12515 26279
rect 12571 26223 12657 26279
rect 12713 26223 12799 26279
rect 12855 26223 12941 26279
rect 12997 26223 13083 26279
rect 13139 26223 13225 26279
rect 13281 26223 13367 26279
rect 13423 26223 13509 26279
rect 13565 26223 13651 26279
rect 13707 26223 13793 26279
rect 13849 26223 13935 26279
rect 13991 26223 14077 26279
rect 14133 26223 14219 26279
rect 14275 26223 14361 26279
rect 14417 26223 14503 26279
rect 14559 26223 14645 26279
rect 14701 26223 14787 26279
rect 14843 26223 14853 26279
rect 151 26137 14853 26223
rect 151 26081 161 26137
rect 217 26081 303 26137
rect 359 26081 445 26137
rect 501 26081 587 26137
rect 643 26081 729 26137
rect 785 26081 871 26137
rect 927 26081 1013 26137
rect 1069 26081 1155 26137
rect 1211 26081 1297 26137
rect 1353 26081 1439 26137
rect 1495 26081 1581 26137
rect 1637 26081 1723 26137
rect 1779 26081 1865 26137
rect 1921 26081 2007 26137
rect 2063 26081 2149 26137
rect 2205 26081 2291 26137
rect 2347 26081 2433 26137
rect 2489 26081 2575 26137
rect 2631 26081 2717 26137
rect 2773 26081 2859 26137
rect 2915 26081 3001 26137
rect 3057 26081 3143 26137
rect 3199 26081 3285 26137
rect 3341 26081 3427 26137
rect 3483 26081 3569 26137
rect 3625 26081 3711 26137
rect 3767 26081 3853 26137
rect 3909 26081 3995 26137
rect 4051 26081 4137 26137
rect 4193 26081 4279 26137
rect 4335 26081 4421 26137
rect 4477 26081 4563 26137
rect 4619 26081 4705 26137
rect 4761 26081 4847 26137
rect 4903 26081 4989 26137
rect 5045 26081 5131 26137
rect 5187 26081 5273 26137
rect 5329 26081 5415 26137
rect 5471 26081 5557 26137
rect 5613 26081 5699 26137
rect 5755 26081 5841 26137
rect 5897 26081 5983 26137
rect 6039 26081 6125 26137
rect 6181 26081 6267 26137
rect 6323 26081 6409 26137
rect 6465 26081 6551 26137
rect 6607 26081 6693 26137
rect 6749 26081 6835 26137
rect 6891 26081 6977 26137
rect 7033 26081 7119 26137
rect 7175 26081 7261 26137
rect 7317 26081 7403 26137
rect 7459 26081 7545 26137
rect 7601 26081 7687 26137
rect 7743 26081 7829 26137
rect 7885 26081 7971 26137
rect 8027 26081 8113 26137
rect 8169 26081 8255 26137
rect 8311 26081 8397 26137
rect 8453 26081 8539 26137
rect 8595 26081 8681 26137
rect 8737 26081 8823 26137
rect 8879 26081 8965 26137
rect 9021 26081 9107 26137
rect 9163 26081 9249 26137
rect 9305 26081 9391 26137
rect 9447 26081 9533 26137
rect 9589 26081 9675 26137
rect 9731 26081 9817 26137
rect 9873 26081 9959 26137
rect 10015 26081 10101 26137
rect 10157 26081 10243 26137
rect 10299 26081 10385 26137
rect 10441 26081 10527 26137
rect 10583 26081 10669 26137
rect 10725 26081 10811 26137
rect 10867 26081 10953 26137
rect 11009 26081 11095 26137
rect 11151 26081 11237 26137
rect 11293 26081 11379 26137
rect 11435 26081 11521 26137
rect 11577 26081 11663 26137
rect 11719 26081 11805 26137
rect 11861 26081 11947 26137
rect 12003 26081 12089 26137
rect 12145 26081 12231 26137
rect 12287 26081 12373 26137
rect 12429 26081 12515 26137
rect 12571 26081 12657 26137
rect 12713 26081 12799 26137
rect 12855 26081 12941 26137
rect 12997 26081 13083 26137
rect 13139 26081 13225 26137
rect 13281 26081 13367 26137
rect 13423 26081 13509 26137
rect 13565 26081 13651 26137
rect 13707 26081 13793 26137
rect 13849 26081 13935 26137
rect 13991 26081 14077 26137
rect 14133 26081 14219 26137
rect 14275 26081 14361 26137
rect 14417 26081 14503 26137
rect 14559 26081 14645 26137
rect 14701 26081 14787 26137
rect 14843 26081 14853 26137
rect 151 25995 14853 26081
rect 151 25939 161 25995
rect 217 25939 303 25995
rect 359 25939 445 25995
rect 501 25939 587 25995
rect 643 25939 729 25995
rect 785 25939 871 25995
rect 927 25939 1013 25995
rect 1069 25939 1155 25995
rect 1211 25939 1297 25995
rect 1353 25939 1439 25995
rect 1495 25939 1581 25995
rect 1637 25939 1723 25995
rect 1779 25939 1865 25995
rect 1921 25939 2007 25995
rect 2063 25939 2149 25995
rect 2205 25939 2291 25995
rect 2347 25939 2433 25995
rect 2489 25939 2575 25995
rect 2631 25939 2717 25995
rect 2773 25939 2859 25995
rect 2915 25939 3001 25995
rect 3057 25939 3143 25995
rect 3199 25939 3285 25995
rect 3341 25939 3427 25995
rect 3483 25939 3569 25995
rect 3625 25939 3711 25995
rect 3767 25939 3853 25995
rect 3909 25939 3995 25995
rect 4051 25939 4137 25995
rect 4193 25939 4279 25995
rect 4335 25939 4421 25995
rect 4477 25939 4563 25995
rect 4619 25939 4705 25995
rect 4761 25939 4847 25995
rect 4903 25939 4989 25995
rect 5045 25939 5131 25995
rect 5187 25939 5273 25995
rect 5329 25939 5415 25995
rect 5471 25939 5557 25995
rect 5613 25939 5699 25995
rect 5755 25939 5841 25995
rect 5897 25939 5983 25995
rect 6039 25939 6125 25995
rect 6181 25939 6267 25995
rect 6323 25939 6409 25995
rect 6465 25939 6551 25995
rect 6607 25939 6693 25995
rect 6749 25939 6835 25995
rect 6891 25939 6977 25995
rect 7033 25939 7119 25995
rect 7175 25939 7261 25995
rect 7317 25939 7403 25995
rect 7459 25939 7545 25995
rect 7601 25939 7687 25995
rect 7743 25939 7829 25995
rect 7885 25939 7971 25995
rect 8027 25939 8113 25995
rect 8169 25939 8255 25995
rect 8311 25939 8397 25995
rect 8453 25939 8539 25995
rect 8595 25939 8681 25995
rect 8737 25939 8823 25995
rect 8879 25939 8965 25995
rect 9021 25939 9107 25995
rect 9163 25939 9249 25995
rect 9305 25939 9391 25995
rect 9447 25939 9533 25995
rect 9589 25939 9675 25995
rect 9731 25939 9817 25995
rect 9873 25939 9959 25995
rect 10015 25939 10101 25995
rect 10157 25939 10243 25995
rect 10299 25939 10385 25995
rect 10441 25939 10527 25995
rect 10583 25939 10669 25995
rect 10725 25939 10811 25995
rect 10867 25939 10953 25995
rect 11009 25939 11095 25995
rect 11151 25939 11237 25995
rect 11293 25939 11379 25995
rect 11435 25939 11521 25995
rect 11577 25939 11663 25995
rect 11719 25939 11805 25995
rect 11861 25939 11947 25995
rect 12003 25939 12089 25995
rect 12145 25939 12231 25995
rect 12287 25939 12373 25995
rect 12429 25939 12515 25995
rect 12571 25939 12657 25995
rect 12713 25939 12799 25995
rect 12855 25939 12941 25995
rect 12997 25939 13083 25995
rect 13139 25939 13225 25995
rect 13281 25939 13367 25995
rect 13423 25939 13509 25995
rect 13565 25939 13651 25995
rect 13707 25939 13793 25995
rect 13849 25939 13935 25995
rect 13991 25939 14077 25995
rect 14133 25939 14219 25995
rect 14275 25939 14361 25995
rect 14417 25939 14503 25995
rect 14559 25939 14645 25995
rect 14701 25939 14787 25995
rect 14843 25939 14853 25995
rect 151 25853 14853 25939
rect 151 25797 161 25853
rect 217 25797 303 25853
rect 359 25797 445 25853
rect 501 25797 587 25853
rect 643 25797 729 25853
rect 785 25797 871 25853
rect 927 25797 1013 25853
rect 1069 25797 1155 25853
rect 1211 25797 1297 25853
rect 1353 25797 1439 25853
rect 1495 25797 1581 25853
rect 1637 25797 1723 25853
rect 1779 25797 1865 25853
rect 1921 25797 2007 25853
rect 2063 25797 2149 25853
rect 2205 25797 2291 25853
rect 2347 25797 2433 25853
rect 2489 25797 2575 25853
rect 2631 25797 2717 25853
rect 2773 25797 2859 25853
rect 2915 25797 3001 25853
rect 3057 25797 3143 25853
rect 3199 25797 3285 25853
rect 3341 25797 3427 25853
rect 3483 25797 3569 25853
rect 3625 25797 3711 25853
rect 3767 25797 3853 25853
rect 3909 25797 3995 25853
rect 4051 25797 4137 25853
rect 4193 25797 4279 25853
rect 4335 25797 4421 25853
rect 4477 25797 4563 25853
rect 4619 25797 4705 25853
rect 4761 25797 4847 25853
rect 4903 25797 4989 25853
rect 5045 25797 5131 25853
rect 5187 25797 5273 25853
rect 5329 25797 5415 25853
rect 5471 25797 5557 25853
rect 5613 25797 5699 25853
rect 5755 25797 5841 25853
rect 5897 25797 5983 25853
rect 6039 25797 6125 25853
rect 6181 25797 6267 25853
rect 6323 25797 6409 25853
rect 6465 25797 6551 25853
rect 6607 25797 6693 25853
rect 6749 25797 6835 25853
rect 6891 25797 6977 25853
rect 7033 25797 7119 25853
rect 7175 25797 7261 25853
rect 7317 25797 7403 25853
rect 7459 25797 7545 25853
rect 7601 25797 7687 25853
rect 7743 25797 7829 25853
rect 7885 25797 7971 25853
rect 8027 25797 8113 25853
rect 8169 25797 8255 25853
rect 8311 25797 8397 25853
rect 8453 25797 8539 25853
rect 8595 25797 8681 25853
rect 8737 25797 8823 25853
rect 8879 25797 8965 25853
rect 9021 25797 9107 25853
rect 9163 25797 9249 25853
rect 9305 25797 9391 25853
rect 9447 25797 9533 25853
rect 9589 25797 9675 25853
rect 9731 25797 9817 25853
rect 9873 25797 9959 25853
rect 10015 25797 10101 25853
rect 10157 25797 10243 25853
rect 10299 25797 10385 25853
rect 10441 25797 10527 25853
rect 10583 25797 10669 25853
rect 10725 25797 10811 25853
rect 10867 25797 10953 25853
rect 11009 25797 11095 25853
rect 11151 25797 11237 25853
rect 11293 25797 11379 25853
rect 11435 25797 11521 25853
rect 11577 25797 11663 25853
rect 11719 25797 11805 25853
rect 11861 25797 11947 25853
rect 12003 25797 12089 25853
rect 12145 25797 12231 25853
rect 12287 25797 12373 25853
rect 12429 25797 12515 25853
rect 12571 25797 12657 25853
rect 12713 25797 12799 25853
rect 12855 25797 12941 25853
rect 12997 25797 13083 25853
rect 13139 25797 13225 25853
rect 13281 25797 13367 25853
rect 13423 25797 13509 25853
rect 13565 25797 13651 25853
rect 13707 25797 13793 25853
rect 13849 25797 13935 25853
rect 13991 25797 14077 25853
rect 14133 25797 14219 25853
rect 14275 25797 14361 25853
rect 14417 25797 14503 25853
rect 14559 25797 14645 25853
rect 14701 25797 14787 25853
rect 14843 25797 14853 25853
rect 151 25711 14853 25797
rect 151 25655 161 25711
rect 217 25655 303 25711
rect 359 25655 445 25711
rect 501 25655 587 25711
rect 643 25655 729 25711
rect 785 25655 871 25711
rect 927 25655 1013 25711
rect 1069 25655 1155 25711
rect 1211 25655 1297 25711
rect 1353 25655 1439 25711
rect 1495 25655 1581 25711
rect 1637 25655 1723 25711
rect 1779 25655 1865 25711
rect 1921 25655 2007 25711
rect 2063 25655 2149 25711
rect 2205 25655 2291 25711
rect 2347 25655 2433 25711
rect 2489 25655 2575 25711
rect 2631 25655 2717 25711
rect 2773 25655 2859 25711
rect 2915 25655 3001 25711
rect 3057 25655 3143 25711
rect 3199 25655 3285 25711
rect 3341 25655 3427 25711
rect 3483 25655 3569 25711
rect 3625 25655 3711 25711
rect 3767 25655 3853 25711
rect 3909 25655 3995 25711
rect 4051 25655 4137 25711
rect 4193 25655 4279 25711
rect 4335 25655 4421 25711
rect 4477 25655 4563 25711
rect 4619 25655 4705 25711
rect 4761 25655 4847 25711
rect 4903 25655 4989 25711
rect 5045 25655 5131 25711
rect 5187 25655 5273 25711
rect 5329 25655 5415 25711
rect 5471 25655 5557 25711
rect 5613 25655 5699 25711
rect 5755 25655 5841 25711
rect 5897 25655 5983 25711
rect 6039 25655 6125 25711
rect 6181 25655 6267 25711
rect 6323 25655 6409 25711
rect 6465 25655 6551 25711
rect 6607 25655 6693 25711
rect 6749 25655 6835 25711
rect 6891 25655 6977 25711
rect 7033 25655 7119 25711
rect 7175 25655 7261 25711
rect 7317 25655 7403 25711
rect 7459 25655 7545 25711
rect 7601 25655 7687 25711
rect 7743 25655 7829 25711
rect 7885 25655 7971 25711
rect 8027 25655 8113 25711
rect 8169 25655 8255 25711
rect 8311 25655 8397 25711
rect 8453 25655 8539 25711
rect 8595 25655 8681 25711
rect 8737 25655 8823 25711
rect 8879 25655 8965 25711
rect 9021 25655 9107 25711
rect 9163 25655 9249 25711
rect 9305 25655 9391 25711
rect 9447 25655 9533 25711
rect 9589 25655 9675 25711
rect 9731 25655 9817 25711
rect 9873 25655 9959 25711
rect 10015 25655 10101 25711
rect 10157 25655 10243 25711
rect 10299 25655 10385 25711
rect 10441 25655 10527 25711
rect 10583 25655 10669 25711
rect 10725 25655 10811 25711
rect 10867 25655 10953 25711
rect 11009 25655 11095 25711
rect 11151 25655 11237 25711
rect 11293 25655 11379 25711
rect 11435 25655 11521 25711
rect 11577 25655 11663 25711
rect 11719 25655 11805 25711
rect 11861 25655 11947 25711
rect 12003 25655 12089 25711
rect 12145 25655 12231 25711
rect 12287 25655 12373 25711
rect 12429 25655 12515 25711
rect 12571 25655 12657 25711
rect 12713 25655 12799 25711
rect 12855 25655 12941 25711
rect 12997 25655 13083 25711
rect 13139 25655 13225 25711
rect 13281 25655 13367 25711
rect 13423 25655 13509 25711
rect 13565 25655 13651 25711
rect 13707 25655 13793 25711
rect 13849 25655 13935 25711
rect 13991 25655 14077 25711
rect 14133 25655 14219 25711
rect 14275 25655 14361 25711
rect 14417 25655 14503 25711
rect 14559 25655 14645 25711
rect 14701 25655 14787 25711
rect 14843 25655 14853 25711
rect 151 25569 14853 25655
rect 151 25513 161 25569
rect 217 25513 303 25569
rect 359 25513 445 25569
rect 501 25513 587 25569
rect 643 25513 729 25569
rect 785 25513 871 25569
rect 927 25513 1013 25569
rect 1069 25513 1155 25569
rect 1211 25513 1297 25569
rect 1353 25513 1439 25569
rect 1495 25513 1581 25569
rect 1637 25513 1723 25569
rect 1779 25513 1865 25569
rect 1921 25513 2007 25569
rect 2063 25513 2149 25569
rect 2205 25513 2291 25569
rect 2347 25513 2433 25569
rect 2489 25513 2575 25569
rect 2631 25513 2717 25569
rect 2773 25513 2859 25569
rect 2915 25513 3001 25569
rect 3057 25513 3143 25569
rect 3199 25513 3285 25569
rect 3341 25513 3427 25569
rect 3483 25513 3569 25569
rect 3625 25513 3711 25569
rect 3767 25513 3853 25569
rect 3909 25513 3995 25569
rect 4051 25513 4137 25569
rect 4193 25513 4279 25569
rect 4335 25513 4421 25569
rect 4477 25513 4563 25569
rect 4619 25513 4705 25569
rect 4761 25513 4847 25569
rect 4903 25513 4989 25569
rect 5045 25513 5131 25569
rect 5187 25513 5273 25569
rect 5329 25513 5415 25569
rect 5471 25513 5557 25569
rect 5613 25513 5699 25569
rect 5755 25513 5841 25569
rect 5897 25513 5983 25569
rect 6039 25513 6125 25569
rect 6181 25513 6267 25569
rect 6323 25513 6409 25569
rect 6465 25513 6551 25569
rect 6607 25513 6693 25569
rect 6749 25513 6835 25569
rect 6891 25513 6977 25569
rect 7033 25513 7119 25569
rect 7175 25513 7261 25569
rect 7317 25513 7403 25569
rect 7459 25513 7545 25569
rect 7601 25513 7687 25569
rect 7743 25513 7829 25569
rect 7885 25513 7971 25569
rect 8027 25513 8113 25569
rect 8169 25513 8255 25569
rect 8311 25513 8397 25569
rect 8453 25513 8539 25569
rect 8595 25513 8681 25569
rect 8737 25513 8823 25569
rect 8879 25513 8965 25569
rect 9021 25513 9107 25569
rect 9163 25513 9249 25569
rect 9305 25513 9391 25569
rect 9447 25513 9533 25569
rect 9589 25513 9675 25569
rect 9731 25513 9817 25569
rect 9873 25513 9959 25569
rect 10015 25513 10101 25569
rect 10157 25513 10243 25569
rect 10299 25513 10385 25569
rect 10441 25513 10527 25569
rect 10583 25513 10669 25569
rect 10725 25513 10811 25569
rect 10867 25513 10953 25569
rect 11009 25513 11095 25569
rect 11151 25513 11237 25569
rect 11293 25513 11379 25569
rect 11435 25513 11521 25569
rect 11577 25513 11663 25569
rect 11719 25513 11805 25569
rect 11861 25513 11947 25569
rect 12003 25513 12089 25569
rect 12145 25513 12231 25569
rect 12287 25513 12373 25569
rect 12429 25513 12515 25569
rect 12571 25513 12657 25569
rect 12713 25513 12799 25569
rect 12855 25513 12941 25569
rect 12997 25513 13083 25569
rect 13139 25513 13225 25569
rect 13281 25513 13367 25569
rect 13423 25513 13509 25569
rect 13565 25513 13651 25569
rect 13707 25513 13793 25569
rect 13849 25513 13935 25569
rect 13991 25513 14077 25569
rect 14133 25513 14219 25569
rect 14275 25513 14361 25569
rect 14417 25513 14503 25569
rect 14559 25513 14645 25569
rect 14701 25513 14787 25569
rect 14843 25513 14853 25569
rect 151 25427 14853 25513
rect 151 25371 161 25427
rect 217 25371 303 25427
rect 359 25371 445 25427
rect 501 25371 587 25427
rect 643 25371 729 25427
rect 785 25371 871 25427
rect 927 25371 1013 25427
rect 1069 25371 1155 25427
rect 1211 25371 1297 25427
rect 1353 25371 1439 25427
rect 1495 25371 1581 25427
rect 1637 25371 1723 25427
rect 1779 25371 1865 25427
rect 1921 25371 2007 25427
rect 2063 25371 2149 25427
rect 2205 25371 2291 25427
rect 2347 25371 2433 25427
rect 2489 25371 2575 25427
rect 2631 25371 2717 25427
rect 2773 25371 2859 25427
rect 2915 25371 3001 25427
rect 3057 25371 3143 25427
rect 3199 25371 3285 25427
rect 3341 25371 3427 25427
rect 3483 25371 3569 25427
rect 3625 25371 3711 25427
rect 3767 25371 3853 25427
rect 3909 25371 3995 25427
rect 4051 25371 4137 25427
rect 4193 25371 4279 25427
rect 4335 25371 4421 25427
rect 4477 25371 4563 25427
rect 4619 25371 4705 25427
rect 4761 25371 4847 25427
rect 4903 25371 4989 25427
rect 5045 25371 5131 25427
rect 5187 25371 5273 25427
rect 5329 25371 5415 25427
rect 5471 25371 5557 25427
rect 5613 25371 5699 25427
rect 5755 25371 5841 25427
rect 5897 25371 5983 25427
rect 6039 25371 6125 25427
rect 6181 25371 6267 25427
rect 6323 25371 6409 25427
rect 6465 25371 6551 25427
rect 6607 25371 6693 25427
rect 6749 25371 6835 25427
rect 6891 25371 6977 25427
rect 7033 25371 7119 25427
rect 7175 25371 7261 25427
rect 7317 25371 7403 25427
rect 7459 25371 7545 25427
rect 7601 25371 7687 25427
rect 7743 25371 7829 25427
rect 7885 25371 7971 25427
rect 8027 25371 8113 25427
rect 8169 25371 8255 25427
rect 8311 25371 8397 25427
rect 8453 25371 8539 25427
rect 8595 25371 8681 25427
rect 8737 25371 8823 25427
rect 8879 25371 8965 25427
rect 9021 25371 9107 25427
rect 9163 25371 9249 25427
rect 9305 25371 9391 25427
rect 9447 25371 9533 25427
rect 9589 25371 9675 25427
rect 9731 25371 9817 25427
rect 9873 25371 9959 25427
rect 10015 25371 10101 25427
rect 10157 25371 10243 25427
rect 10299 25371 10385 25427
rect 10441 25371 10527 25427
rect 10583 25371 10669 25427
rect 10725 25371 10811 25427
rect 10867 25371 10953 25427
rect 11009 25371 11095 25427
rect 11151 25371 11237 25427
rect 11293 25371 11379 25427
rect 11435 25371 11521 25427
rect 11577 25371 11663 25427
rect 11719 25371 11805 25427
rect 11861 25371 11947 25427
rect 12003 25371 12089 25427
rect 12145 25371 12231 25427
rect 12287 25371 12373 25427
rect 12429 25371 12515 25427
rect 12571 25371 12657 25427
rect 12713 25371 12799 25427
rect 12855 25371 12941 25427
rect 12997 25371 13083 25427
rect 13139 25371 13225 25427
rect 13281 25371 13367 25427
rect 13423 25371 13509 25427
rect 13565 25371 13651 25427
rect 13707 25371 13793 25427
rect 13849 25371 13935 25427
rect 13991 25371 14077 25427
rect 14133 25371 14219 25427
rect 14275 25371 14361 25427
rect 14417 25371 14503 25427
rect 14559 25371 14645 25427
rect 14701 25371 14787 25427
rect 14843 25371 14853 25427
rect 151 25285 14853 25371
rect 151 25229 161 25285
rect 217 25229 303 25285
rect 359 25229 445 25285
rect 501 25229 587 25285
rect 643 25229 729 25285
rect 785 25229 871 25285
rect 927 25229 1013 25285
rect 1069 25229 1155 25285
rect 1211 25229 1297 25285
rect 1353 25229 1439 25285
rect 1495 25229 1581 25285
rect 1637 25229 1723 25285
rect 1779 25229 1865 25285
rect 1921 25229 2007 25285
rect 2063 25229 2149 25285
rect 2205 25229 2291 25285
rect 2347 25229 2433 25285
rect 2489 25229 2575 25285
rect 2631 25229 2717 25285
rect 2773 25229 2859 25285
rect 2915 25229 3001 25285
rect 3057 25229 3143 25285
rect 3199 25229 3285 25285
rect 3341 25229 3427 25285
rect 3483 25229 3569 25285
rect 3625 25229 3711 25285
rect 3767 25229 3853 25285
rect 3909 25229 3995 25285
rect 4051 25229 4137 25285
rect 4193 25229 4279 25285
rect 4335 25229 4421 25285
rect 4477 25229 4563 25285
rect 4619 25229 4705 25285
rect 4761 25229 4847 25285
rect 4903 25229 4989 25285
rect 5045 25229 5131 25285
rect 5187 25229 5273 25285
rect 5329 25229 5415 25285
rect 5471 25229 5557 25285
rect 5613 25229 5699 25285
rect 5755 25229 5841 25285
rect 5897 25229 5983 25285
rect 6039 25229 6125 25285
rect 6181 25229 6267 25285
rect 6323 25229 6409 25285
rect 6465 25229 6551 25285
rect 6607 25229 6693 25285
rect 6749 25229 6835 25285
rect 6891 25229 6977 25285
rect 7033 25229 7119 25285
rect 7175 25229 7261 25285
rect 7317 25229 7403 25285
rect 7459 25229 7545 25285
rect 7601 25229 7687 25285
rect 7743 25229 7829 25285
rect 7885 25229 7971 25285
rect 8027 25229 8113 25285
rect 8169 25229 8255 25285
rect 8311 25229 8397 25285
rect 8453 25229 8539 25285
rect 8595 25229 8681 25285
rect 8737 25229 8823 25285
rect 8879 25229 8965 25285
rect 9021 25229 9107 25285
rect 9163 25229 9249 25285
rect 9305 25229 9391 25285
rect 9447 25229 9533 25285
rect 9589 25229 9675 25285
rect 9731 25229 9817 25285
rect 9873 25229 9959 25285
rect 10015 25229 10101 25285
rect 10157 25229 10243 25285
rect 10299 25229 10385 25285
rect 10441 25229 10527 25285
rect 10583 25229 10669 25285
rect 10725 25229 10811 25285
rect 10867 25229 10953 25285
rect 11009 25229 11095 25285
rect 11151 25229 11237 25285
rect 11293 25229 11379 25285
rect 11435 25229 11521 25285
rect 11577 25229 11663 25285
rect 11719 25229 11805 25285
rect 11861 25229 11947 25285
rect 12003 25229 12089 25285
rect 12145 25229 12231 25285
rect 12287 25229 12373 25285
rect 12429 25229 12515 25285
rect 12571 25229 12657 25285
rect 12713 25229 12799 25285
rect 12855 25229 12941 25285
rect 12997 25229 13083 25285
rect 13139 25229 13225 25285
rect 13281 25229 13367 25285
rect 13423 25229 13509 25285
rect 13565 25229 13651 25285
rect 13707 25229 13793 25285
rect 13849 25229 13935 25285
rect 13991 25229 14077 25285
rect 14133 25229 14219 25285
rect 14275 25229 14361 25285
rect 14417 25229 14503 25285
rect 14559 25229 14645 25285
rect 14701 25229 14787 25285
rect 14843 25229 14853 25285
rect 151 25219 14853 25229
rect 151 24963 14853 24973
rect 151 24907 161 24963
rect 217 24907 303 24963
rect 359 24907 445 24963
rect 501 24907 587 24963
rect 643 24907 729 24963
rect 785 24907 871 24963
rect 927 24907 1013 24963
rect 1069 24907 1155 24963
rect 1211 24907 1297 24963
rect 1353 24907 1439 24963
rect 1495 24907 1581 24963
rect 1637 24907 1723 24963
rect 1779 24907 1865 24963
rect 1921 24907 2007 24963
rect 2063 24907 2149 24963
rect 2205 24907 2291 24963
rect 2347 24907 2433 24963
rect 2489 24907 2575 24963
rect 2631 24907 2717 24963
rect 2773 24907 2859 24963
rect 2915 24907 3001 24963
rect 3057 24907 3143 24963
rect 3199 24907 3285 24963
rect 3341 24907 3427 24963
rect 3483 24907 3569 24963
rect 3625 24907 3711 24963
rect 3767 24907 3853 24963
rect 3909 24907 3995 24963
rect 4051 24907 4137 24963
rect 4193 24907 4279 24963
rect 4335 24907 4421 24963
rect 4477 24907 4563 24963
rect 4619 24907 4705 24963
rect 4761 24907 4847 24963
rect 4903 24907 4989 24963
rect 5045 24907 5131 24963
rect 5187 24907 5273 24963
rect 5329 24907 5415 24963
rect 5471 24907 5557 24963
rect 5613 24907 5699 24963
rect 5755 24907 5841 24963
rect 5897 24907 5983 24963
rect 6039 24907 6125 24963
rect 6181 24907 6267 24963
rect 6323 24907 6409 24963
rect 6465 24907 6551 24963
rect 6607 24907 6693 24963
rect 6749 24907 6835 24963
rect 6891 24907 6977 24963
rect 7033 24907 7119 24963
rect 7175 24907 7261 24963
rect 7317 24907 7403 24963
rect 7459 24907 7545 24963
rect 7601 24907 7687 24963
rect 7743 24907 7829 24963
rect 7885 24907 7971 24963
rect 8027 24907 8113 24963
rect 8169 24907 8255 24963
rect 8311 24907 8397 24963
rect 8453 24907 8539 24963
rect 8595 24907 8681 24963
rect 8737 24907 8823 24963
rect 8879 24907 8965 24963
rect 9021 24907 9107 24963
rect 9163 24907 9249 24963
rect 9305 24907 9391 24963
rect 9447 24907 9533 24963
rect 9589 24907 9675 24963
rect 9731 24907 9817 24963
rect 9873 24907 9959 24963
rect 10015 24907 10101 24963
rect 10157 24907 10243 24963
rect 10299 24907 10385 24963
rect 10441 24907 10527 24963
rect 10583 24907 10669 24963
rect 10725 24907 10811 24963
rect 10867 24907 10953 24963
rect 11009 24907 11095 24963
rect 11151 24907 11237 24963
rect 11293 24907 11379 24963
rect 11435 24907 11521 24963
rect 11577 24907 11663 24963
rect 11719 24907 11805 24963
rect 11861 24907 11947 24963
rect 12003 24907 12089 24963
rect 12145 24907 12231 24963
rect 12287 24907 12373 24963
rect 12429 24907 12515 24963
rect 12571 24907 12657 24963
rect 12713 24907 12799 24963
rect 12855 24907 12941 24963
rect 12997 24907 13083 24963
rect 13139 24907 13225 24963
rect 13281 24907 13367 24963
rect 13423 24907 13509 24963
rect 13565 24907 13651 24963
rect 13707 24907 13793 24963
rect 13849 24907 13935 24963
rect 13991 24907 14077 24963
rect 14133 24907 14219 24963
rect 14275 24907 14361 24963
rect 14417 24907 14503 24963
rect 14559 24907 14645 24963
rect 14701 24907 14787 24963
rect 14843 24907 14853 24963
rect 151 24821 14853 24907
rect 151 24765 161 24821
rect 217 24765 303 24821
rect 359 24765 445 24821
rect 501 24765 587 24821
rect 643 24765 729 24821
rect 785 24765 871 24821
rect 927 24765 1013 24821
rect 1069 24765 1155 24821
rect 1211 24765 1297 24821
rect 1353 24765 1439 24821
rect 1495 24765 1581 24821
rect 1637 24765 1723 24821
rect 1779 24765 1865 24821
rect 1921 24765 2007 24821
rect 2063 24765 2149 24821
rect 2205 24765 2291 24821
rect 2347 24765 2433 24821
rect 2489 24765 2575 24821
rect 2631 24765 2717 24821
rect 2773 24765 2859 24821
rect 2915 24765 3001 24821
rect 3057 24765 3143 24821
rect 3199 24765 3285 24821
rect 3341 24765 3427 24821
rect 3483 24765 3569 24821
rect 3625 24765 3711 24821
rect 3767 24765 3853 24821
rect 3909 24765 3995 24821
rect 4051 24765 4137 24821
rect 4193 24765 4279 24821
rect 4335 24765 4421 24821
rect 4477 24765 4563 24821
rect 4619 24765 4705 24821
rect 4761 24765 4847 24821
rect 4903 24765 4989 24821
rect 5045 24765 5131 24821
rect 5187 24765 5273 24821
rect 5329 24765 5415 24821
rect 5471 24765 5557 24821
rect 5613 24765 5699 24821
rect 5755 24765 5841 24821
rect 5897 24765 5983 24821
rect 6039 24765 6125 24821
rect 6181 24765 6267 24821
rect 6323 24765 6409 24821
rect 6465 24765 6551 24821
rect 6607 24765 6693 24821
rect 6749 24765 6835 24821
rect 6891 24765 6977 24821
rect 7033 24765 7119 24821
rect 7175 24765 7261 24821
rect 7317 24765 7403 24821
rect 7459 24765 7545 24821
rect 7601 24765 7687 24821
rect 7743 24765 7829 24821
rect 7885 24765 7971 24821
rect 8027 24765 8113 24821
rect 8169 24765 8255 24821
rect 8311 24765 8397 24821
rect 8453 24765 8539 24821
rect 8595 24765 8681 24821
rect 8737 24765 8823 24821
rect 8879 24765 8965 24821
rect 9021 24765 9107 24821
rect 9163 24765 9249 24821
rect 9305 24765 9391 24821
rect 9447 24765 9533 24821
rect 9589 24765 9675 24821
rect 9731 24765 9817 24821
rect 9873 24765 9959 24821
rect 10015 24765 10101 24821
rect 10157 24765 10243 24821
rect 10299 24765 10385 24821
rect 10441 24765 10527 24821
rect 10583 24765 10669 24821
rect 10725 24765 10811 24821
rect 10867 24765 10953 24821
rect 11009 24765 11095 24821
rect 11151 24765 11237 24821
rect 11293 24765 11379 24821
rect 11435 24765 11521 24821
rect 11577 24765 11663 24821
rect 11719 24765 11805 24821
rect 11861 24765 11947 24821
rect 12003 24765 12089 24821
rect 12145 24765 12231 24821
rect 12287 24765 12373 24821
rect 12429 24765 12515 24821
rect 12571 24765 12657 24821
rect 12713 24765 12799 24821
rect 12855 24765 12941 24821
rect 12997 24765 13083 24821
rect 13139 24765 13225 24821
rect 13281 24765 13367 24821
rect 13423 24765 13509 24821
rect 13565 24765 13651 24821
rect 13707 24765 13793 24821
rect 13849 24765 13935 24821
rect 13991 24765 14077 24821
rect 14133 24765 14219 24821
rect 14275 24765 14361 24821
rect 14417 24765 14503 24821
rect 14559 24765 14645 24821
rect 14701 24765 14787 24821
rect 14843 24765 14853 24821
rect 151 24679 14853 24765
rect 151 24623 161 24679
rect 217 24623 303 24679
rect 359 24623 445 24679
rect 501 24623 587 24679
rect 643 24623 729 24679
rect 785 24623 871 24679
rect 927 24623 1013 24679
rect 1069 24623 1155 24679
rect 1211 24623 1297 24679
rect 1353 24623 1439 24679
rect 1495 24623 1581 24679
rect 1637 24623 1723 24679
rect 1779 24623 1865 24679
rect 1921 24623 2007 24679
rect 2063 24623 2149 24679
rect 2205 24623 2291 24679
rect 2347 24623 2433 24679
rect 2489 24623 2575 24679
rect 2631 24623 2717 24679
rect 2773 24623 2859 24679
rect 2915 24623 3001 24679
rect 3057 24623 3143 24679
rect 3199 24623 3285 24679
rect 3341 24623 3427 24679
rect 3483 24623 3569 24679
rect 3625 24623 3711 24679
rect 3767 24623 3853 24679
rect 3909 24623 3995 24679
rect 4051 24623 4137 24679
rect 4193 24623 4279 24679
rect 4335 24623 4421 24679
rect 4477 24623 4563 24679
rect 4619 24623 4705 24679
rect 4761 24623 4847 24679
rect 4903 24623 4989 24679
rect 5045 24623 5131 24679
rect 5187 24623 5273 24679
rect 5329 24623 5415 24679
rect 5471 24623 5557 24679
rect 5613 24623 5699 24679
rect 5755 24623 5841 24679
rect 5897 24623 5983 24679
rect 6039 24623 6125 24679
rect 6181 24623 6267 24679
rect 6323 24623 6409 24679
rect 6465 24623 6551 24679
rect 6607 24623 6693 24679
rect 6749 24623 6835 24679
rect 6891 24623 6977 24679
rect 7033 24623 7119 24679
rect 7175 24623 7261 24679
rect 7317 24623 7403 24679
rect 7459 24623 7545 24679
rect 7601 24623 7687 24679
rect 7743 24623 7829 24679
rect 7885 24623 7971 24679
rect 8027 24623 8113 24679
rect 8169 24623 8255 24679
rect 8311 24623 8397 24679
rect 8453 24623 8539 24679
rect 8595 24623 8681 24679
rect 8737 24623 8823 24679
rect 8879 24623 8965 24679
rect 9021 24623 9107 24679
rect 9163 24623 9249 24679
rect 9305 24623 9391 24679
rect 9447 24623 9533 24679
rect 9589 24623 9675 24679
rect 9731 24623 9817 24679
rect 9873 24623 9959 24679
rect 10015 24623 10101 24679
rect 10157 24623 10243 24679
rect 10299 24623 10385 24679
rect 10441 24623 10527 24679
rect 10583 24623 10669 24679
rect 10725 24623 10811 24679
rect 10867 24623 10953 24679
rect 11009 24623 11095 24679
rect 11151 24623 11237 24679
rect 11293 24623 11379 24679
rect 11435 24623 11521 24679
rect 11577 24623 11663 24679
rect 11719 24623 11805 24679
rect 11861 24623 11947 24679
rect 12003 24623 12089 24679
rect 12145 24623 12231 24679
rect 12287 24623 12373 24679
rect 12429 24623 12515 24679
rect 12571 24623 12657 24679
rect 12713 24623 12799 24679
rect 12855 24623 12941 24679
rect 12997 24623 13083 24679
rect 13139 24623 13225 24679
rect 13281 24623 13367 24679
rect 13423 24623 13509 24679
rect 13565 24623 13651 24679
rect 13707 24623 13793 24679
rect 13849 24623 13935 24679
rect 13991 24623 14077 24679
rect 14133 24623 14219 24679
rect 14275 24623 14361 24679
rect 14417 24623 14503 24679
rect 14559 24623 14645 24679
rect 14701 24623 14787 24679
rect 14843 24623 14853 24679
rect 151 24537 14853 24623
rect 151 24481 161 24537
rect 217 24481 303 24537
rect 359 24481 445 24537
rect 501 24481 587 24537
rect 643 24481 729 24537
rect 785 24481 871 24537
rect 927 24481 1013 24537
rect 1069 24481 1155 24537
rect 1211 24481 1297 24537
rect 1353 24481 1439 24537
rect 1495 24481 1581 24537
rect 1637 24481 1723 24537
rect 1779 24481 1865 24537
rect 1921 24481 2007 24537
rect 2063 24481 2149 24537
rect 2205 24481 2291 24537
rect 2347 24481 2433 24537
rect 2489 24481 2575 24537
rect 2631 24481 2717 24537
rect 2773 24481 2859 24537
rect 2915 24481 3001 24537
rect 3057 24481 3143 24537
rect 3199 24481 3285 24537
rect 3341 24481 3427 24537
rect 3483 24481 3569 24537
rect 3625 24481 3711 24537
rect 3767 24481 3853 24537
rect 3909 24481 3995 24537
rect 4051 24481 4137 24537
rect 4193 24481 4279 24537
rect 4335 24481 4421 24537
rect 4477 24481 4563 24537
rect 4619 24481 4705 24537
rect 4761 24481 4847 24537
rect 4903 24481 4989 24537
rect 5045 24481 5131 24537
rect 5187 24481 5273 24537
rect 5329 24481 5415 24537
rect 5471 24481 5557 24537
rect 5613 24481 5699 24537
rect 5755 24481 5841 24537
rect 5897 24481 5983 24537
rect 6039 24481 6125 24537
rect 6181 24481 6267 24537
rect 6323 24481 6409 24537
rect 6465 24481 6551 24537
rect 6607 24481 6693 24537
rect 6749 24481 6835 24537
rect 6891 24481 6977 24537
rect 7033 24481 7119 24537
rect 7175 24481 7261 24537
rect 7317 24481 7403 24537
rect 7459 24481 7545 24537
rect 7601 24481 7687 24537
rect 7743 24481 7829 24537
rect 7885 24481 7971 24537
rect 8027 24481 8113 24537
rect 8169 24481 8255 24537
rect 8311 24481 8397 24537
rect 8453 24481 8539 24537
rect 8595 24481 8681 24537
rect 8737 24481 8823 24537
rect 8879 24481 8965 24537
rect 9021 24481 9107 24537
rect 9163 24481 9249 24537
rect 9305 24481 9391 24537
rect 9447 24481 9533 24537
rect 9589 24481 9675 24537
rect 9731 24481 9817 24537
rect 9873 24481 9959 24537
rect 10015 24481 10101 24537
rect 10157 24481 10243 24537
rect 10299 24481 10385 24537
rect 10441 24481 10527 24537
rect 10583 24481 10669 24537
rect 10725 24481 10811 24537
rect 10867 24481 10953 24537
rect 11009 24481 11095 24537
rect 11151 24481 11237 24537
rect 11293 24481 11379 24537
rect 11435 24481 11521 24537
rect 11577 24481 11663 24537
rect 11719 24481 11805 24537
rect 11861 24481 11947 24537
rect 12003 24481 12089 24537
rect 12145 24481 12231 24537
rect 12287 24481 12373 24537
rect 12429 24481 12515 24537
rect 12571 24481 12657 24537
rect 12713 24481 12799 24537
rect 12855 24481 12941 24537
rect 12997 24481 13083 24537
rect 13139 24481 13225 24537
rect 13281 24481 13367 24537
rect 13423 24481 13509 24537
rect 13565 24481 13651 24537
rect 13707 24481 13793 24537
rect 13849 24481 13935 24537
rect 13991 24481 14077 24537
rect 14133 24481 14219 24537
rect 14275 24481 14361 24537
rect 14417 24481 14503 24537
rect 14559 24481 14645 24537
rect 14701 24481 14787 24537
rect 14843 24481 14853 24537
rect 151 24395 14853 24481
rect 151 24339 161 24395
rect 217 24339 303 24395
rect 359 24339 445 24395
rect 501 24339 587 24395
rect 643 24339 729 24395
rect 785 24339 871 24395
rect 927 24339 1013 24395
rect 1069 24339 1155 24395
rect 1211 24339 1297 24395
rect 1353 24339 1439 24395
rect 1495 24339 1581 24395
rect 1637 24339 1723 24395
rect 1779 24339 1865 24395
rect 1921 24339 2007 24395
rect 2063 24339 2149 24395
rect 2205 24339 2291 24395
rect 2347 24339 2433 24395
rect 2489 24339 2575 24395
rect 2631 24339 2717 24395
rect 2773 24339 2859 24395
rect 2915 24339 3001 24395
rect 3057 24339 3143 24395
rect 3199 24339 3285 24395
rect 3341 24339 3427 24395
rect 3483 24339 3569 24395
rect 3625 24339 3711 24395
rect 3767 24339 3853 24395
rect 3909 24339 3995 24395
rect 4051 24339 4137 24395
rect 4193 24339 4279 24395
rect 4335 24339 4421 24395
rect 4477 24339 4563 24395
rect 4619 24339 4705 24395
rect 4761 24339 4847 24395
rect 4903 24339 4989 24395
rect 5045 24339 5131 24395
rect 5187 24339 5273 24395
rect 5329 24339 5415 24395
rect 5471 24339 5557 24395
rect 5613 24339 5699 24395
rect 5755 24339 5841 24395
rect 5897 24339 5983 24395
rect 6039 24339 6125 24395
rect 6181 24339 6267 24395
rect 6323 24339 6409 24395
rect 6465 24339 6551 24395
rect 6607 24339 6693 24395
rect 6749 24339 6835 24395
rect 6891 24339 6977 24395
rect 7033 24339 7119 24395
rect 7175 24339 7261 24395
rect 7317 24339 7403 24395
rect 7459 24339 7545 24395
rect 7601 24339 7687 24395
rect 7743 24339 7829 24395
rect 7885 24339 7971 24395
rect 8027 24339 8113 24395
rect 8169 24339 8255 24395
rect 8311 24339 8397 24395
rect 8453 24339 8539 24395
rect 8595 24339 8681 24395
rect 8737 24339 8823 24395
rect 8879 24339 8965 24395
rect 9021 24339 9107 24395
rect 9163 24339 9249 24395
rect 9305 24339 9391 24395
rect 9447 24339 9533 24395
rect 9589 24339 9675 24395
rect 9731 24339 9817 24395
rect 9873 24339 9959 24395
rect 10015 24339 10101 24395
rect 10157 24339 10243 24395
rect 10299 24339 10385 24395
rect 10441 24339 10527 24395
rect 10583 24339 10669 24395
rect 10725 24339 10811 24395
rect 10867 24339 10953 24395
rect 11009 24339 11095 24395
rect 11151 24339 11237 24395
rect 11293 24339 11379 24395
rect 11435 24339 11521 24395
rect 11577 24339 11663 24395
rect 11719 24339 11805 24395
rect 11861 24339 11947 24395
rect 12003 24339 12089 24395
rect 12145 24339 12231 24395
rect 12287 24339 12373 24395
rect 12429 24339 12515 24395
rect 12571 24339 12657 24395
rect 12713 24339 12799 24395
rect 12855 24339 12941 24395
rect 12997 24339 13083 24395
rect 13139 24339 13225 24395
rect 13281 24339 13367 24395
rect 13423 24339 13509 24395
rect 13565 24339 13651 24395
rect 13707 24339 13793 24395
rect 13849 24339 13935 24395
rect 13991 24339 14077 24395
rect 14133 24339 14219 24395
rect 14275 24339 14361 24395
rect 14417 24339 14503 24395
rect 14559 24339 14645 24395
rect 14701 24339 14787 24395
rect 14843 24339 14853 24395
rect 151 24253 14853 24339
rect 151 24197 161 24253
rect 217 24197 303 24253
rect 359 24197 445 24253
rect 501 24197 587 24253
rect 643 24197 729 24253
rect 785 24197 871 24253
rect 927 24197 1013 24253
rect 1069 24197 1155 24253
rect 1211 24197 1297 24253
rect 1353 24197 1439 24253
rect 1495 24197 1581 24253
rect 1637 24197 1723 24253
rect 1779 24197 1865 24253
rect 1921 24197 2007 24253
rect 2063 24197 2149 24253
rect 2205 24197 2291 24253
rect 2347 24197 2433 24253
rect 2489 24197 2575 24253
rect 2631 24197 2717 24253
rect 2773 24197 2859 24253
rect 2915 24197 3001 24253
rect 3057 24197 3143 24253
rect 3199 24197 3285 24253
rect 3341 24197 3427 24253
rect 3483 24197 3569 24253
rect 3625 24197 3711 24253
rect 3767 24197 3853 24253
rect 3909 24197 3995 24253
rect 4051 24197 4137 24253
rect 4193 24197 4279 24253
rect 4335 24197 4421 24253
rect 4477 24197 4563 24253
rect 4619 24197 4705 24253
rect 4761 24197 4847 24253
rect 4903 24197 4989 24253
rect 5045 24197 5131 24253
rect 5187 24197 5273 24253
rect 5329 24197 5415 24253
rect 5471 24197 5557 24253
rect 5613 24197 5699 24253
rect 5755 24197 5841 24253
rect 5897 24197 5983 24253
rect 6039 24197 6125 24253
rect 6181 24197 6267 24253
rect 6323 24197 6409 24253
rect 6465 24197 6551 24253
rect 6607 24197 6693 24253
rect 6749 24197 6835 24253
rect 6891 24197 6977 24253
rect 7033 24197 7119 24253
rect 7175 24197 7261 24253
rect 7317 24197 7403 24253
rect 7459 24197 7545 24253
rect 7601 24197 7687 24253
rect 7743 24197 7829 24253
rect 7885 24197 7971 24253
rect 8027 24197 8113 24253
rect 8169 24197 8255 24253
rect 8311 24197 8397 24253
rect 8453 24197 8539 24253
rect 8595 24197 8681 24253
rect 8737 24197 8823 24253
rect 8879 24197 8965 24253
rect 9021 24197 9107 24253
rect 9163 24197 9249 24253
rect 9305 24197 9391 24253
rect 9447 24197 9533 24253
rect 9589 24197 9675 24253
rect 9731 24197 9817 24253
rect 9873 24197 9959 24253
rect 10015 24197 10101 24253
rect 10157 24197 10243 24253
rect 10299 24197 10385 24253
rect 10441 24197 10527 24253
rect 10583 24197 10669 24253
rect 10725 24197 10811 24253
rect 10867 24197 10953 24253
rect 11009 24197 11095 24253
rect 11151 24197 11237 24253
rect 11293 24197 11379 24253
rect 11435 24197 11521 24253
rect 11577 24197 11663 24253
rect 11719 24197 11805 24253
rect 11861 24197 11947 24253
rect 12003 24197 12089 24253
rect 12145 24197 12231 24253
rect 12287 24197 12373 24253
rect 12429 24197 12515 24253
rect 12571 24197 12657 24253
rect 12713 24197 12799 24253
rect 12855 24197 12941 24253
rect 12997 24197 13083 24253
rect 13139 24197 13225 24253
rect 13281 24197 13367 24253
rect 13423 24197 13509 24253
rect 13565 24197 13651 24253
rect 13707 24197 13793 24253
rect 13849 24197 13935 24253
rect 13991 24197 14077 24253
rect 14133 24197 14219 24253
rect 14275 24197 14361 24253
rect 14417 24197 14503 24253
rect 14559 24197 14645 24253
rect 14701 24197 14787 24253
rect 14843 24197 14853 24253
rect 151 24111 14853 24197
rect 151 24055 161 24111
rect 217 24055 303 24111
rect 359 24055 445 24111
rect 501 24055 587 24111
rect 643 24055 729 24111
rect 785 24055 871 24111
rect 927 24055 1013 24111
rect 1069 24055 1155 24111
rect 1211 24055 1297 24111
rect 1353 24055 1439 24111
rect 1495 24055 1581 24111
rect 1637 24055 1723 24111
rect 1779 24055 1865 24111
rect 1921 24055 2007 24111
rect 2063 24055 2149 24111
rect 2205 24055 2291 24111
rect 2347 24055 2433 24111
rect 2489 24055 2575 24111
rect 2631 24055 2717 24111
rect 2773 24055 2859 24111
rect 2915 24055 3001 24111
rect 3057 24055 3143 24111
rect 3199 24055 3285 24111
rect 3341 24055 3427 24111
rect 3483 24055 3569 24111
rect 3625 24055 3711 24111
rect 3767 24055 3853 24111
rect 3909 24055 3995 24111
rect 4051 24055 4137 24111
rect 4193 24055 4279 24111
rect 4335 24055 4421 24111
rect 4477 24055 4563 24111
rect 4619 24055 4705 24111
rect 4761 24055 4847 24111
rect 4903 24055 4989 24111
rect 5045 24055 5131 24111
rect 5187 24055 5273 24111
rect 5329 24055 5415 24111
rect 5471 24055 5557 24111
rect 5613 24055 5699 24111
rect 5755 24055 5841 24111
rect 5897 24055 5983 24111
rect 6039 24055 6125 24111
rect 6181 24055 6267 24111
rect 6323 24055 6409 24111
rect 6465 24055 6551 24111
rect 6607 24055 6693 24111
rect 6749 24055 6835 24111
rect 6891 24055 6977 24111
rect 7033 24055 7119 24111
rect 7175 24055 7261 24111
rect 7317 24055 7403 24111
rect 7459 24055 7545 24111
rect 7601 24055 7687 24111
rect 7743 24055 7829 24111
rect 7885 24055 7971 24111
rect 8027 24055 8113 24111
rect 8169 24055 8255 24111
rect 8311 24055 8397 24111
rect 8453 24055 8539 24111
rect 8595 24055 8681 24111
rect 8737 24055 8823 24111
rect 8879 24055 8965 24111
rect 9021 24055 9107 24111
rect 9163 24055 9249 24111
rect 9305 24055 9391 24111
rect 9447 24055 9533 24111
rect 9589 24055 9675 24111
rect 9731 24055 9817 24111
rect 9873 24055 9959 24111
rect 10015 24055 10101 24111
rect 10157 24055 10243 24111
rect 10299 24055 10385 24111
rect 10441 24055 10527 24111
rect 10583 24055 10669 24111
rect 10725 24055 10811 24111
rect 10867 24055 10953 24111
rect 11009 24055 11095 24111
rect 11151 24055 11237 24111
rect 11293 24055 11379 24111
rect 11435 24055 11521 24111
rect 11577 24055 11663 24111
rect 11719 24055 11805 24111
rect 11861 24055 11947 24111
rect 12003 24055 12089 24111
rect 12145 24055 12231 24111
rect 12287 24055 12373 24111
rect 12429 24055 12515 24111
rect 12571 24055 12657 24111
rect 12713 24055 12799 24111
rect 12855 24055 12941 24111
rect 12997 24055 13083 24111
rect 13139 24055 13225 24111
rect 13281 24055 13367 24111
rect 13423 24055 13509 24111
rect 13565 24055 13651 24111
rect 13707 24055 13793 24111
rect 13849 24055 13935 24111
rect 13991 24055 14077 24111
rect 14133 24055 14219 24111
rect 14275 24055 14361 24111
rect 14417 24055 14503 24111
rect 14559 24055 14645 24111
rect 14701 24055 14787 24111
rect 14843 24055 14853 24111
rect 151 23969 14853 24055
rect 151 23913 161 23969
rect 217 23913 303 23969
rect 359 23913 445 23969
rect 501 23913 587 23969
rect 643 23913 729 23969
rect 785 23913 871 23969
rect 927 23913 1013 23969
rect 1069 23913 1155 23969
rect 1211 23913 1297 23969
rect 1353 23913 1439 23969
rect 1495 23913 1581 23969
rect 1637 23913 1723 23969
rect 1779 23913 1865 23969
rect 1921 23913 2007 23969
rect 2063 23913 2149 23969
rect 2205 23913 2291 23969
rect 2347 23913 2433 23969
rect 2489 23913 2575 23969
rect 2631 23913 2717 23969
rect 2773 23913 2859 23969
rect 2915 23913 3001 23969
rect 3057 23913 3143 23969
rect 3199 23913 3285 23969
rect 3341 23913 3427 23969
rect 3483 23913 3569 23969
rect 3625 23913 3711 23969
rect 3767 23913 3853 23969
rect 3909 23913 3995 23969
rect 4051 23913 4137 23969
rect 4193 23913 4279 23969
rect 4335 23913 4421 23969
rect 4477 23913 4563 23969
rect 4619 23913 4705 23969
rect 4761 23913 4847 23969
rect 4903 23913 4989 23969
rect 5045 23913 5131 23969
rect 5187 23913 5273 23969
rect 5329 23913 5415 23969
rect 5471 23913 5557 23969
rect 5613 23913 5699 23969
rect 5755 23913 5841 23969
rect 5897 23913 5983 23969
rect 6039 23913 6125 23969
rect 6181 23913 6267 23969
rect 6323 23913 6409 23969
rect 6465 23913 6551 23969
rect 6607 23913 6693 23969
rect 6749 23913 6835 23969
rect 6891 23913 6977 23969
rect 7033 23913 7119 23969
rect 7175 23913 7261 23969
rect 7317 23913 7403 23969
rect 7459 23913 7545 23969
rect 7601 23913 7687 23969
rect 7743 23913 7829 23969
rect 7885 23913 7971 23969
rect 8027 23913 8113 23969
rect 8169 23913 8255 23969
rect 8311 23913 8397 23969
rect 8453 23913 8539 23969
rect 8595 23913 8681 23969
rect 8737 23913 8823 23969
rect 8879 23913 8965 23969
rect 9021 23913 9107 23969
rect 9163 23913 9249 23969
rect 9305 23913 9391 23969
rect 9447 23913 9533 23969
rect 9589 23913 9675 23969
rect 9731 23913 9817 23969
rect 9873 23913 9959 23969
rect 10015 23913 10101 23969
rect 10157 23913 10243 23969
rect 10299 23913 10385 23969
rect 10441 23913 10527 23969
rect 10583 23913 10669 23969
rect 10725 23913 10811 23969
rect 10867 23913 10953 23969
rect 11009 23913 11095 23969
rect 11151 23913 11237 23969
rect 11293 23913 11379 23969
rect 11435 23913 11521 23969
rect 11577 23913 11663 23969
rect 11719 23913 11805 23969
rect 11861 23913 11947 23969
rect 12003 23913 12089 23969
rect 12145 23913 12231 23969
rect 12287 23913 12373 23969
rect 12429 23913 12515 23969
rect 12571 23913 12657 23969
rect 12713 23913 12799 23969
rect 12855 23913 12941 23969
rect 12997 23913 13083 23969
rect 13139 23913 13225 23969
rect 13281 23913 13367 23969
rect 13423 23913 13509 23969
rect 13565 23913 13651 23969
rect 13707 23913 13793 23969
rect 13849 23913 13935 23969
rect 13991 23913 14077 23969
rect 14133 23913 14219 23969
rect 14275 23913 14361 23969
rect 14417 23913 14503 23969
rect 14559 23913 14645 23969
rect 14701 23913 14787 23969
rect 14843 23913 14853 23969
rect 151 23827 14853 23913
rect 151 23771 161 23827
rect 217 23771 303 23827
rect 359 23771 445 23827
rect 501 23771 587 23827
rect 643 23771 729 23827
rect 785 23771 871 23827
rect 927 23771 1013 23827
rect 1069 23771 1155 23827
rect 1211 23771 1297 23827
rect 1353 23771 1439 23827
rect 1495 23771 1581 23827
rect 1637 23771 1723 23827
rect 1779 23771 1865 23827
rect 1921 23771 2007 23827
rect 2063 23771 2149 23827
rect 2205 23771 2291 23827
rect 2347 23771 2433 23827
rect 2489 23771 2575 23827
rect 2631 23771 2717 23827
rect 2773 23771 2859 23827
rect 2915 23771 3001 23827
rect 3057 23771 3143 23827
rect 3199 23771 3285 23827
rect 3341 23771 3427 23827
rect 3483 23771 3569 23827
rect 3625 23771 3711 23827
rect 3767 23771 3853 23827
rect 3909 23771 3995 23827
rect 4051 23771 4137 23827
rect 4193 23771 4279 23827
rect 4335 23771 4421 23827
rect 4477 23771 4563 23827
rect 4619 23771 4705 23827
rect 4761 23771 4847 23827
rect 4903 23771 4989 23827
rect 5045 23771 5131 23827
rect 5187 23771 5273 23827
rect 5329 23771 5415 23827
rect 5471 23771 5557 23827
rect 5613 23771 5699 23827
rect 5755 23771 5841 23827
rect 5897 23771 5983 23827
rect 6039 23771 6125 23827
rect 6181 23771 6267 23827
rect 6323 23771 6409 23827
rect 6465 23771 6551 23827
rect 6607 23771 6693 23827
rect 6749 23771 6835 23827
rect 6891 23771 6977 23827
rect 7033 23771 7119 23827
rect 7175 23771 7261 23827
rect 7317 23771 7403 23827
rect 7459 23771 7545 23827
rect 7601 23771 7687 23827
rect 7743 23771 7829 23827
rect 7885 23771 7971 23827
rect 8027 23771 8113 23827
rect 8169 23771 8255 23827
rect 8311 23771 8397 23827
rect 8453 23771 8539 23827
rect 8595 23771 8681 23827
rect 8737 23771 8823 23827
rect 8879 23771 8965 23827
rect 9021 23771 9107 23827
rect 9163 23771 9249 23827
rect 9305 23771 9391 23827
rect 9447 23771 9533 23827
rect 9589 23771 9675 23827
rect 9731 23771 9817 23827
rect 9873 23771 9959 23827
rect 10015 23771 10101 23827
rect 10157 23771 10243 23827
rect 10299 23771 10385 23827
rect 10441 23771 10527 23827
rect 10583 23771 10669 23827
rect 10725 23771 10811 23827
rect 10867 23771 10953 23827
rect 11009 23771 11095 23827
rect 11151 23771 11237 23827
rect 11293 23771 11379 23827
rect 11435 23771 11521 23827
rect 11577 23771 11663 23827
rect 11719 23771 11805 23827
rect 11861 23771 11947 23827
rect 12003 23771 12089 23827
rect 12145 23771 12231 23827
rect 12287 23771 12373 23827
rect 12429 23771 12515 23827
rect 12571 23771 12657 23827
rect 12713 23771 12799 23827
rect 12855 23771 12941 23827
rect 12997 23771 13083 23827
rect 13139 23771 13225 23827
rect 13281 23771 13367 23827
rect 13423 23771 13509 23827
rect 13565 23771 13651 23827
rect 13707 23771 13793 23827
rect 13849 23771 13935 23827
rect 13991 23771 14077 23827
rect 14133 23771 14219 23827
rect 14275 23771 14361 23827
rect 14417 23771 14503 23827
rect 14559 23771 14645 23827
rect 14701 23771 14787 23827
rect 14843 23771 14853 23827
rect 151 23685 14853 23771
rect 151 23629 161 23685
rect 217 23629 303 23685
rect 359 23629 445 23685
rect 501 23629 587 23685
rect 643 23629 729 23685
rect 785 23629 871 23685
rect 927 23629 1013 23685
rect 1069 23629 1155 23685
rect 1211 23629 1297 23685
rect 1353 23629 1439 23685
rect 1495 23629 1581 23685
rect 1637 23629 1723 23685
rect 1779 23629 1865 23685
rect 1921 23629 2007 23685
rect 2063 23629 2149 23685
rect 2205 23629 2291 23685
rect 2347 23629 2433 23685
rect 2489 23629 2575 23685
rect 2631 23629 2717 23685
rect 2773 23629 2859 23685
rect 2915 23629 3001 23685
rect 3057 23629 3143 23685
rect 3199 23629 3285 23685
rect 3341 23629 3427 23685
rect 3483 23629 3569 23685
rect 3625 23629 3711 23685
rect 3767 23629 3853 23685
rect 3909 23629 3995 23685
rect 4051 23629 4137 23685
rect 4193 23629 4279 23685
rect 4335 23629 4421 23685
rect 4477 23629 4563 23685
rect 4619 23629 4705 23685
rect 4761 23629 4847 23685
rect 4903 23629 4989 23685
rect 5045 23629 5131 23685
rect 5187 23629 5273 23685
rect 5329 23629 5415 23685
rect 5471 23629 5557 23685
rect 5613 23629 5699 23685
rect 5755 23629 5841 23685
rect 5897 23629 5983 23685
rect 6039 23629 6125 23685
rect 6181 23629 6267 23685
rect 6323 23629 6409 23685
rect 6465 23629 6551 23685
rect 6607 23629 6693 23685
rect 6749 23629 6835 23685
rect 6891 23629 6977 23685
rect 7033 23629 7119 23685
rect 7175 23629 7261 23685
rect 7317 23629 7403 23685
rect 7459 23629 7545 23685
rect 7601 23629 7687 23685
rect 7743 23629 7829 23685
rect 7885 23629 7971 23685
rect 8027 23629 8113 23685
rect 8169 23629 8255 23685
rect 8311 23629 8397 23685
rect 8453 23629 8539 23685
rect 8595 23629 8681 23685
rect 8737 23629 8823 23685
rect 8879 23629 8965 23685
rect 9021 23629 9107 23685
rect 9163 23629 9249 23685
rect 9305 23629 9391 23685
rect 9447 23629 9533 23685
rect 9589 23629 9675 23685
rect 9731 23629 9817 23685
rect 9873 23629 9959 23685
rect 10015 23629 10101 23685
rect 10157 23629 10243 23685
rect 10299 23629 10385 23685
rect 10441 23629 10527 23685
rect 10583 23629 10669 23685
rect 10725 23629 10811 23685
rect 10867 23629 10953 23685
rect 11009 23629 11095 23685
rect 11151 23629 11237 23685
rect 11293 23629 11379 23685
rect 11435 23629 11521 23685
rect 11577 23629 11663 23685
rect 11719 23629 11805 23685
rect 11861 23629 11947 23685
rect 12003 23629 12089 23685
rect 12145 23629 12231 23685
rect 12287 23629 12373 23685
rect 12429 23629 12515 23685
rect 12571 23629 12657 23685
rect 12713 23629 12799 23685
rect 12855 23629 12941 23685
rect 12997 23629 13083 23685
rect 13139 23629 13225 23685
rect 13281 23629 13367 23685
rect 13423 23629 13509 23685
rect 13565 23629 13651 23685
rect 13707 23629 13793 23685
rect 13849 23629 13935 23685
rect 13991 23629 14077 23685
rect 14133 23629 14219 23685
rect 14275 23629 14361 23685
rect 14417 23629 14503 23685
rect 14559 23629 14645 23685
rect 14701 23629 14787 23685
rect 14843 23629 14853 23685
rect 151 23619 14853 23629
rect 151 23341 14853 23351
rect 151 23285 161 23341
rect 217 23285 303 23341
rect 359 23285 445 23341
rect 501 23285 587 23341
rect 643 23285 729 23341
rect 785 23285 871 23341
rect 927 23285 1013 23341
rect 1069 23285 1155 23341
rect 1211 23285 1297 23341
rect 1353 23285 1439 23341
rect 1495 23285 1581 23341
rect 1637 23285 1723 23341
rect 1779 23285 1865 23341
rect 1921 23285 2007 23341
rect 2063 23285 2149 23341
rect 2205 23285 2291 23341
rect 2347 23285 2433 23341
rect 2489 23285 2575 23341
rect 2631 23285 2717 23341
rect 2773 23285 2859 23341
rect 2915 23285 3001 23341
rect 3057 23285 3143 23341
rect 3199 23285 3285 23341
rect 3341 23285 3427 23341
rect 3483 23285 3569 23341
rect 3625 23285 3711 23341
rect 3767 23285 3853 23341
rect 3909 23285 3995 23341
rect 4051 23285 4137 23341
rect 4193 23285 4279 23341
rect 4335 23285 4421 23341
rect 4477 23285 4563 23341
rect 4619 23285 4705 23341
rect 4761 23285 4847 23341
rect 4903 23285 4989 23341
rect 5045 23285 5131 23341
rect 5187 23285 5273 23341
rect 5329 23285 5415 23341
rect 5471 23285 5557 23341
rect 5613 23285 5699 23341
rect 5755 23285 5841 23341
rect 5897 23285 5983 23341
rect 6039 23285 6125 23341
rect 6181 23285 6267 23341
rect 6323 23285 6409 23341
rect 6465 23285 6551 23341
rect 6607 23285 6693 23341
rect 6749 23285 6835 23341
rect 6891 23285 6977 23341
rect 7033 23285 7119 23341
rect 7175 23285 7261 23341
rect 7317 23285 7403 23341
rect 7459 23285 7545 23341
rect 7601 23285 7687 23341
rect 7743 23285 7829 23341
rect 7885 23285 7971 23341
rect 8027 23285 8113 23341
rect 8169 23285 8255 23341
rect 8311 23285 8397 23341
rect 8453 23285 8539 23341
rect 8595 23285 8681 23341
rect 8737 23285 8823 23341
rect 8879 23285 8965 23341
rect 9021 23285 9107 23341
rect 9163 23285 9249 23341
rect 9305 23285 9391 23341
rect 9447 23285 9533 23341
rect 9589 23285 9675 23341
rect 9731 23285 9817 23341
rect 9873 23285 9959 23341
rect 10015 23285 10101 23341
rect 10157 23285 10243 23341
rect 10299 23285 10385 23341
rect 10441 23285 10527 23341
rect 10583 23285 10669 23341
rect 10725 23285 10811 23341
rect 10867 23285 10953 23341
rect 11009 23285 11095 23341
rect 11151 23285 11237 23341
rect 11293 23285 11379 23341
rect 11435 23285 11521 23341
rect 11577 23285 11663 23341
rect 11719 23285 11805 23341
rect 11861 23285 11947 23341
rect 12003 23285 12089 23341
rect 12145 23285 12231 23341
rect 12287 23285 12373 23341
rect 12429 23285 12515 23341
rect 12571 23285 12657 23341
rect 12713 23285 12799 23341
rect 12855 23285 12941 23341
rect 12997 23285 13083 23341
rect 13139 23285 13225 23341
rect 13281 23285 13367 23341
rect 13423 23285 13509 23341
rect 13565 23285 13651 23341
rect 13707 23285 13793 23341
rect 13849 23285 13935 23341
rect 13991 23285 14077 23341
rect 14133 23285 14219 23341
rect 14275 23285 14361 23341
rect 14417 23285 14503 23341
rect 14559 23285 14645 23341
rect 14701 23285 14787 23341
rect 14843 23285 14853 23341
rect 151 23199 14853 23285
rect 151 23143 161 23199
rect 217 23143 303 23199
rect 359 23143 445 23199
rect 501 23143 587 23199
rect 643 23143 729 23199
rect 785 23143 871 23199
rect 927 23143 1013 23199
rect 1069 23143 1155 23199
rect 1211 23143 1297 23199
rect 1353 23143 1439 23199
rect 1495 23143 1581 23199
rect 1637 23143 1723 23199
rect 1779 23143 1865 23199
rect 1921 23143 2007 23199
rect 2063 23143 2149 23199
rect 2205 23143 2291 23199
rect 2347 23143 2433 23199
rect 2489 23143 2575 23199
rect 2631 23143 2717 23199
rect 2773 23143 2859 23199
rect 2915 23143 3001 23199
rect 3057 23143 3143 23199
rect 3199 23143 3285 23199
rect 3341 23143 3427 23199
rect 3483 23143 3569 23199
rect 3625 23143 3711 23199
rect 3767 23143 3853 23199
rect 3909 23143 3995 23199
rect 4051 23143 4137 23199
rect 4193 23143 4279 23199
rect 4335 23143 4421 23199
rect 4477 23143 4563 23199
rect 4619 23143 4705 23199
rect 4761 23143 4847 23199
rect 4903 23143 4989 23199
rect 5045 23143 5131 23199
rect 5187 23143 5273 23199
rect 5329 23143 5415 23199
rect 5471 23143 5557 23199
rect 5613 23143 5699 23199
rect 5755 23143 5841 23199
rect 5897 23143 5983 23199
rect 6039 23143 6125 23199
rect 6181 23143 6267 23199
rect 6323 23143 6409 23199
rect 6465 23143 6551 23199
rect 6607 23143 6693 23199
rect 6749 23143 6835 23199
rect 6891 23143 6977 23199
rect 7033 23143 7119 23199
rect 7175 23143 7261 23199
rect 7317 23143 7403 23199
rect 7459 23143 7545 23199
rect 7601 23143 7687 23199
rect 7743 23143 7829 23199
rect 7885 23143 7971 23199
rect 8027 23143 8113 23199
rect 8169 23143 8255 23199
rect 8311 23143 8397 23199
rect 8453 23143 8539 23199
rect 8595 23143 8681 23199
rect 8737 23143 8823 23199
rect 8879 23143 8965 23199
rect 9021 23143 9107 23199
rect 9163 23143 9249 23199
rect 9305 23143 9391 23199
rect 9447 23143 9533 23199
rect 9589 23143 9675 23199
rect 9731 23143 9817 23199
rect 9873 23143 9959 23199
rect 10015 23143 10101 23199
rect 10157 23143 10243 23199
rect 10299 23143 10385 23199
rect 10441 23143 10527 23199
rect 10583 23143 10669 23199
rect 10725 23143 10811 23199
rect 10867 23143 10953 23199
rect 11009 23143 11095 23199
rect 11151 23143 11237 23199
rect 11293 23143 11379 23199
rect 11435 23143 11521 23199
rect 11577 23143 11663 23199
rect 11719 23143 11805 23199
rect 11861 23143 11947 23199
rect 12003 23143 12089 23199
rect 12145 23143 12231 23199
rect 12287 23143 12373 23199
rect 12429 23143 12515 23199
rect 12571 23143 12657 23199
rect 12713 23143 12799 23199
rect 12855 23143 12941 23199
rect 12997 23143 13083 23199
rect 13139 23143 13225 23199
rect 13281 23143 13367 23199
rect 13423 23143 13509 23199
rect 13565 23143 13651 23199
rect 13707 23143 13793 23199
rect 13849 23143 13935 23199
rect 13991 23143 14077 23199
rect 14133 23143 14219 23199
rect 14275 23143 14361 23199
rect 14417 23143 14503 23199
rect 14559 23143 14645 23199
rect 14701 23143 14787 23199
rect 14843 23143 14853 23199
rect 151 23057 14853 23143
rect 151 23001 161 23057
rect 217 23001 303 23057
rect 359 23001 445 23057
rect 501 23001 587 23057
rect 643 23001 729 23057
rect 785 23001 871 23057
rect 927 23001 1013 23057
rect 1069 23001 1155 23057
rect 1211 23001 1297 23057
rect 1353 23001 1439 23057
rect 1495 23001 1581 23057
rect 1637 23001 1723 23057
rect 1779 23001 1865 23057
rect 1921 23001 2007 23057
rect 2063 23001 2149 23057
rect 2205 23001 2291 23057
rect 2347 23001 2433 23057
rect 2489 23001 2575 23057
rect 2631 23001 2717 23057
rect 2773 23001 2859 23057
rect 2915 23001 3001 23057
rect 3057 23001 3143 23057
rect 3199 23001 3285 23057
rect 3341 23001 3427 23057
rect 3483 23001 3569 23057
rect 3625 23001 3711 23057
rect 3767 23001 3853 23057
rect 3909 23001 3995 23057
rect 4051 23001 4137 23057
rect 4193 23001 4279 23057
rect 4335 23001 4421 23057
rect 4477 23001 4563 23057
rect 4619 23001 4705 23057
rect 4761 23001 4847 23057
rect 4903 23001 4989 23057
rect 5045 23001 5131 23057
rect 5187 23001 5273 23057
rect 5329 23001 5415 23057
rect 5471 23001 5557 23057
rect 5613 23001 5699 23057
rect 5755 23001 5841 23057
rect 5897 23001 5983 23057
rect 6039 23001 6125 23057
rect 6181 23001 6267 23057
rect 6323 23001 6409 23057
rect 6465 23001 6551 23057
rect 6607 23001 6693 23057
rect 6749 23001 6835 23057
rect 6891 23001 6977 23057
rect 7033 23001 7119 23057
rect 7175 23001 7261 23057
rect 7317 23001 7403 23057
rect 7459 23001 7545 23057
rect 7601 23001 7687 23057
rect 7743 23001 7829 23057
rect 7885 23001 7971 23057
rect 8027 23001 8113 23057
rect 8169 23001 8255 23057
rect 8311 23001 8397 23057
rect 8453 23001 8539 23057
rect 8595 23001 8681 23057
rect 8737 23001 8823 23057
rect 8879 23001 8965 23057
rect 9021 23001 9107 23057
rect 9163 23001 9249 23057
rect 9305 23001 9391 23057
rect 9447 23001 9533 23057
rect 9589 23001 9675 23057
rect 9731 23001 9817 23057
rect 9873 23001 9959 23057
rect 10015 23001 10101 23057
rect 10157 23001 10243 23057
rect 10299 23001 10385 23057
rect 10441 23001 10527 23057
rect 10583 23001 10669 23057
rect 10725 23001 10811 23057
rect 10867 23001 10953 23057
rect 11009 23001 11095 23057
rect 11151 23001 11237 23057
rect 11293 23001 11379 23057
rect 11435 23001 11521 23057
rect 11577 23001 11663 23057
rect 11719 23001 11805 23057
rect 11861 23001 11947 23057
rect 12003 23001 12089 23057
rect 12145 23001 12231 23057
rect 12287 23001 12373 23057
rect 12429 23001 12515 23057
rect 12571 23001 12657 23057
rect 12713 23001 12799 23057
rect 12855 23001 12941 23057
rect 12997 23001 13083 23057
rect 13139 23001 13225 23057
rect 13281 23001 13367 23057
rect 13423 23001 13509 23057
rect 13565 23001 13651 23057
rect 13707 23001 13793 23057
rect 13849 23001 13935 23057
rect 13991 23001 14077 23057
rect 14133 23001 14219 23057
rect 14275 23001 14361 23057
rect 14417 23001 14503 23057
rect 14559 23001 14645 23057
rect 14701 23001 14787 23057
rect 14843 23001 14853 23057
rect 151 22915 14853 23001
rect 151 22859 161 22915
rect 217 22859 303 22915
rect 359 22859 445 22915
rect 501 22859 587 22915
rect 643 22859 729 22915
rect 785 22859 871 22915
rect 927 22859 1013 22915
rect 1069 22859 1155 22915
rect 1211 22859 1297 22915
rect 1353 22859 1439 22915
rect 1495 22859 1581 22915
rect 1637 22859 1723 22915
rect 1779 22859 1865 22915
rect 1921 22859 2007 22915
rect 2063 22859 2149 22915
rect 2205 22859 2291 22915
rect 2347 22859 2433 22915
rect 2489 22859 2575 22915
rect 2631 22859 2717 22915
rect 2773 22859 2859 22915
rect 2915 22859 3001 22915
rect 3057 22859 3143 22915
rect 3199 22859 3285 22915
rect 3341 22859 3427 22915
rect 3483 22859 3569 22915
rect 3625 22859 3711 22915
rect 3767 22859 3853 22915
rect 3909 22859 3995 22915
rect 4051 22859 4137 22915
rect 4193 22859 4279 22915
rect 4335 22859 4421 22915
rect 4477 22859 4563 22915
rect 4619 22859 4705 22915
rect 4761 22859 4847 22915
rect 4903 22859 4989 22915
rect 5045 22859 5131 22915
rect 5187 22859 5273 22915
rect 5329 22859 5415 22915
rect 5471 22859 5557 22915
rect 5613 22859 5699 22915
rect 5755 22859 5841 22915
rect 5897 22859 5983 22915
rect 6039 22859 6125 22915
rect 6181 22859 6267 22915
rect 6323 22859 6409 22915
rect 6465 22859 6551 22915
rect 6607 22859 6693 22915
rect 6749 22859 6835 22915
rect 6891 22859 6977 22915
rect 7033 22859 7119 22915
rect 7175 22859 7261 22915
rect 7317 22859 7403 22915
rect 7459 22859 7545 22915
rect 7601 22859 7687 22915
rect 7743 22859 7829 22915
rect 7885 22859 7971 22915
rect 8027 22859 8113 22915
rect 8169 22859 8255 22915
rect 8311 22859 8397 22915
rect 8453 22859 8539 22915
rect 8595 22859 8681 22915
rect 8737 22859 8823 22915
rect 8879 22859 8965 22915
rect 9021 22859 9107 22915
rect 9163 22859 9249 22915
rect 9305 22859 9391 22915
rect 9447 22859 9533 22915
rect 9589 22859 9675 22915
rect 9731 22859 9817 22915
rect 9873 22859 9959 22915
rect 10015 22859 10101 22915
rect 10157 22859 10243 22915
rect 10299 22859 10385 22915
rect 10441 22859 10527 22915
rect 10583 22859 10669 22915
rect 10725 22859 10811 22915
rect 10867 22859 10953 22915
rect 11009 22859 11095 22915
rect 11151 22859 11237 22915
rect 11293 22859 11379 22915
rect 11435 22859 11521 22915
rect 11577 22859 11663 22915
rect 11719 22859 11805 22915
rect 11861 22859 11947 22915
rect 12003 22859 12089 22915
rect 12145 22859 12231 22915
rect 12287 22859 12373 22915
rect 12429 22859 12515 22915
rect 12571 22859 12657 22915
rect 12713 22859 12799 22915
rect 12855 22859 12941 22915
rect 12997 22859 13083 22915
rect 13139 22859 13225 22915
rect 13281 22859 13367 22915
rect 13423 22859 13509 22915
rect 13565 22859 13651 22915
rect 13707 22859 13793 22915
rect 13849 22859 13935 22915
rect 13991 22859 14077 22915
rect 14133 22859 14219 22915
rect 14275 22859 14361 22915
rect 14417 22859 14503 22915
rect 14559 22859 14645 22915
rect 14701 22859 14787 22915
rect 14843 22859 14853 22915
rect 151 22773 14853 22859
rect 151 22717 161 22773
rect 217 22717 303 22773
rect 359 22717 445 22773
rect 501 22717 587 22773
rect 643 22717 729 22773
rect 785 22717 871 22773
rect 927 22717 1013 22773
rect 1069 22717 1155 22773
rect 1211 22717 1297 22773
rect 1353 22717 1439 22773
rect 1495 22717 1581 22773
rect 1637 22717 1723 22773
rect 1779 22717 1865 22773
rect 1921 22717 2007 22773
rect 2063 22717 2149 22773
rect 2205 22717 2291 22773
rect 2347 22717 2433 22773
rect 2489 22717 2575 22773
rect 2631 22717 2717 22773
rect 2773 22717 2859 22773
rect 2915 22717 3001 22773
rect 3057 22717 3143 22773
rect 3199 22717 3285 22773
rect 3341 22717 3427 22773
rect 3483 22717 3569 22773
rect 3625 22717 3711 22773
rect 3767 22717 3853 22773
rect 3909 22717 3995 22773
rect 4051 22717 4137 22773
rect 4193 22717 4279 22773
rect 4335 22717 4421 22773
rect 4477 22717 4563 22773
rect 4619 22717 4705 22773
rect 4761 22717 4847 22773
rect 4903 22717 4989 22773
rect 5045 22717 5131 22773
rect 5187 22717 5273 22773
rect 5329 22717 5415 22773
rect 5471 22717 5557 22773
rect 5613 22717 5699 22773
rect 5755 22717 5841 22773
rect 5897 22717 5983 22773
rect 6039 22717 6125 22773
rect 6181 22717 6267 22773
rect 6323 22717 6409 22773
rect 6465 22717 6551 22773
rect 6607 22717 6693 22773
rect 6749 22717 6835 22773
rect 6891 22717 6977 22773
rect 7033 22717 7119 22773
rect 7175 22717 7261 22773
rect 7317 22717 7403 22773
rect 7459 22717 7545 22773
rect 7601 22717 7687 22773
rect 7743 22717 7829 22773
rect 7885 22717 7971 22773
rect 8027 22717 8113 22773
rect 8169 22717 8255 22773
rect 8311 22717 8397 22773
rect 8453 22717 8539 22773
rect 8595 22717 8681 22773
rect 8737 22717 8823 22773
rect 8879 22717 8965 22773
rect 9021 22717 9107 22773
rect 9163 22717 9249 22773
rect 9305 22717 9391 22773
rect 9447 22717 9533 22773
rect 9589 22717 9675 22773
rect 9731 22717 9817 22773
rect 9873 22717 9959 22773
rect 10015 22717 10101 22773
rect 10157 22717 10243 22773
rect 10299 22717 10385 22773
rect 10441 22717 10527 22773
rect 10583 22717 10669 22773
rect 10725 22717 10811 22773
rect 10867 22717 10953 22773
rect 11009 22717 11095 22773
rect 11151 22717 11237 22773
rect 11293 22717 11379 22773
rect 11435 22717 11521 22773
rect 11577 22717 11663 22773
rect 11719 22717 11805 22773
rect 11861 22717 11947 22773
rect 12003 22717 12089 22773
rect 12145 22717 12231 22773
rect 12287 22717 12373 22773
rect 12429 22717 12515 22773
rect 12571 22717 12657 22773
rect 12713 22717 12799 22773
rect 12855 22717 12941 22773
rect 12997 22717 13083 22773
rect 13139 22717 13225 22773
rect 13281 22717 13367 22773
rect 13423 22717 13509 22773
rect 13565 22717 13651 22773
rect 13707 22717 13793 22773
rect 13849 22717 13935 22773
rect 13991 22717 14077 22773
rect 14133 22717 14219 22773
rect 14275 22717 14361 22773
rect 14417 22717 14503 22773
rect 14559 22717 14645 22773
rect 14701 22717 14787 22773
rect 14843 22717 14853 22773
rect 151 22631 14853 22717
rect 151 22575 161 22631
rect 217 22575 303 22631
rect 359 22575 445 22631
rect 501 22575 587 22631
rect 643 22575 729 22631
rect 785 22575 871 22631
rect 927 22575 1013 22631
rect 1069 22575 1155 22631
rect 1211 22575 1297 22631
rect 1353 22575 1439 22631
rect 1495 22575 1581 22631
rect 1637 22575 1723 22631
rect 1779 22575 1865 22631
rect 1921 22575 2007 22631
rect 2063 22575 2149 22631
rect 2205 22575 2291 22631
rect 2347 22575 2433 22631
rect 2489 22575 2575 22631
rect 2631 22575 2717 22631
rect 2773 22575 2859 22631
rect 2915 22575 3001 22631
rect 3057 22575 3143 22631
rect 3199 22575 3285 22631
rect 3341 22575 3427 22631
rect 3483 22575 3569 22631
rect 3625 22575 3711 22631
rect 3767 22575 3853 22631
rect 3909 22575 3995 22631
rect 4051 22575 4137 22631
rect 4193 22575 4279 22631
rect 4335 22575 4421 22631
rect 4477 22575 4563 22631
rect 4619 22575 4705 22631
rect 4761 22575 4847 22631
rect 4903 22575 4989 22631
rect 5045 22575 5131 22631
rect 5187 22575 5273 22631
rect 5329 22575 5415 22631
rect 5471 22575 5557 22631
rect 5613 22575 5699 22631
rect 5755 22575 5841 22631
rect 5897 22575 5983 22631
rect 6039 22575 6125 22631
rect 6181 22575 6267 22631
rect 6323 22575 6409 22631
rect 6465 22575 6551 22631
rect 6607 22575 6693 22631
rect 6749 22575 6835 22631
rect 6891 22575 6977 22631
rect 7033 22575 7119 22631
rect 7175 22575 7261 22631
rect 7317 22575 7403 22631
rect 7459 22575 7545 22631
rect 7601 22575 7687 22631
rect 7743 22575 7829 22631
rect 7885 22575 7971 22631
rect 8027 22575 8113 22631
rect 8169 22575 8255 22631
rect 8311 22575 8397 22631
rect 8453 22575 8539 22631
rect 8595 22575 8681 22631
rect 8737 22575 8823 22631
rect 8879 22575 8965 22631
rect 9021 22575 9107 22631
rect 9163 22575 9249 22631
rect 9305 22575 9391 22631
rect 9447 22575 9533 22631
rect 9589 22575 9675 22631
rect 9731 22575 9817 22631
rect 9873 22575 9959 22631
rect 10015 22575 10101 22631
rect 10157 22575 10243 22631
rect 10299 22575 10385 22631
rect 10441 22575 10527 22631
rect 10583 22575 10669 22631
rect 10725 22575 10811 22631
rect 10867 22575 10953 22631
rect 11009 22575 11095 22631
rect 11151 22575 11237 22631
rect 11293 22575 11379 22631
rect 11435 22575 11521 22631
rect 11577 22575 11663 22631
rect 11719 22575 11805 22631
rect 11861 22575 11947 22631
rect 12003 22575 12089 22631
rect 12145 22575 12231 22631
rect 12287 22575 12373 22631
rect 12429 22575 12515 22631
rect 12571 22575 12657 22631
rect 12713 22575 12799 22631
rect 12855 22575 12941 22631
rect 12997 22575 13083 22631
rect 13139 22575 13225 22631
rect 13281 22575 13367 22631
rect 13423 22575 13509 22631
rect 13565 22575 13651 22631
rect 13707 22575 13793 22631
rect 13849 22575 13935 22631
rect 13991 22575 14077 22631
rect 14133 22575 14219 22631
rect 14275 22575 14361 22631
rect 14417 22575 14503 22631
rect 14559 22575 14645 22631
rect 14701 22575 14787 22631
rect 14843 22575 14853 22631
rect 151 22489 14853 22575
rect 151 22433 161 22489
rect 217 22433 303 22489
rect 359 22433 445 22489
rect 501 22433 587 22489
rect 643 22433 729 22489
rect 785 22433 871 22489
rect 927 22433 1013 22489
rect 1069 22433 1155 22489
rect 1211 22433 1297 22489
rect 1353 22433 1439 22489
rect 1495 22433 1581 22489
rect 1637 22433 1723 22489
rect 1779 22433 1865 22489
rect 1921 22433 2007 22489
rect 2063 22433 2149 22489
rect 2205 22433 2291 22489
rect 2347 22433 2433 22489
rect 2489 22433 2575 22489
rect 2631 22433 2717 22489
rect 2773 22433 2859 22489
rect 2915 22433 3001 22489
rect 3057 22433 3143 22489
rect 3199 22433 3285 22489
rect 3341 22433 3427 22489
rect 3483 22433 3569 22489
rect 3625 22433 3711 22489
rect 3767 22433 3853 22489
rect 3909 22433 3995 22489
rect 4051 22433 4137 22489
rect 4193 22433 4279 22489
rect 4335 22433 4421 22489
rect 4477 22433 4563 22489
rect 4619 22433 4705 22489
rect 4761 22433 4847 22489
rect 4903 22433 4989 22489
rect 5045 22433 5131 22489
rect 5187 22433 5273 22489
rect 5329 22433 5415 22489
rect 5471 22433 5557 22489
rect 5613 22433 5699 22489
rect 5755 22433 5841 22489
rect 5897 22433 5983 22489
rect 6039 22433 6125 22489
rect 6181 22433 6267 22489
rect 6323 22433 6409 22489
rect 6465 22433 6551 22489
rect 6607 22433 6693 22489
rect 6749 22433 6835 22489
rect 6891 22433 6977 22489
rect 7033 22433 7119 22489
rect 7175 22433 7261 22489
rect 7317 22433 7403 22489
rect 7459 22433 7545 22489
rect 7601 22433 7687 22489
rect 7743 22433 7829 22489
rect 7885 22433 7971 22489
rect 8027 22433 8113 22489
rect 8169 22433 8255 22489
rect 8311 22433 8397 22489
rect 8453 22433 8539 22489
rect 8595 22433 8681 22489
rect 8737 22433 8823 22489
rect 8879 22433 8965 22489
rect 9021 22433 9107 22489
rect 9163 22433 9249 22489
rect 9305 22433 9391 22489
rect 9447 22433 9533 22489
rect 9589 22433 9675 22489
rect 9731 22433 9817 22489
rect 9873 22433 9959 22489
rect 10015 22433 10101 22489
rect 10157 22433 10243 22489
rect 10299 22433 10385 22489
rect 10441 22433 10527 22489
rect 10583 22433 10669 22489
rect 10725 22433 10811 22489
rect 10867 22433 10953 22489
rect 11009 22433 11095 22489
rect 11151 22433 11237 22489
rect 11293 22433 11379 22489
rect 11435 22433 11521 22489
rect 11577 22433 11663 22489
rect 11719 22433 11805 22489
rect 11861 22433 11947 22489
rect 12003 22433 12089 22489
rect 12145 22433 12231 22489
rect 12287 22433 12373 22489
rect 12429 22433 12515 22489
rect 12571 22433 12657 22489
rect 12713 22433 12799 22489
rect 12855 22433 12941 22489
rect 12997 22433 13083 22489
rect 13139 22433 13225 22489
rect 13281 22433 13367 22489
rect 13423 22433 13509 22489
rect 13565 22433 13651 22489
rect 13707 22433 13793 22489
rect 13849 22433 13935 22489
rect 13991 22433 14077 22489
rect 14133 22433 14219 22489
rect 14275 22433 14361 22489
rect 14417 22433 14503 22489
rect 14559 22433 14645 22489
rect 14701 22433 14787 22489
rect 14843 22433 14853 22489
rect 151 22347 14853 22433
rect 151 22291 161 22347
rect 217 22291 303 22347
rect 359 22291 445 22347
rect 501 22291 587 22347
rect 643 22291 729 22347
rect 785 22291 871 22347
rect 927 22291 1013 22347
rect 1069 22291 1155 22347
rect 1211 22291 1297 22347
rect 1353 22291 1439 22347
rect 1495 22291 1581 22347
rect 1637 22291 1723 22347
rect 1779 22291 1865 22347
rect 1921 22291 2007 22347
rect 2063 22291 2149 22347
rect 2205 22291 2291 22347
rect 2347 22291 2433 22347
rect 2489 22291 2575 22347
rect 2631 22291 2717 22347
rect 2773 22291 2859 22347
rect 2915 22291 3001 22347
rect 3057 22291 3143 22347
rect 3199 22291 3285 22347
rect 3341 22291 3427 22347
rect 3483 22291 3569 22347
rect 3625 22291 3711 22347
rect 3767 22291 3853 22347
rect 3909 22291 3995 22347
rect 4051 22291 4137 22347
rect 4193 22291 4279 22347
rect 4335 22291 4421 22347
rect 4477 22291 4563 22347
rect 4619 22291 4705 22347
rect 4761 22291 4847 22347
rect 4903 22291 4989 22347
rect 5045 22291 5131 22347
rect 5187 22291 5273 22347
rect 5329 22291 5415 22347
rect 5471 22291 5557 22347
rect 5613 22291 5699 22347
rect 5755 22291 5841 22347
rect 5897 22291 5983 22347
rect 6039 22291 6125 22347
rect 6181 22291 6267 22347
rect 6323 22291 6409 22347
rect 6465 22291 6551 22347
rect 6607 22291 6693 22347
rect 6749 22291 6835 22347
rect 6891 22291 6977 22347
rect 7033 22291 7119 22347
rect 7175 22291 7261 22347
rect 7317 22291 7403 22347
rect 7459 22291 7545 22347
rect 7601 22291 7687 22347
rect 7743 22291 7829 22347
rect 7885 22291 7971 22347
rect 8027 22291 8113 22347
rect 8169 22291 8255 22347
rect 8311 22291 8397 22347
rect 8453 22291 8539 22347
rect 8595 22291 8681 22347
rect 8737 22291 8823 22347
rect 8879 22291 8965 22347
rect 9021 22291 9107 22347
rect 9163 22291 9249 22347
rect 9305 22291 9391 22347
rect 9447 22291 9533 22347
rect 9589 22291 9675 22347
rect 9731 22291 9817 22347
rect 9873 22291 9959 22347
rect 10015 22291 10101 22347
rect 10157 22291 10243 22347
rect 10299 22291 10385 22347
rect 10441 22291 10527 22347
rect 10583 22291 10669 22347
rect 10725 22291 10811 22347
rect 10867 22291 10953 22347
rect 11009 22291 11095 22347
rect 11151 22291 11237 22347
rect 11293 22291 11379 22347
rect 11435 22291 11521 22347
rect 11577 22291 11663 22347
rect 11719 22291 11805 22347
rect 11861 22291 11947 22347
rect 12003 22291 12089 22347
rect 12145 22291 12231 22347
rect 12287 22291 12373 22347
rect 12429 22291 12515 22347
rect 12571 22291 12657 22347
rect 12713 22291 12799 22347
rect 12855 22291 12941 22347
rect 12997 22291 13083 22347
rect 13139 22291 13225 22347
rect 13281 22291 13367 22347
rect 13423 22291 13509 22347
rect 13565 22291 13651 22347
rect 13707 22291 13793 22347
rect 13849 22291 13935 22347
rect 13991 22291 14077 22347
rect 14133 22291 14219 22347
rect 14275 22291 14361 22347
rect 14417 22291 14503 22347
rect 14559 22291 14645 22347
rect 14701 22291 14787 22347
rect 14843 22291 14853 22347
rect 151 22205 14853 22291
rect 151 22149 161 22205
rect 217 22149 303 22205
rect 359 22149 445 22205
rect 501 22149 587 22205
rect 643 22149 729 22205
rect 785 22149 871 22205
rect 927 22149 1013 22205
rect 1069 22149 1155 22205
rect 1211 22149 1297 22205
rect 1353 22149 1439 22205
rect 1495 22149 1581 22205
rect 1637 22149 1723 22205
rect 1779 22149 1865 22205
rect 1921 22149 2007 22205
rect 2063 22149 2149 22205
rect 2205 22149 2291 22205
rect 2347 22149 2433 22205
rect 2489 22149 2575 22205
rect 2631 22149 2717 22205
rect 2773 22149 2859 22205
rect 2915 22149 3001 22205
rect 3057 22149 3143 22205
rect 3199 22149 3285 22205
rect 3341 22149 3427 22205
rect 3483 22149 3569 22205
rect 3625 22149 3711 22205
rect 3767 22149 3853 22205
rect 3909 22149 3995 22205
rect 4051 22149 4137 22205
rect 4193 22149 4279 22205
rect 4335 22149 4421 22205
rect 4477 22149 4563 22205
rect 4619 22149 4705 22205
rect 4761 22149 4847 22205
rect 4903 22149 4989 22205
rect 5045 22149 5131 22205
rect 5187 22149 5273 22205
rect 5329 22149 5415 22205
rect 5471 22149 5557 22205
rect 5613 22149 5699 22205
rect 5755 22149 5841 22205
rect 5897 22149 5983 22205
rect 6039 22149 6125 22205
rect 6181 22149 6267 22205
rect 6323 22149 6409 22205
rect 6465 22149 6551 22205
rect 6607 22149 6693 22205
rect 6749 22149 6835 22205
rect 6891 22149 6977 22205
rect 7033 22149 7119 22205
rect 7175 22149 7261 22205
rect 7317 22149 7403 22205
rect 7459 22149 7545 22205
rect 7601 22149 7687 22205
rect 7743 22149 7829 22205
rect 7885 22149 7971 22205
rect 8027 22149 8113 22205
rect 8169 22149 8255 22205
rect 8311 22149 8397 22205
rect 8453 22149 8539 22205
rect 8595 22149 8681 22205
rect 8737 22149 8823 22205
rect 8879 22149 8965 22205
rect 9021 22149 9107 22205
rect 9163 22149 9249 22205
rect 9305 22149 9391 22205
rect 9447 22149 9533 22205
rect 9589 22149 9675 22205
rect 9731 22149 9817 22205
rect 9873 22149 9959 22205
rect 10015 22149 10101 22205
rect 10157 22149 10243 22205
rect 10299 22149 10385 22205
rect 10441 22149 10527 22205
rect 10583 22149 10669 22205
rect 10725 22149 10811 22205
rect 10867 22149 10953 22205
rect 11009 22149 11095 22205
rect 11151 22149 11237 22205
rect 11293 22149 11379 22205
rect 11435 22149 11521 22205
rect 11577 22149 11663 22205
rect 11719 22149 11805 22205
rect 11861 22149 11947 22205
rect 12003 22149 12089 22205
rect 12145 22149 12231 22205
rect 12287 22149 12373 22205
rect 12429 22149 12515 22205
rect 12571 22149 12657 22205
rect 12713 22149 12799 22205
rect 12855 22149 12941 22205
rect 12997 22149 13083 22205
rect 13139 22149 13225 22205
rect 13281 22149 13367 22205
rect 13423 22149 13509 22205
rect 13565 22149 13651 22205
rect 13707 22149 13793 22205
rect 13849 22149 13935 22205
rect 13991 22149 14077 22205
rect 14133 22149 14219 22205
rect 14275 22149 14361 22205
rect 14417 22149 14503 22205
rect 14559 22149 14645 22205
rect 14701 22149 14787 22205
rect 14843 22149 14853 22205
rect 151 22063 14853 22149
rect 151 22007 161 22063
rect 217 22007 303 22063
rect 359 22007 445 22063
rect 501 22007 587 22063
rect 643 22007 729 22063
rect 785 22007 871 22063
rect 927 22007 1013 22063
rect 1069 22007 1155 22063
rect 1211 22007 1297 22063
rect 1353 22007 1439 22063
rect 1495 22007 1581 22063
rect 1637 22007 1723 22063
rect 1779 22007 1865 22063
rect 1921 22007 2007 22063
rect 2063 22007 2149 22063
rect 2205 22007 2291 22063
rect 2347 22007 2433 22063
rect 2489 22007 2575 22063
rect 2631 22007 2717 22063
rect 2773 22007 2859 22063
rect 2915 22007 3001 22063
rect 3057 22007 3143 22063
rect 3199 22007 3285 22063
rect 3341 22007 3427 22063
rect 3483 22007 3569 22063
rect 3625 22007 3711 22063
rect 3767 22007 3853 22063
rect 3909 22007 3995 22063
rect 4051 22007 4137 22063
rect 4193 22007 4279 22063
rect 4335 22007 4421 22063
rect 4477 22007 4563 22063
rect 4619 22007 4705 22063
rect 4761 22007 4847 22063
rect 4903 22007 4989 22063
rect 5045 22007 5131 22063
rect 5187 22007 5273 22063
rect 5329 22007 5415 22063
rect 5471 22007 5557 22063
rect 5613 22007 5699 22063
rect 5755 22007 5841 22063
rect 5897 22007 5983 22063
rect 6039 22007 6125 22063
rect 6181 22007 6267 22063
rect 6323 22007 6409 22063
rect 6465 22007 6551 22063
rect 6607 22007 6693 22063
rect 6749 22007 6835 22063
rect 6891 22007 6977 22063
rect 7033 22007 7119 22063
rect 7175 22007 7261 22063
rect 7317 22007 7403 22063
rect 7459 22007 7545 22063
rect 7601 22007 7687 22063
rect 7743 22007 7829 22063
rect 7885 22007 7971 22063
rect 8027 22007 8113 22063
rect 8169 22007 8255 22063
rect 8311 22007 8397 22063
rect 8453 22007 8539 22063
rect 8595 22007 8681 22063
rect 8737 22007 8823 22063
rect 8879 22007 8965 22063
rect 9021 22007 9107 22063
rect 9163 22007 9249 22063
rect 9305 22007 9391 22063
rect 9447 22007 9533 22063
rect 9589 22007 9675 22063
rect 9731 22007 9817 22063
rect 9873 22007 9959 22063
rect 10015 22007 10101 22063
rect 10157 22007 10243 22063
rect 10299 22007 10385 22063
rect 10441 22007 10527 22063
rect 10583 22007 10669 22063
rect 10725 22007 10811 22063
rect 10867 22007 10953 22063
rect 11009 22007 11095 22063
rect 11151 22007 11237 22063
rect 11293 22007 11379 22063
rect 11435 22007 11521 22063
rect 11577 22007 11663 22063
rect 11719 22007 11805 22063
rect 11861 22007 11947 22063
rect 12003 22007 12089 22063
rect 12145 22007 12231 22063
rect 12287 22007 12373 22063
rect 12429 22007 12515 22063
rect 12571 22007 12657 22063
rect 12713 22007 12799 22063
rect 12855 22007 12941 22063
rect 12997 22007 13083 22063
rect 13139 22007 13225 22063
rect 13281 22007 13367 22063
rect 13423 22007 13509 22063
rect 13565 22007 13651 22063
rect 13707 22007 13793 22063
rect 13849 22007 13935 22063
rect 13991 22007 14077 22063
rect 14133 22007 14219 22063
rect 14275 22007 14361 22063
rect 14417 22007 14503 22063
rect 14559 22007 14645 22063
rect 14701 22007 14787 22063
rect 14843 22007 14853 22063
rect 151 21921 14853 22007
rect 151 21865 161 21921
rect 217 21865 303 21921
rect 359 21865 445 21921
rect 501 21865 587 21921
rect 643 21865 729 21921
rect 785 21865 871 21921
rect 927 21865 1013 21921
rect 1069 21865 1155 21921
rect 1211 21865 1297 21921
rect 1353 21865 1439 21921
rect 1495 21865 1581 21921
rect 1637 21865 1723 21921
rect 1779 21865 1865 21921
rect 1921 21865 2007 21921
rect 2063 21865 2149 21921
rect 2205 21865 2291 21921
rect 2347 21865 2433 21921
rect 2489 21865 2575 21921
rect 2631 21865 2717 21921
rect 2773 21865 2859 21921
rect 2915 21865 3001 21921
rect 3057 21865 3143 21921
rect 3199 21865 3285 21921
rect 3341 21865 3427 21921
rect 3483 21865 3569 21921
rect 3625 21865 3711 21921
rect 3767 21865 3853 21921
rect 3909 21865 3995 21921
rect 4051 21865 4137 21921
rect 4193 21865 4279 21921
rect 4335 21865 4421 21921
rect 4477 21865 4563 21921
rect 4619 21865 4705 21921
rect 4761 21865 4847 21921
rect 4903 21865 4989 21921
rect 5045 21865 5131 21921
rect 5187 21865 5273 21921
rect 5329 21865 5415 21921
rect 5471 21865 5557 21921
rect 5613 21865 5699 21921
rect 5755 21865 5841 21921
rect 5897 21865 5983 21921
rect 6039 21865 6125 21921
rect 6181 21865 6267 21921
rect 6323 21865 6409 21921
rect 6465 21865 6551 21921
rect 6607 21865 6693 21921
rect 6749 21865 6835 21921
rect 6891 21865 6977 21921
rect 7033 21865 7119 21921
rect 7175 21865 7261 21921
rect 7317 21865 7403 21921
rect 7459 21865 7545 21921
rect 7601 21865 7687 21921
rect 7743 21865 7829 21921
rect 7885 21865 7971 21921
rect 8027 21865 8113 21921
rect 8169 21865 8255 21921
rect 8311 21865 8397 21921
rect 8453 21865 8539 21921
rect 8595 21865 8681 21921
rect 8737 21865 8823 21921
rect 8879 21865 8965 21921
rect 9021 21865 9107 21921
rect 9163 21865 9249 21921
rect 9305 21865 9391 21921
rect 9447 21865 9533 21921
rect 9589 21865 9675 21921
rect 9731 21865 9817 21921
rect 9873 21865 9959 21921
rect 10015 21865 10101 21921
rect 10157 21865 10243 21921
rect 10299 21865 10385 21921
rect 10441 21865 10527 21921
rect 10583 21865 10669 21921
rect 10725 21865 10811 21921
rect 10867 21865 10953 21921
rect 11009 21865 11095 21921
rect 11151 21865 11237 21921
rect 11293 21865 11379 21921
rect 11435 21865 11521 21921
rect 11577 21865 11663 21921
rect 11719 21865 11805 21921
rect 11861 21865 11947 21921
rect 12003 21865 12089 21921
rect 12145 21865 12231 21921
rect 12287 21865 12373 21921
rect 12429 21865 12515 21921
rect 12571 21865 12657 21921
rect 12713 21865 12799 21921
rect 12855 21865 12941 21921
rect 12997 21865 13083 21921
rect 13139 21865 13225 21921
rect 13281 21865 13367 21921
rect 13423 21865 13509 21921
rect 13565 21865 13651 21921
rect 13707 21865 13793 21921
rect 13849 21865 13935 21921
rect 13991 21865 14077 21921
rect 14133 21865 14219 21921
rect 14275 21865 14361 21921
rect 14417 21865 14503 21921
rect 14559 21865 14645 21921
rect 14701 21865 14787 21921
rect 14843 21865 14853 21921
rect 151 21779 14853 21865
rect 151 21723 161 21779
rect 217 21723 303 21779
rect 359 21723 445 21779
rect 501 21723 587 21779
rect 643 21723 729 21779
rect 785 21723 871 21779
rect 927 21723 1013 21779
rect 1069 21723 1155 21779
rect 1211 21723 1297 21779
rect 1353 21723 1439 21779
rect 1495 21723 1581 21779
rect 1637 21723 1723 21779
rect 1779 21723 1865 21779
rect 1921 21723 2007 21779
rect 2063 21723 2149 21779
rect 2205 21723 2291 21779
rect 2347 21723 2433 21779
rect 2489 21723 2575 21779
rect 2631 21723 2717 21779
rect 2773 21723 2859 21779
rect 2915 21723 3001 21779
rect 3057 21723 3143 21779
rect 3199 21723 3285 21779
rect 3341 21723 3427 21779
rect 3483 21723 3569 21779
rect 3625 21723 3711 21779
rect 3767 21723 3853 21779
rect 3909 21723 3995 21779
rect 4051 21723 4137 21779
rect 4193 21723 4279 21779
rect 4335 21723 4421 21779
rect 4477 21723 4563 21779
rect 4619 21723 4705 21779
rect 4761 21723 4847 21779
rect 4903 21723 4989 21779
rect 5045 21723 5131 21779
rect 5187 21723 5273 21779
rect 5329 21723 5415 21779
rect 5471 21723 5557 21779
rect 5613 21723 5699 21779
rect 5755 21723 5841 21779
rect 5897 21723 5983 21779
rect 6039 21723 6125 21779
rect 6181 21723 6267 21779
rect 6323 21723 6409 21779
rect 6465 21723 6551 21779
rect 6607 21723 6693 21779
rect 6749 21723 6835 21779
rect 6891 21723 6977 21779
rect 7033 21723 7119 21779
rect 7175 21723 7261 21779
rect 7317 21723 7403 21779
rect 7459 21723 7545 21779
rect 7601 21723 7687 21779
rect 7743 21723 7829 21779
rect 7885 21723 7971 21779
rect 8027 21723 8113 21779
rect 8169 21723 8255 21779
rect 8311 21723 8397 21779
rect 8453 21723 8539 21779
rect 8595 21723 8681 21779
rect 8737 21723 8823 21779
rect 8879 21723 8965 21779
rect 9021 21723 9107 21779
rect 9163 21723 9249 21779
rect 9305 21723 9391 21779
rect 9447 21723 9533 21779
rect 9589 21723 9675 21779
rect 9731 21723 9817 21779
rect 9873 21723 9959 21779
rect 10015 21723 10101 21779
rect 10157 21723 10243 21779
rect 10299 21723 10385 21779
rect 10441 21723 10527 21779
rect 10583 21723 10669 21779
rect 10725 21723 10811 21779
rect 10867 21723 10953 21779
rect 11009 21723 11095 21779
rect 11151 21723 11237 21779
rect 11293 21723 11379 21779
rect 11435 21723 11521 21779
rect 11577 21723 11663 21779
rect 11719 21723 11805 21779
rect 11861 21723 11947 21779
rect 12003 21723 12089 21779
rect 12145 21723 12231 21779
rect 12287 21723 12373 21779
rect 12429 21723 12515 21779
rect 12571 21723 12657 21779
rect 12713 21723 12799 21779
rect 12855 21723 12941 21779
rect 12997 21723 13083 21779
rect 13139 21723 13225 21779
rect 13281 21723 13367 21779
rect 13423 21723 13509 21779
rect 13565 21723 13651 21779
rect 13707 21723 13793 21779
rect 13849 21723 13935 21779
rect 13991 21723 14077 21779
rect 14133 21723 14219 21779
rect 14275 21723 14361 21779
rect 14417 21723 14503 21779
rect 14559 21723 14645 21779
rect 14701 21723 14787 21779
rect 14843 21723 14853 21779
rect 151 21637 14853 21723
rect 151 21581 161 21637
rect 217 21581 303 21637
rect 359 21581 445 21637
rect 501 21581 587 21637
rect 643 21581 729 21637
rect 785 21581 871 21637
rect 927 21581 1013 21637
rect 1069 21581 1155 21637
rect 1211 21581 1297 21637
rect 1353 21581 1439 21637
rect 1495 21581 1581 21637
rect 1637 21581 1723 21637
rect 1779 21581 1865 21637
rect 1921 21581 2007 21637
rect 2063 21581 2149 21637
rect 2205 21581 2291 21637
rect 2347 21581 2433 21637
rect 2489 21581 2575 21637
rect 2631 21581 2717 21637
rect 2773 21581 2859 21637
rect 2915 21581 3001 21637
rect 3057 21581 3143 21637
rect 3199 21581 3285 21637
rect 3341 21581 3427 21637
rect 3483 21581 3569 21637
rect 3625 21581 3711 21637
rect 3767 21581 3853 21637
rect 3909 21581 3995 21637
rect 4051 21581 4137 21637
rect 4193 21581 4279 21637
rect 4335 21581 4421 21637
rect 4477 21581 4563 21637
rect 4619 21581 4705 21637
rect 4761 21581 4847 21637
rect 4903 21581 4989 21637
rect 5045 21581 5131 21637
rect 5187 21581 5273 21637
rect 5329 21581 5415 21637
rect 5471 21581 5557 21637
rect 5613 21581 5699 21637
rect 5755 21581 5841 21637
rect 5897 21581 5983 21637
rect 6039 21581 6125 21637
rect 6181 21581 6267 21637
rect 6323 21581 6409 21637
rect 6465 21581 6551 21637
rect 6607 21581 6693 21637
rect 6749 21581 6835 21637
rect 6891 21581 6977 21637
rect 7033 21581 7119 21637
rect 7175 21581 7261 21637
rect 7317 21581 7403 21637
rect 7459 21581 7545 21637
rect 7601 21581 7687 21637
rect 7743 21581 7829 21637
rect 7885 21581 7971 21637
rect 8027 21581 8113 21637
rect 8169 21581 8255 21637
rect 8311 21581 8397 21637
rect 8453 21581 8539 21637
rect 8595 21581 8681 21637
rect 8737 21581 8823 21637
rect 8879 21581 8965 21637
rect 9021 21581 9107 21637
rect 9163 21581 9249 21637
rect 9305 21581 9391 21637
rect 9447 21581 9533 21637
rect 9589 21581 9675 21637
rect 9731 21581 9817 21637
rect 9873 21581 9959 21637
rect 10015 21581 10101 21637
rect 10157 21581 10243 21637
rect 10299 21581 10385 21637
rect 10441 21581 10527 21637
rect 10583 21581 10669 21637
rect 10725 21581 10811 21637
rect 10867 21581 10953 21637
rect 11009 21581 11095 21637
rect 11151 21581 11237 21637
rect 11293 21581 11379 21637
rect 11435 21581 11521 21637
rect 11577 21581 11663 21637
rect 11719 21581 11805 21637
rect 11861 21581 11947 21637
rect 12003 21581 12089 21637
rect 12145 21581 12231 21637
rect 12287 21581 12373 21637
rect 12429 21581 12515 21637
rect 12571 21581 12657 21637
rect 12713 21581 12799 21637
rect 12855 21581 12941 21637
rect 12997 21581 13083 21637
rect 13139 21581 13225 21637
rect 13281 21581 13367 21637
rect 13423 21581 13509 21637
rect 13565 21581 13651 21637
rect 13707 21581 13793 21637
rect 13849 21581 13935 21637
rect 13991 21581 14077 21637
rect 14133 21581 14219 21637
rect 14275 21581 14361 21637
rect 14417 21581 14503 21637
rect 14559 21581 14645 21637
rect 14701 21581 14787 21637
rect 14843 21581 14853 21637
rect 151 21495 14853 21581
rect 151 21439 161 21495
rect 217 21439 303 21495
rect 359 21439 445 21495
rect 501 21439 587 21495
rect 643 21439 729 21495
rect 785 21439 871 21495
rect 927 21439 1013 21495
rect 1069 21439 1155 21495
rect 1211 21439 1297 21495
rect 1353 21439 1439 21495
rect 1495 21439 1581 21495
rect 1637 21439 1723 21495
rect 1779 21439 1865 21495
rect 1921 21439 2007 21495
rect 2063 21439 2149 21495
rect 2205 21439 2291 21495
rect 2347 21439 2433 21495
rect 2489 21439 2575 21495
rect 2631 21439 2717 21495
rect 2773 21439 2859 21495
rect 2915 21439 3001 21495
rect 3057 21439 3143 21495
rect 3199 21439 3285 21495
rect 3341 21439 3427 21495
rect 3483 21439 3569 21495
rect 3625 21439 3711 21495
rect 3767 21439 3853 21495
rect 3909 21439 3995 21495
rect 4051 21439 4137 21495
rect 4193 21439 4279 21495
rect 4335 21439 4421 21495
rect 4477 21439 4563 21495
rect 4619 21439 4705 21495
rect 4761 21439 4847 21495
rect 4903 21439 4989 21495
rect 5045 21439 5131 21495
rect 5187 21439 5273 21495
rect 5329 21439 5415 21495
rect 5471 21439 5557 21495
rect 5613 21439 5699 21495
rect 5755 21439 5841 21495
rect 5897 21439 5983 21495
rect 6039 21439 6125 21495
rect 6181 21439 6267 21495
rect 6323 21439 6409 21495
rect 6465 21439 6551 21495
rect 6607 21439 6693 21495
rect 6749 21439 6835 21495
rect 6891 21439 6977 21495
rect 7033 21439 7119 21495
rect 7175 21439 7261 21495
rect 7317 21439 7403 21495
rect 7459 21439 7545 21495
rect 7601 21439 7687 21495
rect 7743 21439 7829 21495
rect 7885 21439 7971 21495
rect 8027 21439 8113 21495
rect 8169 21439 8255 21495
rect 8311 21439 8397 21495
rect 8453 21439 8539 21495
rect 8595 21439 8681 21495
rect 8737 21439 8823 21495
rect 8879 21439 8965 21495
rect 9021 21439 9107 21495
rect 9163 21439 9249 21495
rect 9305 21439 9391 21495
rect 9447 21439 9533 21495
rect 9589 21439 9675 21495
rect 9731 21439 9817 21495
rect 9873 21439 9959 21495
rect 10015 21439 10101 21495
rect 10157 21439 10243 21495
rect 10299 21439 10385 21495
rect 10441 21439 10527 21495
rect 10583 21439 10669 21495
rect 10725 21439 10811 21495
rect 10867 21439 10953 21495
rect 11009 21439 11095 21495
rect 11151 21439 11237 21495
rect 11293 21439 11379 21495
rect 11435 21439 11521 21495
rect 11577 21439 11663 21495
rect 11719 21439 11805 21495
rect 11861 21439 11947 21495
rect 12003 21439 12089 21495
rect 12145 21439 12231 21495
rect 12287 21439 12373 21495
rect 12429 21439 12515 21495
rect 12571 21439 12657 21495
rect 12713 21439 12799 21495
rect 12855 21439 12941 21495
rect 12997 21439 13083 21495
rect 13139 21439 13225 21495
rect 13281 21439 13367 21495
rect 13423 21439 13509 21495
rect 13565 21439 13651 21495
rect 13707 21439 13793 21495
rect 13849 21439 13935 21495
rect 13991 21439 14077 21495
rect 14133 21439 14219 21495
rect 14275 21439 14361 21495
rect 14417 21439 14503 21495
rect 14559 21439 14645 21495
rect 14701 21439 14787 21495
rect 14843 21439 14853 21495
rect 151 21353 14853 21439
rect 151 21297 161 21353
rect 217 21297 303 21353
rect 359 21297 445 21353
rect 501 21297 587 21353
rect 643 21297 729 21353
rect 785 21297 871 21353
rect 927 21297 1013 21353
rect 1069 21297 1155 21353
rect 1211 21297 1297 21353
rect 1353 21297 1439 21353
rect 1495 21297 1581 21353
rect 1637 21297 1723 21353
rect 1779 21297 1865 21353
rect 1921 21297 2007 21353
rect 2063 21297 2149 21353
rect 2205 21297 2291 21353
rect 2347 21297 2433 21353
rect 2489 21297 2575 21353
rect 2631 21297 2717 21353
rect 2773 21297 2859 21353
rect 2915 21297 3001 21353
rect 3057 21297 3143 21353
rect 3199 21297 3285 21353
rect 3341 21297 3427 21353
rect 3483 21297 3569 21353
rect 3625 21297 3711 21353
rect 3767 21297 3853 21353
rect 3909 21297 3995 21353
rect 4051 21297 4137 21353
rect 4193 21297 4279 21353
rect 4335 21297 4421 21353
rect 4477 21297 4563 21353
rect 4619 21297 4705 21353
rect 4761 21297 4847 21353
rect 4903 21297 4989 21353
rect 5045 21297 5131 21353
rect 5187 21297 5273 21353
rect 5329 21297 5415 21353
rect 5471 21297 5557 21353
rect 5613 21297 5699 21353
rect 5755 21297 5841 21353
rect 5897 21297 5983 21353
rect 6039 21297 6125 21353
rect 6181 21297 6267 21353
rect 6323 21297 6409 21353
rect 6465 21297 6551 21353
rect 6607 21297 6693 21353
rect 6749 21297 6835 21353
rect 6891 21297 6977 21353
rect 7033 21297 7119 21353
rect 7175 21297 7261 21353
rect 7317 21297 7403 21353
rect 7459 21297 7545 21353
rect 7601 21297 7687 21353
rect 7743 21297 7829 21353
rect 7885 21297 7971 21353
rect 8027 21297 8113 21353
rect 8169 21297 8255 21353
rect 8311 21297 8397 21353
rect 8453 21297 8539 21353
rect 8595 21297 8681 21353
rect 8737 21297 8823 21353
rect 8879 21297 8965 21353
rect 9021 21297 9107 21353
rect 9163 21297 9249 21353
rect 9305 21297 9391 21353
rect 9447 21297 9533 21353
rect 9589 21297 9675 21353
rect 9731 21297 9817 21353
rect 9873 21297 9959 21353
rect 10015 21297 10101 21353
rect 10157 21297 10243 21353
rect 10299 21297 10385 21353
rect 10441 21297 10527 21353
rect 10583 21297 10669 21353
rect 10725 21297 10811 21353
rect 10867 21297 10953 21353
rect 11009 21297 11095 21353
rect 11151 21297 11237 21353
rect 11293 21297 11379 21353
rect 11435 21297 11521 21353
rect 11577 21297 11663 21353
rect 11719 21297 11805 21353
rect 11861 21297 11947 21353
rect 12003 21297 12089 21353
rect 12145 21297 12231 21353
rect 12287 21297 12373 21353
rect 12429 21297 12515 21353
rect 12571 21297 12657 21353
rect 12713 21297 12799 21353
rect 12855 21297 12941 21353
rect 12997 21297 13083 21353
rect 13139 21297 13225 21353
rect 13281 21297 13367 21353
rect 13423 21297 13509 21353
rect 13565 21297 13651 21353
rect 13707 21297 13793 21353
rect 13849 21297 13935 21353
rect 13991 21297 14077 21353
rect 14133 21297 14219 21353
rect 14275 21297 14361 21353
rect 14417 21297 14503 21353
rect 14559 21297 14645 21353
rect 14701 21297 14787 21353
rect 14843 21297 14853 21353
rect 151 21211 14853 21297
rect 151 21155 161 21211
rect 217 21155 303 21211
rect 359 21155 445 21211
rect 501 21155 587 21211
rect 643 21155 729 21211
rect 785 21155 871 21211
rect 927 21155 1013 21211
rect 1069 21155 1155 21211
rect 1211 21155 1297 21211
rect 1353 21155 1439 21211
rect 1495 21155 1581 21211
rect 1637 21155 1723 21211
rect 1779 21155 1865 21211
rect 1921 21155 2007 21211
rect 2063 21155 2149 21211
rect 2205 21155 2291 21211
rect 2347 21155 2433 21211
rect 2489 21155 2575 21211
rect 2631 21155 2717 21211
rect 2773 21155 2859 21211
rect 2915 21155 3001 21211
rect 3057 21155 3143 21211
rect 3199 21155 3285 21211
rect 3341 21155 3427 21211
rect 3483 21155 3569 21211
rect 3625 21155 3711 21211
rect 3767 21155 3853 21211
rect 3909 21155 3995 21211
rect 4051 21155 4137 21211
rect 4193 21155 4279 21211
rect 4335 21155 4421 21211
rect 4477 21155 4563 21211
rect 4619 21155 4705 21211
rect 4761 21155 4847 21211
rect 4903 21155 4989 21211
rect 5045 21155 5131 21211
rect 5187 21155 5273 21211
rect 5329 21155 5415 21211
rect 5471 21155 5557 21211
rect 5613 21155 5699 21211
rect 5755 21155 5841 21211
rect 5897 21155 5983 21211
rect 6039 21155 6125 21211
rect 6181 21155 6267 21211
rect 6323 21155 6409 21211
rect 6465 21155 6551 21211
rect 6607 21155 6693 21211
rect 6749 21155 6835 21211
rect 6891 21155 6977 21211
rect 7033 21155 7119 21211
rect 7175 21155 7261 21211
rect 7317 21155 7403 21211
rect 7459 21155 7545 21211
rect 7601 21155 7687 21211
rect 7743 21155 7829 21211
rect 7885 21155 7971 21211
rect 8027 21155 8113 21211
rect 8169 21155 8255 21211
rect 8311 21155 8397 21211
rect 8453 21155 8539 21211
rect 8595 21155 8681 21211
rect 8737 21155 8823 21211
rect 8879 21155 8965 21211
rect 9021 21155 9107 21211
rect 9163 21155 9249 21211
rect 9305 21155 9391 21211
rect 9447 21155 9533 21211
rect 9589 21155 9675 21211
rect 9731 21155 9817 21211
rect 9873 21155 9959 21211
rect 10015 21155 10101 21211
rect 10157 21155 10243 21211
rect 10299 21155 10385 21211
rect 10441 21155 10527 21211
rect 10583 21155 10669 21211
rect 10725 21155 10811 21211
rect 10867 21155 10953 21211
rect 11009 21155 11095 21211
rect 11151 21155 11237 21211
rect 11293 21155 11379 21211
rect 11435 21155 11521 21211
rect 11577 21155 11663 21211
rect 11719 21155 11805 21211
rect 11861 21155 11947 21211
rect 12003 21155 12089 21211
rect 12145 21155 12231 21211
rect 12287 21155 12373 21211
rect 12429 21155 12515 21211
rect 12571 21155 12657 21211
rect 12713 21155 12799 21211
rect 12855 21155 12941 21211
rect 12997 21155 13083 21211
rect 13139 21155 13225 21211
rect 13281 21155 13367 21211
rect 13423 21155 13509 21211
rect 13565 21155 13651 21211
rect 13707 21155 13793 21211
rect 13849 21155 13935 21211
rect 13991 21155 14077 21211
rect 14133 21155 14219 21211
rect 14275 21155 14361 21211
rect 14417 21155 14503 21211
rect 14559 21155 14645 21211
rect 14701 21155 14787 21211
rect 14843 21155 14853 21211
rect 151 21069 14853 21155
rect 151 21013 161 21069
rect 217 21013 303 21069
rect 359 21013 445 21069
rect 501 21013 587 21069
rect 643 21013 729 21069
rect 785 21013 871 21069
rect 927 21013 1013 21069
rect 1069 21013 1155 21069
rect 1211 21013 1297 21069
rect 1353 21013 1439 21069
rect 1495 21013 1581 21069
rect 1637 21013 1723 21069
rect 1779 21013 1865 21069
rect 1921 21013 2007 21069
rect 2063 21013 2149 21069
rect 2205 21013 2291 21069
rect 2347 21013 2433 21069
rect 2489 21013 2575 21069
rect 2631 21013 2717 21069
rect 2773 21013 2859 21069
rect 2915 21013 3001 21069
rect 3057 21013 3143 21069
rect 3199 21013 3285 21069
rect 3341 21013 3427 21069
rect 3483 21013 3569 21069
rect 3625 21013 3711 21069
rect 3767 21013 3853 21069
rect 3909 21013 3995 21069
rect 4051 21013 4137 21069
rect 4193 21013 4279 21069
rect 4335 21013 4421 21069
rect 4477 21013 4563 21069
rect 4619 21013 4705 21069
rect 4761 21013 4847 21069
rect 4903 21013 4989 21069
rect 5045 21013 5131 21069
rect 5187 21013 5273 21069
rect 5329 21013 5415 21069
rect 5471 21013 5557 21069
rect 5613 21013 5699 21069
rect 5755 21013 5841 21069
rect 5897 21013 5983 21069
rect 6039 21013 6125 21069
rect 6181 21013 6267 21069
rect 6323 21013 6409 21069
rect 6465 21013 6551 21069
rect 6607 21013 6693 21069
rect 6749 21013 6835 21069
rect 6891 21013 6977 21069
rect 7033 21013 7119 21069
rect 7175 21013 7261 21069
rect 7317 21013 7403 21069
rect 7459 21013 7545 21069
rect 7601 21013 7687 21069
rect 7743 21013 7829 21069
rect 7885 21013 7971 21069
rect 8027 21013 8113 21069
rect 8169 21013 8255 21069
rect 8311 21013 8397 21069
rect 8453 21013 8539 21069
rect 8595 21013 8681 21069
rect 8737 21013 8823 21069
rect 8879 21013 8965 21069
rect 9021 21013 9107 21069
rect 9163 21013 9249 21069
rect 9305 21013 9391 21069
rect 9447 21013 9533 21069
rect 9589 21013 9675 21069
rect 9731 21013 9817 21069
rect 9873 21013 9959 21069
rect 10015 21013 10101 21069
rect 10157 21013 10243 21069
rect 10299 21013 10385 21069
rect 10441 21013 10527 21069
rect 10583 21013 10669 21069
rect 10725 21013 10811 21069
rect 10867 21013 10953 21069
rect 11009 21013 11095 21069
rect 11151 21013 11237 21069
rect 11293 21013 11379 21069
rect 11435 21013 11521 21069
rect 11577 21013 11663 21069
rect 11719 21013 11805 21069
rect 11861 21013 11947 21069
rect 12003 21013 12089 21069
rect 12145 21013 12231 21069
rect 12287 21013 12373 21069
rect 12429 21013 12515 21069
rect 12571 21013 12657 21069
rect 12713 21013 12799 21069
rect 12855 21013 12941 21069
rect 12997 21013 13083 21069
rect 13139 21013 13225 21069
rect 13281 21013 13367 21069
rect 13423 21013 13509 21069
rect 13565 21013 13651 21069
rect 13707 21013 13793 21069
rect 13849 21013 13935 21069
rect 13991 21013 14077 21069
rect 14133 21013 14219 21069
rect 14275 21013 14361 21069
rect 14417 21013 14503 21069
rect 14559 21013 14645 21069
rect 14701 21013 14787 21069
rect 14843 21013 14853 21069
rect 151 20927 14853 21013
rect 151 20871 161 20927
rect 217 20871 303 20927
rect 359 20871 445 20927
rect 501 20871 587 20927
rect 643 20871 729 20927
rect 785 20871 871 20927
rect 927 20871 1013 20927
rect 1069 20871 1155 20927
rect 1211 20871 1297 20927
rect 1353 20871 1439 20927
rect 1495 20871 1581 20927
rect 1637 20871 1723 20927
rect 1779 20871 1865 20927
rect 1921 20871 2007 20927
rect 2063 20871 2149 20927
rect 2205 20871 2291 20927
rect 2347 20871 2433 20927
rect 2489 20871 2575 20927
rect 2631 20871 2717 20927
rect 2773 20871 2859 20927
rect 2915 20871 3001 20927
rect 3057 20871 3143 20927
rect 3199 20871 3285 20927
rect 3341 20871 3427 20927
rect 3483 20871 3569 20927
rect 3625 20871 3711 20927
rect 3767 20871 3853 20927
rect 3909 20871 3995 20927
rect 4051 20871 4137 20927
rect 4193 20871 4279 20927
rect 4335 20871 4421 20927
rect 4477 20871 4563 20927
rect 4619 20871 4705 20927
rect 4761 20871 4847 20927
rect 4903 20871 4989 20927
rect 5045 20871 5131 20927
rect 5187 20871 5273 20927
rect 5329 20871 5415 20927
rect 5471 20871 5557 20927
rect 5613 20871 5699 20927
rect 5755 20871 5841 20927
rect 5897 20871 5983 20927
rect 6039 20871 6125 20927
rect 6181 20871 6267 20927
rect 6323 20871 6409 20927
rect 6465 20871 6551 20927
rect 6607 20871 6693 20927
rect 6749 20871 6835 20927
rect 6891 20871 6977 20927
rect 7033 20871 7119 20927
rect 7175 20871 7261 20927
rect 7317 20871 7403 20927
rect 7459 20871 7545 20927
rect 7601 20871 7687 20927
rect 7743 20871 7829 20927
rect 7885 20871 7971 20927
rect 8027 20871 8113 20927
rect 8169 20871 8255 20927
rect 8311 20871 8397 20927
rect 8453 20871 8539 20927
rect 8595 20871 8681 20927
rect 8737 20871 8823 20927
rect 8879 20871 8965 20927
rect 9021 20871 9107 20927
rect 9163 20871 9249 20927
rect 9305 20871 9391 20927
rect 9447 20871 9533 20927
rect 9589 20871 9675 20927
rect 9731 20871 9817 20927
rect 9873 20871 9959 20927
rect 10015 20871 10101 20927
rect 10157 20871 10243 20927
rect 10299 20871 10385 20927
rect 10441 20871 10527 20927
rect 10583 20871 10669 20927
rect 10725 20871 10811 20927
rect 10867 20871 10953 20927
rect 11009 20871 11095 20927
rect 11151 20871 11237 20927
rect 11293 20871 11379 20927
rect 11435 20871 11521 20927
rect 11577 20871 11663 20927
rect 11719 20871 11805 20927
rect 11861 20871 11947 20927
rect 12003 20871 12089 20927
rect 12145 20871 12231 20927
rect 12287 20871 12373 20927
rect 12429 20871 12515 20927
rect 12571 20871 12657 20927
rect 12713 20871 12799 20927
rect 12855 20871 12941 20927
rect 12997 20871 13083 20927
rect 13139 20871 13225 20927
rect 13281 20871 13367 20927
rect 13423 20871 13509 20927
rect 13565 20871 13651 20927
rect 13707 20871 13793 20927
rect 13849 20871 13935 20927
rect 13991 20871 14077 20927
rect 14133 20871 14219 20927
rect 14275 20871 14361 20927
rect 14417 20871 14503 20927
rect 14559 20871 14645 20927
rect 14701 20871 14787 20927
rect 14843 20871 14853 20927
rect 151 20785 14853 20871
rect 151 20729 161 20785
rect 217 20729 303 20785
rect 359 20729 445 20785
rect 501 20729 587 20785
rect 643 20729 729 20785
rect 785 20729 871 20785
rect 927 20729 1013 20785
rect 1069 20729 1155 20785
rect 1211 20729 1297 20785
rect 1353 20729 1439 20785
rect 1495 20729 1581 20785
rect 1637 20729 1723 20785
rect 1779 20729 1865 20785
rect 1921 20729 2007 20785
rect 2063 20729 2149 20785
rect 2205 20729 2291 20785
rect 2347 20729 2433 20785
rect 2489 20729 2575 20785
rect 2631 20729 2717 20785
rect 2773 20729 2859 20785
rect 2915 20729 3001 20785
rect 3057 20729 3143 20785
rect 3199 20729 3285 20785
rect 3341 20729 3427 20785
rect 3483 20729 3569 20785
rect 3625 20729 3711 20785
rect 3767 20729 3853 20785
rect 3909 20729 3995 20785
rect 4051 20729 4137 20785
rect 4193 20729 4279 20785
rect 4335 20729 4421 20785
rect 4477 20729 4563 20785
rect 4619 20729 4705 20785
rect 4761 20729 4847 20785
rect 4903 20729 4989 20785
rect 5045 20729 5131 20785
rect 5187 20729 5273 20785
rect 5329 20729 5415 20785
rect 5471 20729 5557 20785
rect 5613 20729 5699 20785
rect 5755 20729 5841 20785
rect 5897 20729 5983 20785
rect 6039 20729 6125 20785
rect 6181 20729 6267 20785
rect 6323 20729 6409 20785
rect 6465 20729 6551 20785
rect 6607 20729 6693 20785
rect 6749 20729 6835 20785
rect 6891 20729 6977 20785
rect 7033 20729 7119 20785
rect 7175 20729 7261 20785
rect 7317 20729 7403 20785
rect 7459 20729 7545 20785
rect 7601 20729 7687 20785
rect 7743 20729 7829 20785
rect 7885 20729 7971 20785
rect 8027 20729 8113 20785
rect 8169 20729 8255 20785
rect 8311 20729 8397 20785
rect 8453 20729 8539 20785
rect 8595 20729 8681 20785
rect 8737 20729 8823 20785
rect 8879 20729 8965 20785
rect 9021 20729 9107 20785
rect 9163 20729 9249 20785
rect 9305 20729 9391 20785
rect 9447 20729 9533 20785
rect 9589 20729 9675 20785
rect 9731 20729 9817 20785
rect 9873 20729 9959 20785
rect 10015 20729 10101 20785
rect 10157 20729 10243 20785
rect 10299 20729 10385 20785
rect 10441 20729 10527 20785
rect 10583 20729 10669 20785
rect 10725 20729 10811 20785
rect 10867 20729 10953 20785
rect 11009 20729 11095 20785
rect 11151 20729 11237 20785
rect 11293 20729 11379 20785
rect 11435 20729 11521 20785
rect 11577 20729 11663 20785
rect 11719 20729 11805 20785
rect 11861 20729 11947 20785
rect 12003 20729 12089 20785
rect 12145 20729 12231 20785
rect 12287 20729 12373 20785
rect 12429 20729 12515 20785
rect 12571 20729 12657 20785
rect 12713 20729 12799 20785
rect 12855 20729 12941 20785
rect 12997 20729 13083 20785
rect 13139 20729 13225 20785
rect 13281 20729 13367 20785
rect 13423 20729 13509 20785
rect 13565 20729 13651 20785
rect 13707 20729 13793 20785
rect 13849 20729 13935 20785
rect 13991 20729 14077 20785
rect 14133 20729 14219 20785
rect 14275 20729 14361 20785
rect 14417 20729 14503 20785
rect 14559 20729 14645 20785
rect 14701 20729 14787 20785
rect 14843 20729 14853 20785
rect 151 20643 14853 20729
rect 151 20587 161 20643
rect 217 20587 303 20643
rect 359 20587 445 20643
rect 501 20587 587 20643
rect 643 20587 729 20643
rect 785 20587 871 20643
rect 927 20587 1013 20643
rect 1069 20587 1155 20643
rect 1211 20587 1297 20643
rect 1353 20587 1439 20643
rect 1495 20587 1581 20643
rect 1637 20587 1723 20643
rect 1779 20587 1865 20643
rect 1921 20587 2007 20643
rect 2063 20587 2149 20643
rect 2205 20587 2291 20643
rect 2347 20587 2433 20643
rect 2489 20587 2575 20643
rect 2631 20587 2717 20643
rect 2773 20587 2859 20643
rect 2915 20587 3001 20643
rect 3057 20587 3143 20643
rect 3199 20587 3285 20643
rect 3341 20587 3427 20643
rect 3483 20587 3569 20643
rect 3625 20587 3711 20643
rect 3767 20587 3853 20643
rect 3909 20587 3995 20643
rect 4051 20587 4137 20643
rect 4193 20587 4279 20643
rect 4335 20587 4421 20643
rect 4477 20587 4563 20643
rect 4619 20587 4705 20643
rect 4761 20587 4847 20643
rect 4903 20587 4989 20643
rect 5045 20587 5131 20643
rect 5187 20587 5273 20643
rect 5329 20587 5415 20643
rect 5471 20587 5557 20643
rect 5613 20587 5699 20643
rect 5755 20587 5841 20643
rect 5897 20587 5983 20643
rect 6039 20587 6125 20643
rect 6181 20587 6267 20643
rect 6323 20587 6409 20643
rect 6465 20587 6551 20643
rect 6607 20587 6693 20643
rect 6749 20587 6835 20643
rect 6891 20587 6977 20643
rect 7033 20587 7119 20643
rect 7175 20587 7261 20643
rect 7317 20587 7403 20643
rect 7459 20587 7545 20643
rect 7601 20587 7687 20643
rect 7743 20587 7829 20643
rect 7885 20587 7971 20643
rect 8027 20587 8113 20643
rect 8169 20587 8255 20643
rect 8311 20587 8397 20643
rect 8453 20587 8539 20643
rect 8595 20587 8681 20643
rect 8737 20587 8823 20643
rect 8879 20587 8965 20643
rect 9021 20587 9107 20643
rect 9163 20587 9249 20643
rect 9305 20587 9391 20643
rect 9447 20587 9533 20643
rect 9589 20587 9675 20643
rect 9731 20587 9817 20643
rect 9873 20587 9959 20643
rect 10015 20587 10101 20643
rect 10157 20587 10243 20643
rect 10299 20587 10385 20643
rect 10441 20587 10527 20643
rect 10583 20587 10669 20643
rect 10725 20587 10811 20643
rect 10867 20587 10953 20643
rect 11009 20587 11095 20643
rect 11151 20587 11237 20643
rect 11293 20587 11379 20643
rect 11435 20587 11521 20643
rect 11577 20587 11663 20643
rect 11719 20587 11805 20643
rect 11861 20587 11947 20643
rect 12003 20587 12089 20643
rect 12145 20587 12231 20643
rect 12287 20587 12373 20643
rect 12429 20587 12515 20643
rect 12571 20587 12657 20643
rect 12713 20587 12799 20643
rect 12855 20587 12941 20643
rect 12997 20587 13083 20643
rect 13139 20587 13225 20643
rect 13281 20587 13367 20643
rect 13423 20587 13509 20643
rect 13565 20587 13651 20643
rect 13707 20587 13793 20643
rect 13849 20587 13935 20643
rect 13991 20587 14077 20643
rect 14133 20587 14219 20643
rect 14275 20587 14361 20643
rect 14417 20587 14503 20643
rect 14559 20587 14645 20643
rect 14701 20587 14787 20643
rect 14843 20587 14853 20643
rect 151 20501 14853 20587
rect 151 20445 161 20501
rect 217 20445 303 20501
rect 359 20445 445 20501
rect 501 20445 587 20501
rect 643 20445 729 20501
rect 785 20445 871 20501
rect 927 20445 1013 20501
rect 1069 20445 1155 20501
rect 1211 20445 1297 20501
rect 1353 20445 1439 20501
rect 1495 20445 1581 20501
rect 1637 20445 1723 20501
rect 1779 20445 1865 20501
rect 1921 20445 2007 20501
rect 2063 20445 2149 20501
rect 2205 20445 2291 20501
rect 2347 20445 2433 20501
rect 2489 20445 2575 20501
rect 2631 20445 2717 20501
rect 2773 20445 2859 20501
rect 2915 20445 3001 20501
rect 3057 20445 3143 20501
rect 3199 20445 3285 20501
rect 3341 20445 3427 20501
rect 3483 20445 3569 20501
rect 3625 20445 3711 20501
rect 3767 20445 3853 20501
rect 3909 20445 3995 20501
rect 4051 20445 4137 20501
rect 4193 20445 4279 20501
rect 4335 20445 4421 20501
rect 4477 20445 4563 20501
rect 4619 20445 4705 20501
rect 4761 20445 4847 20501
rect 4903 20445 4989 20501
rect 5045 20445 5131 20501
rect 5187 20445 5273 20501
rect 5329 20445 5415 20501
rect 5471 20445 5557 20501
rect 5613 20445 5699 20501
rect 5755 20445 5841 20501
rect 5897 20445 5983 20501
rect 6039 20445 6125 20501
rect 6181 20445 6267 20501
rect 6323 20445 6409 20501
rect 6465 20445 6551 20501
rect 6607 20445 6693 20501
rect 6749 20445 6835 20501
rect 6891 20445 6977 20501
rect 7033 20445 7119 20501
rect 7175 20445 7261 20501
rect 7317 20445 7403 20501
rect 7459 20445 7545 20501
rect 7601 20445 7687 20501
rect 7743 20445 7829 20501
rect 7885 20445 7971 20501
rect 8027 20445 8113 20501
rect 8169 20445 8255 20501
rect 8311 20445 8397 20501
rect 8453 20445 8539 20501
rect 8595 20445 8681 20501
rect 8737 20445 8823 20501
rect 8879 20445 8965 20501
rect 9021 20445 9107 20501
rect 9163 20445 9249 20501
rect 9305 20445 9391 20501
rect 9447 20445 9533 20501
rect 9589 20445 9675 20501
rect 9731 20445 9817 20501
rect 9873 20445 9959 20501
rect 10015 20445 10101 20501
rect 10157 20445 10243 20501
rect 10299 20445 10385 20501
rect 10441 20445 10527 20501
rect 10583 20445 10669 20501
rect 10725 20445 10811 20501
rect 10867 20445 10953 20501
rect 11009 20445 11095 20501
rect 11151 20445 11237 20501
rect 11293 20445 11379 20501
rect 11435 20445 11521 20501
rect 11577 20445 11663 20501
rect 11719 20445 11805 20501
rect 11861 20445 11947 20501
rect 12003 20445 12089 20501
rect 12145 20445 12231 20501
rect 12287 20445 12373 20501
rect 12429 20445 12515 20501
rect 12571 20445 12657 20501
rect 12713 20445 12799 20501
rect 12855 20445 12941 20501
rect 12997 20445 13083 20501
rect 13139 20445 13225 20501
rect 13281 20445 13367 20501
rect 13423 20445 13509 20501
rect 13565 20445 13651 20501
rect 13707 20445 13793 20501
rect 13849 20445 13935 20501
rect 13991 20445 14077 20501
rect 14133 20445 14219 20501
rect 14275 20445 14361 20501
rect 14417 20445 14503 20501
rect 14559 20445 14645 20501
rect 14701 20445 14787 20501
rect 14843 20445 14853 20501
rect 151 20435 14853 20445
rect 151 20141 14853 20151
rect 151 20085 161 20141
rect 217 20085 303 20141
rect 359 20085 445 20141
rect 501 20085 587 20141
rect 643 20085 729 20141
rect 785 20085 871 20141
rect 927 20085 1013 20141
rect 1069 20085 1155 20141
rect 1211 20085 1297 20141
rect 1353 20085 1439 20141
rect 1495 20085 1581 20141
rect 1637 20085 1723 20141
rect 1779 20085 1865 20141
rect 1921 20085 2007 20141
rect 2063 20085 2149 20141
rect 2205 20085 2291 20141
rect 2347 20085 2433 20141
rect 2489 20085 2575 20141
rect 2631 20085 2717 20141
rect 2773 20085 2859 20141
rect 2915 20085 3001 20141
rect 3057 20085 3143 20141
rect 3199 20085 3285 20141
rect 3341 20085 3427 20141
rect 3483 20085 3569 20141
rect 3625 20085 3711 20141
rect 3767 20085 3853 20141
rect 3909 20085 3995 20141
rect 4051 20085 4137 20141
rect 4193 20085 4279 20141
rect 4335 20085 4421 20141
rect 4477 20085 4563 20141
rect 4619 20085 4705 20141
rect 4761 20085 4847 20141
rect 4903 20085 4989 20141
rect 5045 20085 5131 20141
rect 5187 20085 5273 20141
rect 5329 20085 5415 20141
rect 5471 20085 5557 20141
rect 5613 20085 5699 20141
rect 5755 20085 5841 20141
rect 5897 20085 5983 20141
rect 6039 20085 6125 20141
rect 6181 20085 6267 20141
rect 6323 20085 6409 20141
rect 6465 20085 6551 20141
rect 6607 20085 6693 20141
rect 6749 20085 6835 20141
rect 6891 20085 6977 20141
rect 7033 20085 7119 20141
rect 7175 20085 7261 20141
rect 7317 20085 7403 20141
rect 7459 20085 7545 20141
rect 7601 20085 7687 20141
rect 7743 20085 7829 20141
rect 7885 20085 7971 20141
rect 8027 20085 8113 20141
rect 8169 20085 8255 20141
rect 8311 20085 8397 20141
rect 8453 20085 8539 20141
rect 8595 20085 8681 20141
rect 8737 20085 8823 20141
rect 8879 20085 8965 20141
rect 9021 20085 9107 20141
rect 9163 20085 9249 20141
rect 9305 20085 9391 20141
rect 9447 20085 9533 20141
rect 9589 20085 9675 20141
rect 9731 20085 9817 20141
rect 9873 20085 9959 20141
rect 10015 20085 10101 20141
rect 10157 20085 10243 20141
rect 10299 20085 10385 20141
rect 10441 20085 10527 20141
rect 10583 20085 10669 20141
rect 10725 20085 10811 20141
rect 10867 20085 10953 20141
rect 11009 20085 11095 20141
rect 11151 20085 11237 20141
rect 11293 20085 11379 20141
rect 11435 20085 11521 20141
rect 11577 20085 11663 20141
rect 11719 20085 11805 20141
rect 11861 20085 11947 20141
rect 12003 20085 12089 20141
rect 12145 20085 12231 20141
rect 12287 20085 12373 20141
rect 12429 20085 12515 20141
rect 12571 20085 12657 20141
rect 12713 20085 12799 20141
rect 12855 20085 12941 20141
rect 12997 20085 13083 20141
rect 13139 20085 13225 20141
rect 13281 20085 13367 20141
rect 13423 20085 13509 20141
rect 13565 20085 13651 20141
rect 13707 20085 13793 20141
rect 13849 20085 13935 20141
rect 13991 20085 14077 20141
rect 14133 20085 14219 20141
rect 14275 20085 14361 20141
rect 14417 20085 14503 20141
rect 14559 20085 14645 20141
rect 14701 20085 14787 20141
rect 14843 20085 14853 20141
rect 151 19999 14853 20085
rect 151 19943 161 19999
rect 217 19943 303 19999
rect 359 19943 445 19999
rect 501 19943 587 19999
rect 643 19943 729 19999
rect 785 19943 871 19999
rect 927 19943 1013 19999
rect 1069 19943 1155 19999
rect 1211 19943 1297 19999
rect 1353 19943 1439 19999
rect 1495 19943 1581 19999
rect 1637 19943 1723 19999
rect 1779 19943 1865 19999
rect 1921 19943 2007 19999
rect 2063 19943 2149 19999
rect 2205 19943 2291 19999
rect 2347 19943 2433 19999
rect 2489 19943 2575 19999
rect 2631 19943 2717 19999
rect 2773 19943 2859 19999
rect 2915 19943 3001 19999
rect 3057 19943 3143 19999
rect 3199 19943 3285 19999
rect 3341 19943 3427 19999
rect 3483 19943 3569 19999
rect 3625 19943 3711 19999
rect 3767 19943 3853 19999
rect 3909 19943 3995 19999
rect 4051 19943 4137 19999
rect 4193 19943 4279 19999
rect 4335 19943 4421 19999
rect 4477 19943 4563 19999
rect 4619 19943 4705 19999
rect 4761 19943 4847 19999
rect 4903 19943 4989 19999
rect 5045 19943 5131 19999
rect 5187 19943 5273 19999
rect 5329 19943 5415 19999
rect 5471 19943 5557 19999
rect 5613 19943 5699 19999
rect 5755 19943 5841 19999
rect 5897 19943 5983 19999
rect 6039 19943 6125 19999
rect 6181 19943 6267 19999
rect 6323 19943 6409 19999
rect 6465 19943 6551 19999
rect 6607 19943 6693 19999
rect 6749 19943 6835 19999
rect 6891 19943 6977 19999
rect 7033 19943 7119 19999
rect 7175 19943 7261 19999
rect 7317 19943 7403 19999
rect 7459 19943 7545 19999
rect 7601 19943 7687 19999
rect 7743 19943 7829 19999
rect 7885 19943 7971 19999
rect 8027 19943 8113 19999
rect 8169 19943 8255 19999
rect 8311 19943 8397 19999
rect 8453 19943 8539 19999
rect 8595 19943 8681 19999
rect 8737 19943 8823 19999
rect 8879 19943 8965 19999
rect 9021 19943 9107 19999
rect 9163 19943 9249 19999
rect 9305 19943 9391 19999
rect 9447 19943 9533 19999
rect 9589 19943 9675 19999
rect 9731 19943 9817 19999
rect 9873 19943 9959 19999
rect 10015 19943 10101 19999
rect 10157 19943 10243 19999
rect 10299 19943 10385 19999
rect 10441 19943 10527 19999
rect 10583 19943 10669 19999
rect 10725 19943 10811 19999
rect 10867 19943 10953 19999
rect 11009 19943 11095 19999
rect 11151 19943 11237 19999
rect 11293 19943 11379 19999
rect 11435 19943 11521 19999
rect 11577 19943 11663 19999
rect 11719 19943 11805 19999
rect 11861 19943 11947 19999
rect 12003 19943 12089 19999
rect 12145 19943 12231 19999
rect 12287 19943 12373 19999
rect 12429 19943 12515 19999
rect 12571 19943 12657 19999
rect 12713 19943 12799 19999
rect 12855 19943 12941 19999
rect 12997 19943 13083 19999
rect 13139 19943 13225 19999
rect 13281 19943 13367 19999
rect 13423 19943 13509 19999
rect 13565 19943 13651 19999
rect 13707 19943 13793 19999
rect 13849 19943 13935 19999
rect 13991 19943 14077 19999
rect 14133 19943 14219 19999
rect 14275 19943 14361 19999
rect 14417 19943 14503 19999
rect 14559 19943 14645 19999
rect 14701 19943 14787 19999
rect 14843 19943 14853 19999
rect 151 19857 14853 19943
rect 151 19801 161 19857
rect 217 19801 303 19857
rect 359 19801 445 19857
rect 501 19801 587 19857
rect 643 19801 729 19857
rect 785 19801 871 19857
rect 927 19801 1013 19857
rect 1069 19801 1155 19857
rect 1211 19801 1297 19857
rect 1353 19801 1439 19857
rect 1495 19801 1581 19857
rect 1637 19801 1723 19857
rect 1779 19801 1865 19857
rect 1921 19801 2007 19857
rect 2063 19801 2149 19857
rect 2205 19801 2291 19857
rect 2347 19801 2433 19857
rect 2489 19801 2575 19857
rect 2631 19801 2717 19857
rect 2773 19801 2859 19857
rect 2915 19801 3001 19857
rect 3057 19801 3143 19857
rect 3199 19801 3285 19857
rect 3341 19801 3427 19857
rect 3483 19801 3569 19857
rect 3625 19801 3711 19857
rect 3767 19801 3853 19857
rect 3909 19801 3995 19857
rect 4051 19801 4137 19857
rect 4193 19801 4279 19857
rect 4335 19801 4421 19857
rect 4477 19801 4563 19857
rect 4619 19801 4705 19857
rect 4761 19801 4847 19857
rect 4903 19801 4989 19857
rect 5045 19801 5131 19857
rect 5187 19801 5273 19857
rect 5329 19801 5415 19857
rect 5471 19801 5557 19857
rect 5613 19801 5699 19857
rect 5755 19801 5841 19857
rect 5897 19801 5983 19857
rect 6039 19801 6125 19857
rect 6181 19801 6267 19857
rect 6323 19801 6409 19857
rect 6465 19801 6551 19857
rect 6607 19801 6693 19857
rect 6749 19801 6835 19857
rect 6891 19801 6977 19857
rect 7033 19801 7119 19857
rect 7175 19801 7261 19857
rect 7317 19801 7403 19857
rect 7459 19801 7545 19857
rect 7601 19801 7687 19857
rect 7743 19801 7829 19857
rect 7885 19801 7971 19857
rect 8027 19801 8113 19857
rect 8169 19801 8255 19857
rect 8311 19801 8397 19857
rect 8453 19801 8539 19857
rect 8595 19801 8681 19857
rect 8737 19801 8823 19857
rect 8879 19801 8965 19857
rect 9021 19801 9107 19857
rect 9163 19801 9249 19857
rect 9305 19801 9391 19857
rect 9447 19801 9533 19857
rect 9589 19801 9675 19857
rect 9731 19801 9817 19857
rect 9873 19801 9959 19857
rect 10015 19801 10101 19857
rect 10157 19801 10243 19857
rect 10299 19801 10385 19857
rect 10441 19801 10527 19857
rect 10583 19801 10669 19857
rect 10725 19801 10811 19857
rect 10867 19801 10953 19857
rect 11009 19801 11095 19857
rect 11151 19801 11237 19857
rect 11293 19801 11379 19857
rect 11435 19801 11521 19857
rect 11577 19801 11663 19857
rect 11719 19801 11805 19857
rect 11861 19801 11947 19857
rect 12003 19801 12089 19857
rect 12145 19801 12231 19857
rect 12287 19801 12373 19857
rect 12429 19801 12515 19857
rect 12571 19801 12657 19857
rect 12713 19801 12799 19857
rect 12855 19801 12941 19857
rect 12997 19801 13083 19857
rect 13139 19801 13225 19857
rect 13281 19801 13367 19857
rect 13423 19801 13509 19857
rect 13565 19801 13651 19857
rect 13707 19801 13793 19857
rect 13849 19801 13935 19857
rect 13991 19801 14077 19857
rect 14133 19801 14219 19857
rect 14275 19801 14361 19857
rect 14417 19801 14503 19857
rect 14559 19801 14645 19857
rect 14701 19801 14787 19857
rect 14843 19801 14853 19857
rect 151 19715 14853 19801
rect 151 19659 161 19715
rect 217 19659 303 19715
rect 359 19659 445 19715
rect 501 19659 587 19715
rect 643 19659 729 19715
rect 785 19659 871 19715
rect 927 19659 1013 19715
rect 1069 19659 1155 19715
rect 1211 19659 1297 19715
rect 1353 19659 1439 19715
rect 1495 19659 1581 19715
rect 1637 19659 1723 19715
rect 1779 19659 1865 19715
rect 1921 19659 2007 19715
rect 2063 19659 2149 19715
rect 2205 19659 2291 19715
rect 2347 19659 2433 19715
rect 2489 19659 2575 19715
rect 2631 19659 2717 19715
rect 2773 19659 2859 19715
rect 2915 19659 3001 19715
rect 3057 19659 3143 19715
rect 3199 19659 3285 19715
rect 3341 19659 3427 19715
rect 3483 19659 3569 19715
rect 3625 19659 3711 19715
rect 3767 19659 3853 19715
rect 3909 19659 3995 19715
rect 4051 19659 4137 19715
rect 4193 19659 4279 19715
rect 4335 19659 4421 19715
rect 4477 19659 4563 19715
rect 4619 19659 4705 19715
rect 4761 19659 4847 19715
rect 4903 19659 4989 19715
rect 5045 19659 5131 19715
rect 5187 19659 5273 19715
rect 5329 19659 5415 19715
rect 5471 19659 5557 19715
rect 5613 19659 5699 19715
rect 5755 19659 5841 19715
rect 5897 19659 5983 19715
rect 6039 19659 6125 19715
rect 6181 19659 6267 19715
rect 6323 19659 6409 19715
rect 6465 19659 6551 19715
rect 6607 19659 6693 19715
rect 6749 19659 6835 19715
rect 6891 19659 6977 19715
rect 7033 19659 7119 19715
rect 7175 19659 7261 19715
rect 7317 19659 7403 19715
rect 7459 19659 7545 19715
rect 7601 19659 7687 19715
rect 7743 19659 7829 19715
rect 7885 19659 7971 19715
rect 8027 19659 8113 19715
rect 8169 19659 8255 19715
rect 8311 19659 8397 19715
rect 8453 19659 8539 19715
rect 8595 19659 8681 19715
rect 8737 19659 8823 19715
rect 8879 19659 8965 19715
rect 9021 19659 9107 19715
rect 9163 19659 9249 19715
rect 9305 19659 9391 19715
rect 9447 19659 9533 19715
rect 9589 19659 9675 19715
rect 9731 19659 9817 19715
rect 9873 19659 9959 19715
rect 10015 19659 10101 19715
rect 10157 19659 10243 19715
rect 10299 19659 10385 19715
rect 10441 19659 10527 19715
rect 10583 19659 10669 19715
rect 10725 19659 10811 19715
rect 10867 19659 10953 19715
rect 11009 19659 11095 19715
rect 11151 19659 11237 19715
rect 11293 19659 11379 19715
rect 11435 19659 11521 19715
rect 11577 19659 11663 19715
rect 11719 19659 11805 19715
rect 11861 19659 11947 19715
rect 12003 19659 12089 19715
rect 12145 19659 12231 19715
rect 12287 19659 12373 19715
rect 12429 19659 12515 19715
rect 12571 19659 12657 19715
rect 12713 19659 12799 19715
rect 12855 19659 12941 19715
rect 12997 19659 13083 19715
rect 13139 19659 13225 19715
rect 13281 19659 13367 19715
rect 13423 19659 13509 19715
rect 13565 19659 13651 19715
rect 13707 19659 13793 19715
rect 13849 19659 13935 19715
rect 13991 19659 14077 19715
rect 14133 19659 14219 19715
rect 14275 19659 14361 19715
rect 14417 19659 14503 19715
rect 14559 19659 14645 19715
rect 14701 19659 14787 19715
rect 14843 19659 14853 19715
rect 151 19573 14853 19659
rect 151 19517 161 19573
rect 217 19517 303 19573
rect 359 19517 445 19573
rect 501 19517 587 19573
rect 643 19517 729 19573
rect 785 19517 871 19573
rect 927 19517 1013 19573
rect 1069 19517 1155 19573
rect 1211 19517 1297 19573
rect 1353 19517 1439 19573
rect 1495 19517 1581 19573
rect 1637 19517 1723 19573
rect 1779 19517 1865 19573
rect 1921 19517 2007 19573
rect 2063 19517 2149 19573
rect 2205 19517 2291 19573
rect 2347 19517 2433 19573
rect 2489 19517 2575 19573
rect 2631 19517 2717 19573
rect 2773 19517 2859 19573
rect 2915 19517 3001 19573
rect 3057 19517 3143 19573
rect 3199 19517 3285 19573
rect 3341 19517 3427 19573
rect 3483 19517 3569 19573
rect 3625 19517 3711 19573
rect 3767 19517 3853 19573
rect 3909 19517 3995 19573
rect 4051 19517 4137 19573
rect 4193 19517 4279 19573
rect 4335 19517 4421 19573
rect 4477 19517 4563 19573
rect 4619 19517 4705 19573
rect 4761 19517 4847 19573
rect 4903 19517 4989 19573
rect 5045 19517 5131 19573
rect 5187 19517 5273 19573
rect 5329 19517 5415 19573
rect 5471 19517 5557 19573
rect 5613 19517 5699 19573
rect 5755 19517 5841 19573
rect 5897 19517 5983 19573
rect 6039 19517 6125 19573
rect 6181 19517 6267 19573
rect 6323 19517 6409 19573
rect 6465 19517 6551 19573
rect 6607 19517 6693 19573
rect 6749 19517 6835 19573
rect 6891 19517 6977 19573
rect 7033 19517 7119 19573
rect 7175 19517 7261 19573
rect 7317 19517 7403 19573
rect 7459 19517 7545 19573
rect 7601 19517 7687 19573
rect 7743 19517 7829 19573
rect 7885 19517 7971 19573
rect 8027 19517 8113 19573
rect 8169 19517 8255 19573
rect 8311 19517 8397 19573
rect 8453 19517 8539 19573
rect 8595 19517 8681 19573
rect 8737 19517 8823 19573
rect 8879 19517 8965 19573
rect 9021 19517 9107 19573
rect 9163 19517 9249 19573
rect 9305 19517 9391 19573
rect 9447 19517 9533 19573
rect 9589 19517 9675 19573
rect 9731 19517 9817 19573
rect 9873 19517 9959 19573
rect 10015 19517 10101 19573
rect 10157 19517 10243 19573
rect 10299 19517 10385 19573
rect 10441 19517 10527 19573
rect 10583 19517 10669 19573
rect 10725 19517 10811 19573
rect 10867 19517 10953 19573
rect 11009 19517 11095 19573
rect 11151 19517 11237 19573
rect 11293 19517 11379 19573
rect 11435 19517 11521 19573
rect 11577 19517 11663 19573
rect 11719 19517 11805 19573
rect 11861 19517 11947 19573
rect 12003 19517 12089 19573
rect 12145 19517 12231 19573
rect 12287 19517 12373 19573
rect 12429 19517 12515 19573
rect 12571 19517 12657 19573
rect 12713 19517 12799 19573
rect 12855 19517 12941 19573
rect 12997 19517 13083 19573
rect 13139 19517 13225 19573
rect 13281 19517 13367 19573
rect 13423 19517 13509 19573
rect 13565 19517 13651 19573
rect 13707 19517 13793 19573
rect 13849 19517 13935 19573
rect 13991 19517 14077 19573
rect 14133 19517 14219 19573
rect 14275 19517 14361 19573
rect 14417 19517 14503 19573
rect 14559 19517 14645 19573
rect 14701 19517 14787 19573
rect 14843 19517 14853 19573
rect 151 19431 14853 19517
rect 151 19375 161 19431
rect 217 19375 303 19431
rect 359 19375 445 19431
rect 501 19375 587 19431
rect 643 19375 729 19431
rect 785 19375 871 19431
rect 927 19375 1013 19431
rect 1069 19375 1155 19431
rect 1211 19375 1297 19431
rect 1353 19375 1439 19431
rect 1495 19375 1581 19431
rect 1637 19375 1723 19431
rect 1779 19375 1865 19431
rect 1921 19375 2007 19431
rect 2063 19375 2149 19431
rect 2205 19375 2291 19431
rect 2347 19375 2433 19431
rect 2489 19375 2575 19431
rect 2631 19375 2717 19431
rect 2773 19375 2859 19431
rect 2915 19375 3001 19431
rect 3057 19375 3143 19431
rect 3199 19375 3285 19431
rect 3341 19375 3427 19431
rect 3483 19375 3569 19431
rect 3625 19375 3711 19431
rect 3767 19375 3853 19431
rect 3909 19375 3995 19431
rect 4051 19375 4137 19431
rect 4193 19375 4279 19431
rect 4335 19375 4421 19431
rect 4477 19375 4563 19431
rect 4619 19375 4705 19431
rect 4761 19375 4847 19431
rect 4903 19375 4989 19431
rect 5045 19375 5131 19431
rect 5187 19375 5273 19431
rect 5329 19375 5415 19431
rect 5471 19375 5557 19431
rect 5613 19375 5699 19431
rect 5755 19375 5841 19431
rect 5897 19375 5983 19431
rect 6039 19375 6125 19431
rect 6181 19375 6267 19431
rect 6323 19375 6409 19431
rect 6465 19375 6551 19431
rect 6607 19375 6693 19431
rect 6749 19375 6835 19431
rect 6891 19375 6977 19431
rect 7033 19375 7119 19431
rect 7175 19375 7261 19431
rect 7317 19375 7403 19431
rect 7459 19375 7545 19431
rect 7601 19375 7687 19431
rect 7743 19375 7829 19431
rect 7885 19375 7971 19431
rect 8027 19375 8113 19431
rect 8169 19375 8255 19431
rect 8311 19375 8397 19431
rect 8453 19375 8539 19431
rect 8595 19375 8681 19431
rect 8737 19375 8823 19431
rect 8879 19375 8965 19431
rect 9021 19375 9107 19431
rect 9163 19375 9249 19431
rect 9305 19375 9391 19431
rect 9447 19375 9533 19431
rect 9589 19375 9675 19431
rect 9731 19375 9817 19431
rect 9873 19375 9959 19431
rect 10015 19375 10101 19431
rect 10157 19375 10243 19431
rect 10299 19375 10385 19431
rect 10441 19375 10527 19431
rect 10583 19375 10669 19431
rect 10725 19375 10811 19431
rect 10867 19375 10953 19431
rect 11009 19375 11095 19431
rect 11151 19375 11237 19431
rect 11293 19375 11379 19431
rect 11435 19375 11521 19431
rect 11577 19375 11663 19431
rect 11719 19375 11805 19431
rect 11861 19375 11947 19431
rect 12003 19375 12089 19431
rect 12145 19375 12231 19431
rect 12287 19375 12373 19431
rect 12429 19375 12515 19431
rect 12571 19375 12657 19431
rect 12713 19375 12799 19431
rect 12855 19375 12941 19431
rect 12997 19375 13083 19431
rect 13139 19375 13225 19431
rect 13281 19375 13367 19431
rect 13423 19375 13509 19431
rect 13565 19375 13651 19431
rect 13707 19375 13793 19431
rect 13849 19375 13935 19431
rect 13991 19375 14077 19431
rect 14133 19375 14219 19431
rect 14275 19375 14361 19431
rect 14417 19375 14503 19431
rect 14559 19375 14645 19431
rect 14701 19375 14787 19431
rect 14843 19375 14853 19431
rect 151 19289 14853 19375
rect 151 19233 161 19289
rect 217 19233 303 19289
rect 359 19233 445 19289
rect 501 19233 587 19289
rect 643 19233 729 19289
rect 785 19233 871 19289
rect 927 19233 1013 19289
rect 1069 19233 1155 19289
rect 1211 19233 1297 19289
rect 1353 19233 1439 19289
rect 1495 19233 1581 19289
rect 1637 19233 1723 19289
rect 1779 19233 1865 19289
rect 1921 19233 2007 19289
rect 2063 19233 2149 19289
rect 2205 19233 2291 19289
rect 2347 19233 2433 19289
rect 2489 19233 2575 19289
rect 2631 19233 2717 19289
rect 2773 19233 2859 19289
rect 2915 19233 3001 19289
rect 3057 19233 3143 19289
rect 3199 19233 3285 19289
rect 3341 19233 3427 19289
rect 3483 19233 3569 19289
rect 3625 19233 3711 19289
rect 3767 19233 3853 19289
rect 3909 19233 3995 19289
rect 4051 19233 4137 19289
rect 4193 19233 4279 19289
rect 4335 19233 4421 19289
rect 4477 19233 4563 19289
rect 4619 19233 4705 19289
rect 4761 19233 4847 19289
rect 4903 19233 4989 19289
rect 5045 19233 5131 19289
rect 5187 19233 5273 19289
rect 5329 19233 5415 19289
rect 5471 19233 5557 19289
rect 5613 19233 5699 19289
rect 5755 19233 5841 19289
rect 5897 19233 5983 19289
rect 6039 19233 6125 19289
rect 6181 19233 6267 19289
rect 6323 19233 6409 19289
rect 6465 19233 6551 19289
rect 6607 19233 6693 19289
rect 6749 19233 6835 19289
rect 6891 19233 6977 19289
rect 7033 19233 7119 19289
rect 7175 19233 7261 19289
rect 7317 19233 7403 19289
rect 7459 19233 7545 19289
rect 7601 19233 7687 19289
rect 7743 19233 7829 19289
rect 7885 19233 7971 19289
rect 8027 19233 8113 19289
rect 8169 19233 8255 19289
rect 8311 19233 8397 19289
rect 8453 19233 8539 19289
rect 8595 19233 8681 19289
rect 8737 19233 8823 19289
rect 8879 19233 8965 19289
rect 9021 19233 9107 19289
rect 9163 19233 9249 19289
rect 9305 19233 9391 19289
rect 9447 19233 9533 19289
rect 9589 19233 9675 19289
rect 9731 19233 9817 19289
rect 9873 19233 9959 19289
rect 10015 19233 10101 19289
rect 10157 19233 10243 19289
rect 10299 19233 10385 19289
rect 10441 19233 10527 19289
rect 10583 19233 10669 19289
rect 10725 19233 10811 19289
rect 10867 19233 10953 19289
rect 11009 19233 11095 19289
rect 11151 19233 11237 19289
rect 11293 19233 11379 19289
rect 11435 19233 11521 19289
rect 11577 19233 11663 19289
rect 11719 19233 11805 19289
rect 11861 19233 11947 19289
rect 12003 19233 12089 19289
rect 12145 19233 12231 19289
rect 12287 19233 12373 19289
rect 12429 19233 12515 19289
rect 12571 19233 12657 19289
rect 12713 19233 12799 19289
rect 12855 19233 12941 19289
rect 12997 19233 13083 19289
rect 13139 19233 13225 19289
rect 13281 19233 13367 19289
rect 13423 19233 13509 19289
rect 13565 19233 13651 19289
rect 13707 19233 13793 19289
rect 13849 19233 13935 19289
rect 13991 19233 14077 19289
rect 14133 19233 14219 19289
rect 14275 19233 14361 19289
rect 14417 19233 14503 19289
rect 14559 19233 14645 19289
rect 14701 19233 14787 19289
rect 14843 19233 14853 19289
rect 151 19147 14853 19233
rect 151 19091 161 19147
rect 217 19091 303 19147
rect 359 19091 445 19147
rect 501 19091 587 19147
rect 643 19091 729 19147
rect 785 19091 871 19147
rect 927 19091 1013 19147
rect 1069 19091 1155 19147
rect 1211 19091 1297 19147
rect 1353 19091 1439 19147
rect 1495 19091 1581 19147
rect 1637 19091 1723 19147
rect 1779 19091 1865 19147
rect 1921 19091 2007 19147
rect 2063 19091 2149 19147
rect 2205 19091 2291 19147
rect 2347 19091 2433 19147
rect 2489 19091 2575 19147
rect 2631 19091 2717 19147
rect 2773 19091 2859 19147
rect 2915 19091 3001 19147
rect 3057 19091 3143 19147
rect 3199 19091 3285 19147
rect 3341 19091 3427 19147
rect 3483 19091 3569 19147
rect 3625 19091 3711 19147
rect 3767 19091 3853 19147
rect 3909 19091 3995 19147
rect 4051 19091 4137 19147
rect 4193 19091 4279 19147
rect 4335 19091 4421 19147
rect 4477 19091 4563 19147
rect 4619 19091 4705 19147
rect 4761 19091 4847 19147
rect 4903 19091 4989 19147
rect 5045 19091 5131 19147
rect 5187 19091 5273 19147
rect 5329 19091 5415 19147
rect 5471 19091 5557 19147
rect 5613 19091 5699 19147
rect 5755 19091 5841 19147
rect 5897 19091 5983 19147
rect 6039 19091 6125 19147
rect 6181 19091 6267 19147
rect 6323 19091 6409 19147
rect 6465 19091 6551 19147
rect 6607 19091 6693 19147
rect 6749 19091 6835 19147
rect 6891 19091 6977 19147
rect 7033 19091 7119 19147
rect 7175 19091 7261 19147
rect 7317 19091 7403 19147
rect 7459 19091 7545 19147
rect 7601 19091 7687 19147
rect 7743 19091 7829 19147
rect 7885 19091 7971 19147
rect 8027 19091 8113 19147
rect 8169 19091 8255 19147
rect 8311 19091 8397 19147
rect 8453 19091 8539 19147
rect 8595 19091 8681 19147
rect 8737 19091 8823 19147
rect 8879 19091 8965 19147
rect 9021 19091 9107 19147
rect 9163 19091 9249 19147
rect 9305 19091 9391 19147
rect 9447 19091 9533 19147
rect 9589 19091 9675 19147
rect 9731 19091 9817 19147
rect 9873 19091 9959 19147
rect 10015 19091 10101 19147
rect 10157 19091 10243 19147
rect 10299 19091 10385 19147
rect 10441 19091 10527 19147
rect 10583 19091 10669 19147
rect 10725 19091 10811 19147
rect 10867 19091 10953 19147
rect 11009 19091 11095 19147
rect 11151 19091 11237 19147
rect 11293 19091 11379 19147
rect 11435 19091 11521 19147
rect 11577 19091 11663 19147
rect 11719 19091 11805 19147
rect 11861 19091 11947 19147
rect 12003 19091 12089 19147
rect 12145 19091 12231 19147
rect 12287 19091 12373 19147
rect 12429 19091 12515 19147
rect 12571 19091 12657 19147
rect 12713 19091 12799 19147
rect 12855 19091 12941 19147
rect 12997 19091 13083 19147
rect 13139 19091 13225 19147
rect 13281 19091 13367 19147
rect 13423 19091 13509 19147
rect 13565 19091 13651 19147
rect 13707 19091 13793 19147
rect 13849 19091 13935 19147
rect 13991 19091 14077 19147
rect 14133 19091 14219 19147
rect 14275 19091 14361 19147
rect 14417 19091 14503 19147
rect 14559 19091 14645 19147
rect 14701 19091 14787 19147
rect 14843 19091 14853 19147
rect 151 19005 14853 19091
rect 151 18949 161 19005
rect 217 18949 303 19005
rect 359 18949 445 19005
rect 501 18949 587 19005
rect 643 18949 729 19005
rect 785 18949 871 19005
rect 927 18949 1013 19005
rect 1069 18949 1155 19005
rect 1211 18949 1297 19005
rect 1353 18949 1439 19005
rect 1495 18949 1581 19005
rect 1637 18949 1723 19005
rect 1779 18949 1865 19005
rect 1921 18949 2007 19005
rect 2063 18949 2149 19005
rect 2205 18949 2291 19005
rect 2347 18949 2433 19005
rect 2489 18949 2575 19005
rect 2631 18949 2717 19005
rect 2773 18949 2859 19005
rect 2915 18949 3001 19005
rect 3057 18949 3143 19005
rect 3199 18949 3285 19005
rect 3341 18949 3427 19005
rect 3483 18949 3569 19005
rect 3625 18949 3711 19005
rect 3767 18949 3853 19005
rect 3909 18949 3995 19005
rect 4051 18949 4137 19005
rect 4193 18949 4279 19005
rect 4335 18949 4421 19005
rect 4477 18949 4563 19005
rect 4619 18949 4705 19005
rect 4761 18949 4847 19005
rect 4903 18949 4989 19005
rect 5045 18949 5131 19005
rect 5187 18949 5273 19005
rect 5329 18949 5415 19005
rect 5471 18949 5557 19005
rect 5613 18949 5699 19005
rect 5755 18949 5841 19005
rect 5897 18949 5983 19005
rect 6039 18949 6125 19005
rect 6181 18949 6267 19005
rect 6323 18949 6409 19005
rect 6465 18949 6551 19005
rect 6607 18949 6693 19005
rect 6749 18949 6835 19005
rect 6891 18949 6977 19005
rect 7033 18949 7119 19005
rect 7175 18949 7261 19005
rect 7317 18949 7403 19005
rect 7459 18949 7545 19005
rect 7601 18949 7687 19005
rect 7743 18949 7829 19005
rect 7885 18949 7971 19005
rect 8027 18949 8113 19005
rect 8169 18949 8255 19005
rect 8311 18949 8397 19005
rect 8453 18949 8539 19005
rect 8595 18949 8681 19005
rect 8737 18949 8823 19005
rect 8879 18949 8965 19005
rect 9021 18949 9107 19005
rect 9163 18949 9249 19005
rect 9305 18949 9391 19005
rect 9447 18949 9533 19005
rect 9589 18949 9675 19005
rect 9731 18949 9817 19005
rect 9873 18949 9959 19005
rect 10015 18949 10101 19005
rect 10157 18949 10243 19005
rect 10299 18949 10385 19005
rect 10441 18949 10527 19005
rect 10583 18949 10669 19005
rect 10725 18949 10811 19005
rect 10867 18949 10953 19005
rect 11009 18949 11095 19005
rect 11151 18949 11237 19005
rect 11293 18949 11379 19005
rect 11435 18949 11521 19005
rect 11577 18949 11663 19005
rect 11719 18949 11805 19005
rect 11861 18949 11947 19005
rect 12003 18949 12089 19005
rect 12145 18949 12231 19005
rect 12287 18949 12373 19005
rect 12429 18949 12515 19005
rect 12571 18949 12657 19005
rect 12713 18949 12799 19005
rect 12855 18949 12941 19005
rect 12997 18949 13083 19005
rect 13139 18949 13225 19005
rect 13281 18949 13367 19005
rect 13423 18949 13509 19005
rect 13565 18949 13651 19005
rect 13707 18949 13793 19005
rect 13849 18949 13935 19005
rect 13991 18949 14077 19005
rect 14133 18949 14219 19005
rect 14275 18949 14361 19005
rect 14417 18949 14503 19005
rect 14559 18949 14645 19005
rect 14701 18949 14787 19005
rect 14843 18949 14853 19005
rect 151 18863 14853 18949
rect 151 18807 161 18863
rect 217 18807 303 18863
rect 359 18807 445 18863
rect 501 18807 587 18863
rect 643 18807 729 18863
rect 785 18807 871 18863
rect 927 18807 1013 18863
rect 1069 18807 1155 18863
rect 1211 18807 1297 18863
rect 1353 18807 1439 18863
rect 1495 18807 1581 18863
rect 1637 18807 1723 18863
rect 1779 18807 1865 18863
rect 1921 18807 2007 18863
rect 2063 18807 2149 18863
rect 2205 18807 2291 18863
rect 2347 18807 2433 18863
rect 2489 18807 2575 18863
rect 2631 18807 2717 18863
rect 2773 18807 2859 18863
rect 2915 18807 3001 18863
rect 3057 18807 3143 18863
rect 3199 18807 3285 18863
rect 3341 18807 3427 18863
rect 3483 18807 3569 18863
rect 3625 18807 3711 18863
rect 3767 18807 3853 18863
rect 3909 18807 3995 18863
rect 4051 18807 4137 18863
rect 4193 18807 4279 18863
rect 4335 18807 4421 18863
rect 4477 18807 4563 18863
rect 4619 18807 4705 18863
rect 4761 18807 4847 18863
rect 4903 18807 4989 18863
rect 5045 18807 5131 18863
rect 5187 18807 5273 18863
rect 5329 18807 5415 18863
rect 5471 18807 5557 18863
rect 5613 18807 5699 18863
rect 5755 18807 5841 18863
rect 5897 18807 5983 18863
rect 6039 18807 6125 18863
rect 6181 18807 6267 18863
rect 6323 18807 6409 18863
rect 6465 18807 6551 18863
rect 6607 18807 6693 18863
rect 6749 18807 6835 18863
rect 6891 18807 6977 18863
rect 7033 18807 7119 18863
rect 7175 18807 7261 18863
rect 7317 18807 7403 18863
rect 7459 18807 7545 18863
rect 7601 18807 7687 18863
rect 7743 18807 7829 18863
rect 7885 18807 7971 18863
rect 8027 18807 8113 18863
rect 8169 18807 8255 18863
rect 8311 18807 8397 18863
rect 8453 18807 8539 18863
rect 8595 18807 8681 18863
rect 8737 18807 8823 18863
rect 8879 18807 8965 18863
rect 9021 18807 9107 18863
rect 9163 18807 9249 18863
rect 9305 18807 9391 18863
rect 9447 18807 9533 18863
rect 9589 18807 9675 18863
rect 9731 18807 9817 18863
rect 9873 18807 9959 18863
rect 10015 18807 10101 18863
rect 10157 18807 10243 18863
rect 10299 18807 10385 18863
rect 10441 18807 10527 18863
rect 10583 18807 10669 18863
rect 10725 18807 10811 18863
rect 10867 18807 10953 18863
rect 11009 18807 11095 18863
rect 11151 18807 11237 18863
rect 11293 18807 11379 18863
rect 11435 18807 11521 18863
rect 11577 18807 11663 18863
rect 11719 18807 11805 18863
rect 11861 18807 11947 18863
rect 12003 18807 12089 18863
rect 12145 18807 12231 18863
rect 12287 18807 12373 18863
rect 12429 18807 12515 18863
rect 12571 18807 12657 18863
rect 12713 18807 12799 18863
rect 12855 18807 12941 18863
rect 12997 18807 13083 18863
rect 13139 18807 13225 18863
rect 13281 18807 13367 18863
rect 13423 18807 13509 18863
rect 13565 18807 13651 18863
rect 13707 18807 13793 18863
rect 13849 18807 13935 18863
rect 13991 18807 14077 18863
rect 14133 18807 14219 18863
rect 14275 18807 14361 18863
rect 14417 18807 14503 18863
rect 14559 18807 14645 18863
rect 14701 18807 14787 18863
rect 14843 18807 14853 18863
rect 151 18721 14853 18807
rect 151 18665 161 18721
rect 217 18665 303 18721
rect 359 18665 445 18721
rect 501 18665 587 18721
rect 643 18665 729 18721
rect 785 18665 871 18721
rect 927 18665 1013 18721
rect 1069 18665 1155 18721
rect 1211 18665 1297 18721
rect 1353 18665 1439 18721
rect 1495 18665 1581 18721
rect 1637 18665 1723 18721
rect 1779 18665 1865 18721
rect 1921 18665 2007 18721
rect 2063 18665 2149 18721
rect 2205 18665 2291 18721
rect 2347 18665 2433 18721
rect 2489 18665 2575 18721
rect 2631 18665 2717 18721
rect 2773 18665 2859 18721
rect 2915 18665 3001 18721
rect 3057 18665 3143 18721
rect 3199 18665 3285 18721
rect 3341 18665 3427 18721
rect 3483 18665 3569 18721
rect 3625 18665 3711 18721
rect 3767 18665 3853 18721
rect 3909 18665 3995 18721
rect 4051 18665 4137 18721
rect 4193 18665 4279 18721
rect 4335 18665 4421 18721
rect 4477 18665 4563 18721
rect 4619 18665 4705 18721
rect 4761 18665 4847 18721
rect 4903 18665 4989 18721
rect 5045 18665 5131 18721
rect 5187 18665 5273 18721
rect 5329 18665 5415 18721
rect 5471 18665 5557 18721
rect 5613 18665 5699 18721
rect 5755 18665 5841 18721
rect 5897 18665 5983 18721
rect 6039 18665 6125 18721
rect 6181 18665 6267 18721
rect 6323 18665 6409 18721
rect 6465 18665 6551 18721
rect 6607 18665 6693 18721
rect 6749 18665 6835 18721
rect 6891 18665 6977 18721
rect 7033 18665 7119 18721
rect 7175 18665 7261 18721
rect 7317 18665 7403 18721
rect 7459 18665 7545 18721
rect 7601 18665 7687 18721
rect 7743 18665 7829 18721
rect 7885 18665 7971 18721
rect 8027 18665 8113 18721
rect 8169 18665 8255 18721
rect 8311 18665 8397 18721
rect 8453 18665 8539 18721
rect 8595 18665 8681 18721
rect 8737 18665 8823 18721
rect 8879 18665 8965 18721
rect 9021 18665 9107 18721
rect 9163 18665 9249 18721
rect 9305 18665 9391 18721
rect 9447 18665 9533 18721
rect 9589 18665 9675 18721
rect 9731 18665 9817 18721
rect 9873 18665 9959 18721
rect 10015 18665 10101 18721
rect 10157 18665 10243 18721
rect 10299 18665 10385 18721
rect 10441 18665 10527 18721
rect 10583 18665 10669 18721
rect 10725 18665 10811 18721
rect 10867 18665 10953 18721
rect 11009 18665 11095 18721
rect 11151 18665 11237 18721
rect 11293 18665 11379 18721
rect 11435 18665 11521 18721
rect 11577 18665 11663 18721
rect 11719 18665 11805 18721
rect 11861 18665 11947 18721
rect 12003 18665 12089 18721
rect 12145 18665 12231 18721
rect 12287 18665 12373 18721
rect 12429 18665 12515 18721
rect 12571 18665 12657 18721
rect 12713 18665 12799 18721
rect 12855 18665 12941 18721
rect 12997 18665 13083 18721
rect 13139 18665 13225 18721
rect 13281 18665 13367 18721
rect 13423 18665 13509 18721
rect 13565 18665 13651 18721
rect 13707 18665 13793 18721
rect 13849 18665 13935 18721
rect 13991 18665 14077 18721
rect 14133 18665 14219 18721
rect 14275 18665 14361 18721
rect 14417 18665 14503 18721
rect 14559 18665 14645 18721
rect 14701 18665 14787 18721
rect 14843 18665 14853 18721
rect 151 18579 14853 18665
rect 151 18523 161 18579
rect 217 18523 303 18579
rect 359 18523 445 18579
rect 501 18523 587 18579
rect 643 18523 729 18579
rect 785 18523 871 18579
rect 927 18523 1013 18579
rect 1069 18523 1155 18579
rect 1211 18523 1297 18579
rect 1353 18523 1439 18579
rect 1495 18523 1581 18579
rect 1637 18523 1723 18579
rect 1779 18523 1865 18579
rect 1921 18523 2007 18579
rect 2063 18523 2149 18579
rect 2205 18523 2291 18579
rect 2347 18523 2433 18579
rect 2489 18523 2575 18579
rect 2631 18523 2717 18579
rect 2773 18523 2859 18579
rect 2915 18523 3001 18579
rect 3057 18523 3143 18579
rect 3199 18523 3285 18579
rect 3341 18523 3427 18579
rect 3483 18523 3569 18579
rect 3625 18523 3711 18579
rect 3767 18523 3853 18579
rect 3909 18523 3995 18579
rect 4051 18523 4137 18579
rect 4193 18523 4279 18579
rect 4335 18523 4421 18579
rect 4477 18523 4563 18579
rect 4619 18523 4705 18579
rect 4761 18523 4847 18579
rect 4903 18523 4989 18579
rect 5045 18523 5131 18579
rect 5187 18523 5273 18579
rect 5329 18523 5415 18579
rect 5471 18523 5557 18579
rect 5613 18523 5699 18579
rect 5755 18523 5841 18579
rect 5897 18523 5983 18579
rect 6039 18523 6125 18579
rect 6181 18523 6267 18579
rect 6323 18523 6409 18579
rect 6465 18523 6551 18579
rect 6607 18523 6693 18579
rect 6749 18523 6835 18579
rect 6891 18523 6977 18579
rect 7033 18523 7119 18579
rect 7175 18523 7261 18579
rect 7317 18523 7403 18579
rect 7459 18523 7545 18579
rect 7601 18523 7687 18579
rect 7743 18523 7829 18579
rect 7885 18523 7971 18579
rect 8027 18523 8113 18579
rect 8169 18523 8255 18579
rect 8311 18523 8397 18579
rect 8453 18523 8539 18579
rect 8595 18523 8681 18579
rect 8737 18523 8823 18579
rect 8879 18523 8965 18579
rect 9021 18523 9107 18579
rect 9163 18523 9249 18579
rect 9305 18523 9391 18579
rect 9447 18523 9533 18579
rect 9589 18523 9675 18579
rect 9731 18523 9817 18579
rect 9873 18523 9959 18579
rect 10015 18523 10101 18579
rect 10157 18523 10243 18579
rect 10299 18523 10385 18579
rect 10441 18523 10527 18579
rect 10583 18523 10669 18579
rect 10725 18523 10811 18579
rect 10867 18523 10953 18579
rect 11009 18523 11095 18579
rect 11151 18523 11237 18579
rect 11293 18523 11379 18579
rect 11435 18523 11521 18579
rect 11577 18523 11663 18579
rect 11719 18523 11805 18579
rect 11861 18523 11947 18579
rect 12003 18523 12089 18579
rect 12145 18523 12231 18579
rect 12287 18523 12373 18579
rect 12429 18523 12515 18579
rect 12571 18523 12657 18579
rect 12713 18523 12799 18579
rect 12855 18523 12941 18579
rect 12997 18523 13083 18579
rect 13139 18523 13225 18579
rect 13281 18523 13367 18579
rect 13423 18523 13509 18579
rect 13565 18523 13651 18579
rect 13707 18523 13793 18579
rect 13849 18523 13935 18579
rect 13991 18523 14077 18579
rect 14133 18523 14219 18579
rect 14275 18523 14361 18579
rect 14417 18523 14503 18579
rect 14559 18523 14645 18579
rect 14701 18523 14787 18579
rect 14843 18523 14853 18579
rect 151 18437 14853 18523
rect 151 18381 161 18437
rect 217 18381 303 18437
rect 359 18381 445 18437
rect 501 18381 587 18437
rect 643 18381 729 18437
rect 785 18381 871 18437
rect 927 18381 1013 18437
rect 1069 18381 1155 18437
rect 1211 18381 1297 18437
rect 1353 18381 1439 18437
rect 1495 18381 1581 18437
rect 1637 18381 1723 18437
rect 1779 18381 1865 18437
rect 1921 18381 2007 18437
rect 2063 18381 2149 18437
rect 2205 18381 2291 18437
rect 2347 18381 2433 18437
rect 2489 18381 2575 18437
rect 2631 18381 2717 18437
rect 2773 18381 2859 18437
rect 2915 18381 3001 18437
rect 3057 18381 3143 18437
rect 3199 18381 3285 18437
rect 3341 18381 3427 18437
rect 3483 18381 3569 18437
rect 3625 18381 3711 18437
rect 3767 18381 3853 18437
rect 3909 18381 3995 18437
rect 4051 18381 4137 18437
rect 4193 18381 4279 18437
rect 4335 18381 4421 18437
rect 4477 18381 4563 18437
rect 4619 18381 4705 18437
rect 4761 18381 4847 18437
rect 4903 18381 4989 18437
rect 5045 18381 5131 18437
rect 5187 18381 5273 18437
rect 5329 18381 5415 18437
rect 5471 18381 5557 18437
rect 5613 18381 5699 18437
rect 5755 18381 5841 18437
rect 5897 18381 5983 18437
rect 6039 18381 6125 18437
rect 6181 18381 6267 18437
rect 6323 18381 6409 18437
rect 6465 18381 6551 18437
rect 6607 18381 6693 18437
rect 6749 18381 6835 18437
rect 6891 18381 6977 18437
rect 7033 18381 7119 18437
rect 7175 18381 7261 18437
rect 7317 18381 7403 18437
rect 7459 18381 7545 18437
rect 7601 18381 7687 18437
rect 7743 18381 7829 18437
rect 7885 18381 7971 18437
rect 8027 18381 8113 18437
rect 8169 18381 8255 18437
rect 8311 18381 8397 18437
rect 8453 18381 8539 18437
rect 8595 18381 8681 18437
rect 8737 18381 8823 18437
rect 8879 18381 8965 18437
rect 9021 18381 9107 18437
rect 9163 18381 9249 18437
rect 9305 18381 9391 18437
rect 9447 18381 9533 18437
rect 9589 18381 9675 18437
rect 9731 18381 9817 18437
rect 9873 18381 9959 18437
rect 10015 18381 10101 18437
rect 10157 18381 10243 18437
rect 10299 18381 10385 18437
rect 10441 18381 10527 18437
rect 10583 18381 10669 18437
rect 10725 18381 10811 18437
rect 10867 18381 10953 18437
rect 11009 18381 11095 18437
rect 11151 18381 11237 18437
rect 11293 18381 11379 18437
rect 11435 18381 11521 18437
rect 11577 18381 11663 18437
rect 11719 18381 11805 18437
rect 11861 18381 11947 18437
rect 12003 18381 12089 18437
rect 12145 18381 12231 18437
rect 12287 18381 12373 18437
rect 12429 18381 12515 18437
rect 12571 18381 12657 18437
rect 12713 18381 12799 18437
rect 12855 18381 12941 18437
rect 12997 18381 13083 18437
rect 13139 18381 13225 18437
rect 13281 18381 13367 18437
rect 13423 18381 13509 18437
rect 13565 18381 13651 18437
rect 13707 18381 13793 18437
rect 13849 18381 13935 18437
rect 13991 18381 14077 18437
rect 14133 18381 14219 18437
rect 14275 18381 14361 18437
rect 14417 18381 14503 18437
rect 14559 18381 14645 18437
rect 14701 18381 14787 18437
rect 14843 18381 14853 18437
rect 151 18295 14853 18381
rect 151 18239 161 18295
rect 217 18239 303 18295
rect 359 18239 445 18295
rect 501 18239 587 18295
rect 643 18239 729 18295
rect 785 18239 871 18295
rect 927 18239 1013 18295
rect 1069 18239 1155 18295
rect 1211 18239 1297 18295
rect 1353 18239 1439 18295
rect 1495 18239 1581 18295
rect 1637 18239 1723 18295
rect 1779 18239 1865 18295
rect 1921 18239 2007 18295
rect 2063 18239 2149 18295
rect 2205 18239 2291 18295
rect 2347 18239 2433 18295
rect 2489 18239 2575 18295
rect 2631 18239 2717 18295
rect 2773 18239 2859 18295
rect 2915 18239 3001 18295
rect 3057 18239 3143 18295
rect 3199 18239 3285 18295
rect 3341 18239 3427 18295
rect 3483 18239 3569 18295
rect 3625 18239 3711 18295
rect 3767 18239 3853 18295
rect 3909 18239 3995 18295
rect 4051 18239 4137 18295
rect 4193 18239 4279 18295
rect 4335 18239 4421 18295
rect 4477 18239 4563 18295
rect 4619 18239 4705 18295
rect 4761 18239 4847 18295
rect 4903 18239 4989 18295
rect 5045 18239 5131 18295
rect 5187 18239 5273 18295
rect 5329 18239 5415 18295
rect 5471 18239 5557 18295
rect 5613 18239 5699 18295
rect 5755 18239 5841 18295
rect 5897 18239 5983 18295
rect 6039 18239 6125 18295
rect 6181 18239 6267 18295
rect 6323 18239 6409 18295
rect 6465 18239 6551 18295
rect 6607 18239 6693 18295
rect 6749 18239 6835 18295
rect 6891 18239 6977 18295
rect 7033 18239 7119 18295
rect 7175 18239 7261 18295
rect 7317 18239 7403 18295
rect 7459 18239 7545 18295
rect 7601 18239 7687 18295
rect 7743 18239 7829 18295
rect 7885 18239 7971 18295
rect 8027 18239 8113 18295
rect 8169 18239 8255 18295
rect 8311 18239 8397 18295
rect 8453 18239 8539 18295
rect 8595 18239 8681 18295
rect 8737 18239 8823 18295
rect 8879 18239 8965 18295
rect 9021 18239 9107 18295
rect 9163 18239 9249 18295
rect 9305 18239 9391 18295
rect 9447 18239 9533 18295
rect 9589 18239 9675 18295
rect 9731 18239 9817 18295
rect 9873 18239 9959 18295
rect 10015 18239 10101 18295
rect 10157 18239 10243 18295
rect 10299 18239 10385 18295
rect 10441 18239 10527 18295
rect 10583 18239 10669 18295
rect 10725 18239 10811 18295
rect 10867 18239 10953 18295
rect 11009 18239 11095 18295
rect 11151 18239 11237 18295
rect 11293 18239 11379 18295
rect 11435 18239 11521 18295
rect 11577 18239 11663 18295
rect 11719 18239 11805 18295
rect 11861 18239 11947 18295
rect 12003 18239 12089 18295
rect 12145 18239 12231 18295
rect 12287 18239 12373 18295
rect 12429 18239 12515 18295
rect 12571 18239 12657 18295
rect 12713 18239 12799 18295
rect 12855 18239 12941 18295
rect 12997 18239 13083 18295
rect 13139 18239 13225 18295
rect 13281 18239 13367 18295
rect 13423 18239 13509 18295
rect 13565 18239 13651 18295
rect 13707 18239 13793 18295
rect 13849 18239 13935 18295
rect 13991 18239 14077 18295
rect 14133 18239 14219 18295
rect 14275 18239 14361 18295
rect 14417 18239 14503 18295
rect 14559 18239 14645 18295
rect 14701 18239 14787 18295
rect 14843 18239 14853 18295
rect 151 18153 14853 18239
rect 151 18097 161 18153
rect 217 18097 303 18153
rect 359 18097 445 18153
rect 501 18097 587 18153
rect 643 18097 729 18153
rect 785 18097 871 18153
rect 927 18097 1013 18153
rect 1069 18097 1155 18153
rect 1211 18097 1297 18153
rect 1353 18097 1439 18153
rect 1495 18097 1581 18153
rect 1637 18097 1723 18153
rect 1779 18097 1865 18153
rect 1921 18097 2007 18153
rect 2063 18097 2149 18153
rect 2205 18097 2291 18153
rect 2347 18097 2433 18153
rect 2489 18097 2575 18153
rect 2631 18097 2717 18153
rect 2773 18097 2859 18153
rect 2915 18097 3001 18153
rect 3057 18097 3143 18153
rect 3199 18097 3285 18153
rect 3341 18097 3427 18153
rect 3483 18097 3569 18153
rect 3625 18097 3711 18153
rect 3767 18097 3853 18153
rect 3909 18097 3995 18153
rect 4051 18097 4137 18153
rect 4193 18097 4279 18153
rect 4335 18097 4421 18153
rect 4477 18097 4563 18153
rect 4619 18097 4705 18153
rect 4761 18097 4847 18153
rect 4903 18097 4989 18153
rect 5045 18097 5131 18153
rect 5187 18097 5273 18153
rect 5329 18097 5415 18153
rect 5471 18097 5557 18153
rect 5613 18097 5699 18153
rect 5755 18097 5841 18153
rect 5897 18097 5983 18153
rect 6039 18097 6125 18153
rect 6181 18097 6267 18153
rect 6323 18097 6409 18153
rect 6465 18097 6551 18153
rect 6607 18097 6693 18153
rect 6749 18097 6835 18153
rect 6891 18097 6977 18153
rect 7033 18097 7119 18153
rect 7175 18097 7261 18153
rect 7317 18097 7403 18153
rect 7459 18097 7545 18153
rect 7601 18097 7687 18153
rect 7743 18097 7829 18153
rect 7885 18097 7971 18153
rect 8027 18097 8113 18153
rect 8169 18097 8255 18153
rect 8311 18097 8397 18153
rect 8453 18097 8539 18153
rect 8595 18097 8681 18153
rect 8737 18097 8823 18153
rect 8879 18097 8965 18153
rect 9021 18097 9107 18153
rect 9163 18097 9249 18153
rect 9305 18097 9391 18153
rect 9447 18097 9533 18153
rect 9589 18097 9675 18153
rect 9731 18097 9817 18153
rect 9873 18097 9959 18153
rect 10015 18097 10101 18153
rect 10157 18097 10243 18153
rect 10299 18097 10385 18153
rect 10441 18097 10527 18153
rect 10583 18097 10669 18153
rect 10725 18097 10811 18153
rect 10867 18097 10953 18153
rect 11009 18097 11095 18153
rect 11151 18097 11237 18153
rect 11293 18097 11379 18153
rect 11435 18097 11521 18153
rect 11577 18097 11663 18153
rect 11719 18097 11805 18153
rect 11861 18097 11947 18153
rect 12003 18097 12089 18153
rect 12145 18097 12231 18153
rect 12287 18097 12373 18153
rect 12429 18097 12515 18153
rect 12571 18097 12657 18153
rect 12713 18097 12799 18153
rect 12855 18097 12941 18153
rect 12997 18097 13083 18153
rect 13139 18097 13225 18153
rect 13281 18097 13367 18153
rect 13423 18097 13509 18153
rect 13565 18097 13651 18153
rect 13707 18097 13793 18153
rect 13849 18097 13935 18153
rect 13991 18097 14077 18153
rect 14133 18097 14219 18153
rect 14275 18097 14361 18153
rect 14417 18097 14503 18153
rect 14559 18097 14645 18153
rect 14701 18097 14787 18153
rect 14843 18097 14853 18153
rect 151 18011 14853 18097
rect 151 17955 161 18011
rect 217 17955 303 18011
rect 359 17955 445 18011
rect 501 17955 587 18011
rect 643 17955 729 18011
rect 785 17955 871 18011
rect 927 17955 1013 18011
rect 1069 17955 1155 18011
rect 1211 17955 1297 18011
rect 1353 17955 1439 18011
rect 1495 17955 1581 18011
rect 1637 17955 1723 18011
rect 1779 17955 1865 18011
rect 1921 17955 2007 18011
rect 2063 17955 2149 18011
rect 2205 17955 2291 18011
rect 2347 17955 2433 18011
rect 2489 17955 2575 18011
rect 2631 17955 2717 18011
rect 2773 17955 2859 18011
rect 2915 17955 3001 18011
rect 3057 17955 3143 18011
rect 3199 17955 3285 18011
rect 3341 17955 3427 18011
rect 3483 17955 3569 18011
rect 3625 17955 3711 18011
rect 3767 17955 3853 18011
rect 3909 17955 3995 18011
rect 4051 17955 4137 18011
rect 4193 17955 4279 18011
rect 4335 17955 4421 18011
rect 4477 17955 4563 18011
rect 4619 17955 4705 18011
rect 4761 17955 4847 18011
rect 4903 17955 4989 18011
rect 5045 17955 5131 18011
rect 5187 17955 5273 18011
rect 5329 17955 5415 18011
rect 5471 17955 5557 18011
rect 5613 17955 5699 18011
rect 5755 17955 5841 18011
rect 5897 17955 5983 18011
rect 6039 17955 6125 18011
rect 6181 17955 6267 18011
rect 6323 17955 6409 18011
rect 6465 17955 6551 18011
rect 6607 17955 6693 18011
rect 6749 17955 6835 18011
rect 6891 17955 6977 18011
rect 7033 17955 7119 18011
rect 7175 17955 7261 18011
rect 7317 17955 7403 18011
rect 7459 17955 7545 18011
rect 7601 17955 7687 18011
rect 7743 17955 7829 18011
rect 7885 17955 7971 18011
rect 8027 17955 8113 18011
rect 8169 17955 8255 18011
rect 8311 17955 8397 18011
rect 8453 17955 8539 18011
rect 8595 17955 8681 18011
rect 8737 17955 8823 18011
rect 8879 17955 8965 18011
rect 9021 17955 9107 18011
rect 9163 17955 9249 18011
rect 9305 17955 9391 18011
rect 9447 17955 9533 18011
rect 9589 17955 9675 18011
rect 9731 17955 9817 18011
rect 9873 17955 9959 18011
rect 10015 17955 10101 18011
rect 10157 17955 10243 18011
rect 10299 17955 10385 18011
rect 10441 17955 10527 18011
rect 10583 17955 10669 18011
rect 10725 17955 10811 18011
rect 10867 17955 10953 18011
rect 11009 17955 11095 18011
rect 11151 17955 11237 18011
rect 11293 17955 11379 18011
rect 11435 17955 11521 18011
rect 11577 17955 11663 18011
rect 11719 17955 11805 18011
rect 11861 17955 11947 18011
rect 12003 17955 12089 18011
rect 12145 17955 12231 18011
rect 12287 17955 12373 18011
rect 12429 17955 12515 18011
rect 12571 17955 12657 18011
rect 12713 17955 12799 18011
rect 12855 17955 12941 18011
rect 12997 17955 13083 18011
rect 13139 17955 13225 18011
rect 13281 17955 13367 18011
rect 13423 17955 13509 18011
rect 13565 17955 13651 18011
rect 13707 17955 13793 18011
rect 13849 17955 13935 18011
rect 13991 17955 14077 18011
rect 14133 17955 14219 18011
rect 14275 17955 14361 18011
rect 14417 17955 14503 18011
rect 14559 17955 14645 18011
rect 14701 17955 14787 18011
rect 14843 17955 14853 18011
rect 151 17869 14853 17955
rect 151 17813 161 17869
rect 217 17813 303 17869
rect 359 17813 445 17869
rect 501 17813 587 17869
rect 643 17813 729 17869
rect 785 17813 871 17869
rect 927 17813 1013 17869
rect 1069 17813 1155 17869
rect 1211 17813 1297 17869
rect 1353 17813 1439 17869
rect 1495 17813 1581 17869
rect 1637 17813 1723 17869
rect 1779 17813 1865 17869
rect 1921 17813 2007 17869
rect 2063 17813 2149 17869
rect 2205 17813 2291 17869
rect 2347 17813 2433 17869
rect 2489 17813 2575 17869
rect 2631 17813 2717 17869
rect 2773 17813 2859 17869
rect 2915 17813 3001 17869
rect 3057 17813 3143 17869
rect 3199 17813 3285 17869
rect 3341 17813 3427 17869
rect 3483 17813 3569 17869
rect 3625 17813 3711 17869
rect 3767 17813 3853 17869
rect 3909 17813 3995 17869
rect 4051 17813 4137 17869
rect 4193 17813 4279 17869
rect 4335 17813 4421 17869
rect 4477 17813 4563 17869
rect 4619 17813 4705 17869
rect 4761 17813 4847 17869
rect 4903 17813 4989 17869
rect 5045 17813 5131 17869
rect 5187 17813 5273 17869
rect 5329 17813 5415 17869
rect 5471 17813 5557 17869
rect 5613 17813 5699 17869
rect 5755 17813 5841 17869
rect 5897 17813 5983 17869
rect 6039 17813 6125 17869
rect 6181 17813 6267 17869
rect 6323 17813 6409 17869
rect 6465 17813 6551 17869
rect 6607 17813 6693 17869
rect 6749 17813 6835 17869
rect 6891 17813 6977 17869
rect 7033 17813 7119 17869
rect 7175 17813 7261 17869
rect 7317 17813 7403 17869
rect 7459 17813 7545 17869
rect 7601 17813 7687 17869
rect 7743 17813 7829 17869
rect 7885 17813 7971 17869
rect 8027 17813 8113 17869
rect 8169 17813 8255 17869
rect 8311 17813 8397 17869
rect 8453 17813 8539 17869
rect 8595 17813 8681 17869
rect 8737 17813 8823 17869
rect 8879 17813 8965 17869
rect 9021 17813 9107 17869
rect 9163 17813 9249 17869
rect 9305 17813 9391 17869
rect 9447 17813 9533 17869
rect 9589 17813 9675 17869
rect 9731 17813 9817 17869
rect 9873 17813 9959 17869
rect 10015 17813 10101 17869
rect 10157 17813 10243 17869
rect 10299 17813 10385 17869
rect 10441 17813 10527 17869
rect 10583 17813 10669 17869
rect 10725 17813 10811 17869
rect 10867 17813 10953 17869
rect 11009 17813 11095 17869
rect 11151 17813 11237 17869
rect 11293 17813 11379 17869
rect 11435 17813 11521 17869
rect 11577 17813 11663 17869
rect 11719 17813 11805 17869
rect 11861 17813 11947 17869
rect 12003 17813 12089 17869
rect 12145 17813 12231 17869
rect 12287 17813 12373 17869
rect 12429 17813 12515 17869
rect 12571 17813 12657 17869
rect 12713 17813 12799 17869
rect 12855 17813 12941 17869
rect 12997 17813 13083 17869
rect 13139 17813 13225 17869
rect 13281 17813 13367 17869
rect 13423 17813 13509 17869
rect 13565 17813 13651 17869
rect 13707 17813 13793 17869
rect 13849 17813 13935 17869
rect 13991 17813 14077 17869
rect 14133 17813 14219 17869
rect 14275 17813 14361 17869
rect 14417 17813 14503 17869
rect 14559 17813 14645 17869
rect 14701 17813 14787 17869
rect 14843 17813 14853 17869
rect 151 17727 14853 17813
rect 151 17671 161 17727
rect 217 17671 303 17727
rect 359 17671 445 17727
rect 501 17671 587 17727
rect 643 17671 729 17727
rect 785 17671 871 17727
rect 927 17671 1013 17727
rect 1069 17671 1155 17727
rect 1211 17671 1297 17727
rect 1353 17671 1439 17727
rect 1495 17671 1581 17727
rect 1637 17671 1723 17727
rect 1779 17671 1865 17727
rect 1921 17671 2007 17727
rect 2063 17671 2149 17727
rect 2205 17671 2291 17727
rect 2347 17671 2433 17727
rect 2489 17671 2575 17727
rect 2631 17671 2717 17727
rect 2773 17671 2859 17727
rect 2915 17671 3001 17727
rect 3057 17671 3143 17727
rect 3199 17671 3285 17727
rect 3341 17671 3427 17727
rect 3483 17671 3569 17727
rect 3625 17671 3711 17727
rect 3767 17671 3853 17727
rect 3909 17671 3995 17727
rect 4051 17671 4137 17727
rect 4193 17671 4279 17727
rect 4335 17671 4421 17727
rect 4477 17671 4563 17727
rect 4619 17671 4705 17727
rect 4761 17671 4847 17727
rect 4903 17671 4989 17727
rect 5045 17671 5131 17727
rect 5187 17671 5273 17727
rect 5329 17671 5415 17727
rect 5471 17671 5557 17727
rect 5613 17671 5699 17727
rect 5755 17671 5841 17727
rect 5897 17671 5983 17727
rect 6039 17671 6125 17727
rect 6181 17671 6267 17727
rect 6323 17671 6409 17727
rect 6465 17671 6551 17727
rect 6607 17671 6693 17727
rect 6749 17671 6835 17727
rect 6891 17671 6977 17727
rect 7033 17671 7119 17727
rect 7175 17671 7261 17727
rect 7317 17671 7403 17727
rect 7459 17671 7545 17727
rect 7601 17671 7687 17727
rect 7743 17671 7829 17727
rect 7885 17671 7971 17727
rect 8027 17671 8113 17727
rect 8169 17671 8255 17727
rect 8311 17671 8397 17727
rect 8453 17671 8539 17727
rect 8595 17671 8681 17727
rect 8737 17671 8823 17727
rect 8879 17671 8965 17727
rect 9021 17671 9107 17727
rect 9163 17671 9249 17727
rect 9305 17671 9391 17727
rect 9447 17671 9533 17727
rect 9589 17671 9675 17727
rect 9731 17671 9817 17727
rect 9873 17671 9959 17727
rect 10015 17671 10101 17727
rect 10157 17671 10243 17727
rect 10299 17671 10385 17727
rect 10441 17671 10527 17727
rect 10583 17671 10669 17727
rect 10725 17671 10811 17727
rect 10867 17671 10953 17727
rect 11009 17671 11095 17727
rect 11151 17671 11237 17727
rect 11293 17671 11379 17727
rect 11435 17671 11521 17727
rect 11577 17671 11663 17727
rect 11719 17671 11805 17727
rect 11861 17671 11947 17727
rect 12003 17671 12089 17727
rect 12145 17671 12231 17727
rect 12287 17671 12373 17727
rect 12429 17671 12515 17727
rect 12571 17671 12657 17727
rect 12713 17671 12799 17727
rect 12855 17671 12941 17727
rect 12997 17671 13083 17727
rect 13139 17671 13225 17727
rect 13281 17671 13367 17727
rect 13423 17671 13509 17727
rect 13565 17671 13651 17727
rect 13707 17671 13793 17727
rect 13849 17671 13935 17727
rect 13991 17671 14077 17727
rect 14133 17671 14219 17727
rect 14275 17671 14361 17727
rect 14417 17671 14503 17727
rect 14559 17671 14645 17727
rect 14701 17671 14787 17727
rect 14843 17671 14853 17727
rect 151 17585 14853 17671
rect 151 17529 161 17585
rect 217 17529 303 17585
rect 359 17529 445 17585
rect 501 17529 587 17585
rect 643 17529 729 17585
rect 785 17529 871 17585
rect 927 17529 1013 17585
rect 1069 17529 1155 17585
rect 1211 17529 1297 17585
rect 1353 17529 1439 17585
rect 1495 17529 1581 17585
rect 1637 17529 1723 17585
rect 1779 17529 1865 17585
rect 1921 17529 2007 17585
rect 2063 17529 2149 17585
rect 2205 17529 2291 17585
rect 2347 17529 2433 17585
rect 2489 17529 2575 17585
rect 2631 17529 2717 17585
rect 2773 17529 2859 17585
rect 2915 17529 3001 17585
rect 3057 17529 3143 17585
rect 3199 17529 3285 17585
rect 3341 17529 3427 17585
rect 3483 17529 3569 17585
rect 3625 17529 3711 17585
rect 3767 17529 3853 17585
rect 3909 17529 3995 17585
rect 4051 17529 4137 17585
rect 4193 17529 4279 17585
rect 4335 17529 4421 17585
rect 4477 17529 4563 17585
rect 4619 17529 4705 17585
rect 4761 17529 4847 17585
rect 4903 17529 4989 17585
rect 5045 17529 5131 17585
rect 5187 17529 5273 17585
rect 5329 17529 5415 17585
rect 5471 17529 5557 17585
rect 5613 17529 5699 17585
rect 5755 17529 5841 17585
rect 5897 17529 5983 17585
rect 6039 17529 6125 17585
rect 6181 17529 6267 17585
rect 6323 17529 6409 17585
rect 6465 17529 6551 17585
rect 6607 17529 6693 17585
rect 6749 17529 6835 17585
rect 6891 17529 6977 17585
rect 7033 17529 7119 17585
rect 7175 17529 7261 17585
rect 7317 17529 7403 17585
rect 7459 17529 7545 17585
rect 7601 17529 7687 17585
rect 7743 17529 7829 17585
rect 7885 17529 7971 17585
rect 8027 17529 8113 17585
rect 8169 17529 8255 17585
rect 8311 17529 8397 17585
rect 8453 17529 8539 17585
rect 8595 17529 8681 17585
rect 8737 17529 8823 17585
rect 8879 17529 8965 17585
rect 9021 17529 9107 17585
rect 9163 17529 9249 17585
rect 9305 17529 9391 17585
rect 9447 17529 9533 17585
rect 9589 17529 9675 17585
rect 9731 17529 9817 17585
rect 9873 17529 9959 17585
rect 10015 17529 10101 17585
rect 10157 17529 10243 17585
rect 10299 17529 10385 17585
rect 10441 17529 10527 17585
rect 10583 17529 10669 17585
rect 10725 17529 10811 17585
rect 10867 17529 10953 17585
rect 11009 17529 11095 17585
rect 11151 17529 11237 17585
rect 11293 17529 11379 17585
rect 11435 17529 11521 17585
rect 11577 17529 11663 17585
rect 11719 17529 11805 17585
rect 11861 17529 11947 17585
rect 12003 17529 12089 17585
rect 12145 17529 12231 17585
rect 12287 17529 12373 17585
rect 12429 17529 12515 17585
rect 12571 17529 12657 17585
rect 12713 17529 12799 17585
rect 12855 17529 12941 17585
rect 12997 17529 13083 17585
rect 13139 17529 13225 17585
rect 13281 17529 13367 17585
rect 13423 17529 13509 17585
rect 13565 17529 13651 17585
rect 13707 17529 13793 17585
rect 13849 17529 13935 17585
rect 13991 17529 14077 17585
rect 14133 17529 14219 17585
rect 14275 17529 14361 17585
rect 14417 17529 14503 17585
rect 14559 17529 14645 17585
rect 14701 17529 14787 17585
rect 14843 17529 14853 17585
rect 151 17443 14853 17529
rect 151 17387 161 17443
rect 217 17387 303 17443
rect 359 17387 445 17443
rect 501 17387 587 17443
rect 643 17387 729 17443
rect 785 17387 871 17443
rect 927 17387 1013 17443
rect 1069 17387 1155 17443
rect 1211 17387 1297 17443
rect 1353 17387 1439 17443
rect 1495 17387 1581 17443
rect 1637 17387 1723 17443
rect 1779 17387 1865 17443
rect 1921 17387 2007 17443
rect 2063 17387 2149 17443
rect 2205 17387 2291 17443
rect 2347 17387 2433 17443
rect 2489 17387 2575 17443
rect 2631 17387 2717 17443
rect 2773 17387 2859 17443
rect 2915 17387 3001 17443
rect 3057 17387 3143 17443
rect 3199 17387 3285 17443
rect 3341 17387 3427 17443
rect 3483 17387 3569 17443
rect 3625 17387 3711 17443
rect 3767 17387 3853 17443
rect 3909 17387 3995 17443
rect 4051 17387 4137 17443
rect 4193 17387 4279 17443
rect 4335 17387 4421 17443
rect 4477 17387 4563 17443
rect 4619 17387 4705 17443
rect 4761 17387 4847 17443
rect 4903 17387 4989 17443
rect 5045 17387 5131 17443
rect 5187 17387 5273 17443
rect 5329 17387 5415 17443
rect 5471 17387 5557 17443
rect 5613 17387 5699 17443
rect 5755 17387 5841 17443
rect 5897 17387 5983 17443
rect 6039 17387 6125 17443
rect 6181 17387 6267 17443
rect 6323 17387 6409 17443
rect 6465 17387 6551 17443
rect 6607 17387 6693 17443
rect 6749 17387 6835 17443
rect 6891 17387 6977 17443
rect 7033 17387 7119 17443
rect 7175 17387 7261 17443
rect 7317 17387 7403 17443
rect 7459 17387 7545 17443
rect 7601 17387 7687 17443
rect 7743 17387 7829 17443
rect 7885 17387 7971 17443
rect 8027 17387 8113 17443
rect 8169 17387 8255 17443
rect 8311 17387 8397 17443
rect 8453 17387 8539 17443
rect 8595 17387 8681 17443
rect 8737 17387 8823 17443
rect 8879 17387 8965 17443
rect 9021 17387 9107 17443
rect 9163 17387 9249 17443
rect 9305 17387 9391 17443
rect 9447 17387 9533 17443
rect 9589 17387 9675 17443
rect 9731 17387 9817 17443
rect 9873 17387 9959 17443
rect 10015 17387 10101 17443
rect 10157 17387 10243 17443
rect 10299 17387 10385 17443
rect 10441 17387 10527 17443
rect 10583 17387 10669 17443
rect 10725 17387 10811 17443
rect 10867 17387 10953 17443
rect 11009 17387 11095 17443
rect 11151 17387 11237 17443
rect 11293 17387 11379 17443
rect 11435 17387 11521 17443
rect 11577 17387 11663 17443
rect 11719 17387 11805 17443
rect 11861 17387 11947 17443
rect 12003 17387 12089 17443
rect 12145 17387 12231 17443
rect 12287 17387 12373 17443
rect 12429 17387 12515 17443
rect 12571 17387 12657 17443
rect 12713 17387 12799 17443
rect 12855 17387 12941 17443
rect 12997 17387 13083 17443
rect 13139 17387 13225 17443
rect 13281 17387 13367 17443
rect 13423 17387 13509 17443
rect 13565 17387 13651 17443
rect 13707 17387 13793 17443
rect 13849 17387 13935 17443
rect 13991 17387 14077 17443
rect 14133 17387 14219 17443
rect 14275 17387 14361 17443
rect 14417 17387 14503 17443
rect 14559 17387 14645 17443
rect 14701 17387 14787 17443
rect 14843 17387 14853 17443
rect 151 17301 14853 17387
rect 151 17245 161 17301
rect 217 17245 303 17301
rect 359 17245 445 17301
rect 501 17245 587 17301
rect 643 17245 729 17301
rect 785 17245 871 17301
rect 927 17245 1013 17301
rect 1069 17245 1155 17301
rect 1211 17245 1297 17301
rect 1353 17245 1439 17301
rect 1495 17245 1581 17301
rect 1637 17245 1723 17301
rect 1779 17245 1865 17301
rect 1921 17245 2007 17301
rect 2063 17245 2149 17301
rect 2205 17245 2291 17301
rect 2347 17245 2433 17301
rect 2489 17245 2575 17301
rect 2631 17245 2717 17301
rect 2773 17245 2859 17301
rect 2915 17245 3001 17301
rect 3057 17245 3143 17301
rect 3199 17245 3285 17301
rect 3341 17245 3427 17301
rect 3483 17245 3569 17301
rect 3625 17245 3711 17301
rect 3767 17245 3853 17301
rect 3909 17245 3995 17301
rect 4051 17245 4137 17301
rect 4193 17245 4279 17301
rect 4335 17245 4421 17301
rect 4477 17245 4563 17301
rect 4619 17245 4705 17301
rect 4761 17245 4847 17301
rect 4903 17245 4989 17301
rect 5045 17245 5131 17301
rect 5187 17245 5273 17301
rect 5329 17245 5415 17301
rect 5471 17245 5557 17301
rect 5613 17245 5699 17301
rect 5755 17245 5841 17301
rect 5897 17245 5983 17301
rect 6039 17245 6125 17301
rect 6181 17245 6267 17301
rect 6323 17245 6409 17301
rect 6465 17245 6551 17301
rect 6607 17245 6693 17301
rect 6749 17245 6835 17301
rect 6891 17245 6977 17301
rect 7033 17245 7119 17301
rect 7175 17245 7261 17301
rect 7317 17245 7403 17301
rect 7459 17245 7545 17301
rect 7601 17245 7687 17301
rect 7743 17245 7829 17301
rect 7885 17245 7971 17301
rect 8027 17245 8113 17301
rect 8169 17245 8255 17301
rect 8311 17245 8397 17301
rect 8453 17245 8539 17301
rect 8595 17245 8681 17301
rect 8737 17245 8823 17301
rect 8879 17245 8965 17301
rect 9021 17245 9107 17301
rect 9163 17245 9249 17301
rect 9305 17245 9391 17301
rect 9447 17245 9533 17301
rect 9589 17245 9675 17301
rect 9731 17245 9817 17301
rect 9873 17245 9959 17301
rect 10015 17245 10101 17301
rect 10157 17245 10243 17301
rect 10299 17245 10385 17301
rect 10441 17245 10527 17301
rect 10583 17245 10669 17301
rect 10725 17245 10811 17301
rect 10867 17245 10953 17301
rect 11009 17245 11095 17301
rect 11151 17245 11237 17301
rect 11293 17245 11379 17301
rect 11435 17245 11521 17301
rect 11577 17245 11663 17301
rect 11719 17245 11805 17301
rect 11861 17245 11947 17301
rect 12003 17245 12089 17301
rect 12145 17245 12231 17301
rect 12287 17245 12373 17301
rect 12429 17245 12515 17301
rect 12571 17245 12657 17301
rect 12713 17245 12799 17301
rect 12855 17245 12941 17301
rect 12997 17245 13083 17301
rect 13139 17245 13225 17301
rect 13281 17245 13367 17301
rect 13423 17245 13509 17301
rect 13565 17245 13651 17301
rect 13707 17245 13793 17301
rect 13849 17245 13935 17301
rect 13991 17245 14077 17301
rect 14133 17245 14219 17301
rect 14275 17245 14361 17301
rect 14417 17245 14503 17301
rect 14559 17245 14645 17301
rect 14701 17245 14787 17301
rect 14843 17245 14853 17301
rect 151 17235 14853 17245
rect 151 16941 14853 16951
rect 151 16885 161 16941
rect 217 16885 303 16941
rect 359 16885 445 16941
rect 501 16885 587 16941
rect 643 16885 729 16941
rect 785 16885 871 16941
rect 927 16885 1013 16941
rect 1069 16885 1155 16941
rect 1211 16885 1297 16941
rect 1353 16885 1439 16941
rect 1495 16885 1581 16941
rect 1637 16885 1723 16941
rect 1779 16885 1865 16941
rect 1921 16885 2007 16941
rect 2063 16885 2149 16941
rect 2205 16885 2291 16941
rect 2347 16885 2433 16941
rect 2489 16885 2575 16941
rect 2631 16885 2717 16941
rect 2773 16885 2859 16941
rect 2915 16885 3001 16941
rect 3057 16885 3143 16941
rect 3199 16885 3285 16941
rect 3341 16885 3427 16941
rect 3483 16885 3569 16941
rect 3625 16885 3711 16941
rect 3767 16885 3853 16941
rect 3909 16885 3995 16941
rect 4051 16885 4137 16941
rect 4193 16885 4279 16941
rect 4335 16885 4421 16941
rect 4477 16885 4563 16941
rect 4619 16885 4705 16941
rect 4761 16885 4847 16941
rect 4903 16885 4989 16941
rect 5045 16885 5131 16941
rect 5187 16885 5273 16941
rect 5329 16885 5415 16941
rect 5471 16885 5557 16941
rect 5613 16885 5699 16941
rect 5755 16885 5841 16941
rect 5897 16885 5983 16941
rect 6039 16885 6125 16941
rect 6181 16885 6267 16941
rect 6323 16885 6409 16941
rect 6465 16885 6551 16941
rect 6607 16885 6693 16941
rect 6749 16885 6835 16941
rect 6891 16885 6977 16941
rect 7033 16885 7119 16941
rect 7175 16885 7261 16941
rect 7317 16885 7403 16941
rect 7459 16885 7545 16941
rect 7601 16885 7687 16941
rect 7743 16885 7829 16941
rect 7885 16885 7971 16941
rect 8027 16885 8113 16941
rect 8169 16885 8255 16941
rect 8311 16885 8397 16941
rect 8453 16885 8539 16941
rect 8595 16885 8681 16941
rect 8737 16885 8823 16941
rect 8879 16885 8965 16941
rect 9021 16885 9107 16941
rect 9163 16885 9249 16941
rect 9305 16885 9391 16941
rect 9447 16885 9533 16941
rect 9589 16885 9675 16941
rect 9731 16885 9817 16941
rect 9873 16885 9959 16941
rect 10015 16885 10101 16941
rect 10157 16885 10243 16941
rect 10299 16885 10385 16941
rect 10441 16885 10527 16941
rect 10583 16885 10669 16941
rect 10725 16885 10811 16941
rect 10867 16885 10953 16941
rect 11009 16885 11095 16941
rect 11151 16885 11237 16941
rect 11293 16885 11379 16941
rect 11435 16885 11521 16941
rect 11577 16885 11663 16941
rect 11719 16885 11805 16941
rect 11861 16885 11947 16941
rect 12003 16885 12089 16941
rect 12145 16885 12231 16941
rect 12287 16885 12373 16941
rect 12429 16885 12515 16941
rect 12571 16885 12657 16941
rect 12713 16885 12799 16941
rect 12855 16885 12941 16941
rect 12997 16885 13083 16941
rect 13139 16885 13225 16941
rect 13281 16885 13367 16941
rect 13423 16885 13509 16941
rect 13565 16885 13651 16941
rect 13707 16885 13793 16941
rect 13849 16885 13935 16941
rect 13991 16885 14077 16941
rect 14133 16885 14219 16941
rect 14275 16885 14361 16941
rect 14417 16885 14503 16941
rect 14559 16885 14645 16941
rect 14701 16885 14787 16941
rect 14843 16885 14853 16941
rect 151 16799 14853 16885
rect 151 16743 161 16799
rect 217 16743 303 16799
rect 359 16743 445 16799
rect 501 16743 587 16799
rect 643 16743 729 16799
rect 785 16743 871 16799
rect 927 16743 1013 16799
rect 1069 16743 1155 16799
rect 1211 16743 1297 16799
rect 1353 16743 1439 16799
rect 1495 16743 1581 16799
rect 1637 16743 1723 16799
rect 1779 16743 1865 16799
rect 1921 16743 2007 16799
rect 2063 16743 2149 16799
rect 2205 16743 2291 16799
rect 2347 16743 2433 16799
rect 2489 16743 2575 16799
rect 2631 16743 2717 16799
rect 2773 16743 2859 16799
rect 2915 16743 3001 16799
rect 3057 16743 3143 16799
rect 3199 16743 3285 16799
rect 3341 16743 3427 16799
rect 3483 16743 3569 16799
rect 3625 16743 3711 16799
rect 3767 16743 3853 16799
rect 3909 16743 3995 16799
rect 4051 16743 4137 16799
rect 4193 16743 4279 16799
rect 4335 16743 4421 16799
rect 4477 16743 4563 16799
rect 4619 16743 4705 16799
rect 4761 16743 4847 16799
rect 4903 16743 4989 16799
rect 5045 16743 5131 16799
rect 5187 16743 5273 16799
rect 5329 16743 5415 16799
rect 5471 16743 5557 16799
rect 5613 16743 5699 16799
rect 5755 16743 5841 16799
rect 5897 16743 5983 16799
rect 6039 16743 6125 16799
rect 6181 16743 6267 16799
rect 6323 16743 6409 16799
rect 6465 16743 6551 16799
rect 6607 16743 6693 16799
rect 6749 16743 6835 16799
rect 6891 16743 6977 16799
rect 7033 16743 7119 16799
rect 7175 16743 7261 16799
rect 7317 16743 7403 16799
rect 7459 16743 7545 16799
rect 7601 16743 7687 16799
rect 7743 16743 7829 16799
rect 7885 16743 7971 16799
rect 8027 16743 8113 16799
rect 8169 16743 8255 16799
rect 8311 16743 8397 16799
rect 8453 16743 8539 16799
rect 8595 16743 8681 16799
rect 8737 16743 8823 16799
rect 8879 16743 8965 16799
rect 9021 16743 9107 16799
rect 9163 16743 9249 16799
rect 9305 16743 9391 16799
rect 9447 16743 9533 16799
rect 9589 16743 9675 16799
rect 9731 16743 9817 16799
rect 9873 16743 9959 16799
rect 10015 16743 10101 16799
rect 10157 16743 10243 16799
rect 10299 16743 10385 16799
rect 10441 16743 10527 16799
rect 10583 16743 10669 16799
rect 10725 16743 10811 16799
rect 10867 16743 10953 16799
rect 11009 16743 11095 16799
rect 11151 16743 11237 16799
rect 11293 16743 11379 16799
rect 11435 16743 11521 16799
rect 11577 16743 11663 16799
rect 11719 16743 11805 16799
rect 11861 16743 11947 16799
rect 12003 16743 12089 16799
rect 12145 16743 12231 16799
rect 12287 16743 12373 16799
rect 12429 16743 12515 16799
rect 12571 16743 12657 16799
rect 12713 16743 12799 16799
rect 12855 16743 12941 16799
rect 12997 16743 13083 16799
rect 13139 16743 13225 16799
rect 13281 16743 13367 16799
rect 13423 16743 13509 16799
rect 13565 16743 13651 16799
rect 13707 16743 13793 16799
rect 13849 16743 13935 16799
rect 13991 16743 14077 16799
rect 14133 16743 14219 16799
rect 14275 16743 14361 16799
rect 14417 16743 14503 16799
rect 14559 16743 14645 16799
rect 14701 16743 14787 16799
rect 14843 16743 14853 16799
rect 151 16657 14853 16743
rect 151 16601 161 16657
rect 217 16601 303 16657
rect 359 16601 445 16657
rect 501 16601 587 16657
rect 643 16601 729 16657
rect 785 16601 871 16657
rect 927 16601 1013 16657
rect 1069 16601 1155 16657
rect 1211 16601 1297 16657
rect 1353 16601 1439 16657
rect 1495 16601 1581 16657
rect 1637 16601 1723 16657
rect 1779 16601 1865 16657
rect 1921 16601 2007 16657
rect 2063 16601 2149 16657
rect 2205 16601 2291 16657
rect 2347 16601 2433 16657
rect 2489 16601 2575 16657
rect 2631 16601 2717 16657
rect 2773 16601 2859 16657
rect 2915 16601 3001 16657
rect 3057 16601 3143 16657
rect 3199 16601 3285 16657
rect 3341 16601 3427 16657
rect 3483 16601 3569 16657
rect 3625 16601 3711 16657
rect 3767 16601 3853 16657
rect 3909 16601 3995 16657
rect 4051 16601 4137 16657
rect 4193 16601 4279 16657
rect 4335 16601 4421 16657
rect 4477 16601 4563 16657
rect 4619 16601 4705 16657
rect 4761 16601 4847 16657
rect 4903 16601 4989 16657
rect 5045 16601 5131 16657
rect 5187 16601 5273 16657
rect 5329 16601 5415 16657
rect 5471 16601 5557 16657
rect 5613 16601 5699 16657
rect 5755 16601 5841 16657
rect 5897 16601 5983 16657
rect 6039 16601 6125 16657
rect 6181 16601 6267 16657
rect 6323 16601 6409 16657
rect 6465 16601 6551 16657
rect 6607 16601 6693 16657
rect 6749 16601 6835 16657
rect 6891 16601 6977 16657
rect 7033 16601 7119 16657
rect 7175 16601 7261 16657
rect 7317 16601 7403 16657
rect 7459 16601 7545 16657
rect 7601 16601 7687 16657
rect 7743 16601 7829 16657
rect 7885 16601 7971 16657
rect 8027 16601 8113 16657
rect 8169 16601 8255 16657
rect 8311 16601 8397 16657
rect 8453 16601 8539 16657
rect 8595 16601 8681 16657
rect 8737 16601 8823 16657
rect 8879 16601 8965 16657
rect 9021 16601 9107 16657
rect 9163 16601 9249 16657
rect 9305 16601 9391 16657
rect 9447 16601 9533 16657
rect 9589 16601 9675 16657
rect 9731 16601 9817 16657
rect 9873 16601 9959 16657
rect 10015 16601 10101 16657
rect 10157 16601 10243 16657
rect 10299 16601 10385 16657
rect 10441 16601 10527 16657
rect 10583 16601 10669 16657
rect 10725 16601 10811 16657
rect 10867 16601 10953 16657
rect 11009 16601 11095 16657
rect 11151 16601 11237 16657
rect 11293 16601 11379 16657
rect 11435 16601 11521 16657
rect 11577 16601 11663 16657
rect 11719 16601 11805 16657
rect 11861 16601 11947 16657
rect 12003 16601 12089 16657
rect 12145 16601 12231 16657
rect 12287 16601 12373 16657
rect 12429 16601 12515 16657
rect 12571 16601 12657 16657
rect 12713 16601 12799 16657
rect 12855 16601 12941 16657
rect 12997 16601 13083 16657
rect 13139 16601 13225 16657
rect 13281 16601 13367 16657
rect 13423 16601 13509 16657
rect 13565 16601 13651 16657
rect 13707 16601 13793 16657
rect 13849 16601 13935 16657
rect 13991 16601 14077 16657
rect 14133 16601 14219 16657
rect 14275 16601 14361 16657
rect 14417 16601 14503 16657
rect 14559 16601 14645 16657
rect 14701 16601 14787 16657
rect 14843 16601 14853 16657
rect 151 16515 14853 16601
rect 151 16459 161 16515
rect 217 16459 303 16515
rect 359 16459 445 16515
rect 501 16459 587 16515
rect 643 16459 729 16515
rect 785 16459 871 16515
rect 927 16459 1013 16515
rect 1069 16459 1155 16515
rect 1211 16459 1297 16515
rect 1353 16459 1439 16515
rect 1495 16459 1581 16515
rect 1637 16459 1723 16515
rect 1779 16459 1865 16515
rect 1921 16459 2007 16515
rect 2063 16459 2149 16515
rect 2205 16459 2291 16515
rect 2347 16459 2433 16515
rect 2489 16459 2575 16515
rect 2631 16459 2717 16515
rect 2773 16459 2859 16515
rect 2915 16459 3001 16515
rect 3057 16459 3143 16515
rect 3199 16459 3285 16515
rect 3341 16459 3427 16515
rect 3483 16459 3569 16515
rect 3625 16459 3711 16515
rect 3767 16459 3853 16515
rect 3909 16459 3995 16515
rect 4051 16459 4137 16515
rect 4193 16459 4279 16515
rect 4335 16459 4421 16515
rect 4477 16459 4563 16515
rect 4619 16459 4705 16515
rect 4761 16459 4847 16515
rect 4903 16459 4989 16515
rect 5045 16459 5131 16515
rect 5187 16459 5273 16515
rect 5329 16459 5415 16515
rect 5471 16459 5557 16515
rect 5613 16459 5699 16515
rect 5755 16459 5841 16515
rect 5897 16459 5983 16515
rect 6039 16459 6125 16515
rect 6181 16459 6267 16515
rect 6323 16459 6409 16515
rect 6465 16459 6551 16515
rect 6607 16459 6693 16515
rect 6749 16459 6835 16515
rect 6891 16459 6977 16515
rect 7033 16459 7119 16515
rect 7175 16459 7261 16515
rect 7317 16459 7403 16515
rect 7459 16459 7545 16515
rect 7601 16459 7687 16515
rect 7743 16459 7829 16515
rect 7885 16459 7971 16515
rect 8027 16459 8113 16515
rect 8169 16459 8255 16515
rect 8311 16459 8397 16515
rect 8453 16459 8539 16515
rect 8595 16459 8681 16515
rect 8737 16459 8823 16515
rect 8879 16459 8965 16515
rect 9021 16459 9107 16515
rect 9163 16459 9249 16515
rect 9305 16459 9391 16515
rect 9447 16459 9533 16515
rect 9589 16459 9675 16515
rect 9731 16459 9817 16515
rect 9873 16459 9959 16515
rect 10015 16459 10101 16515
rect 10157 16459 10243 16515
rect 10299 16459 10385 16515
rect 10441 16459 10527 16515
rect 10583 16459 10669 16515
rect 10725 16459 10811 16515
rect 10867 16459 10953 16515
rect 11009 16459 11095 16515
rect 11151 16459 11237 16515
rect 11293 16459 11379 16515
rect 11435 16459 11521 16515
rect 11577 16459 11663 16515
rect 11719 16459 11805 16515
rect 11861 16459 11947 16515
rect 12003 16459 12089 16515
rect 12145 16459 12231 16515
rect 12287 16459 12373 16515
rect 12429 16459 12515 16515
rect 12571 16459 12657 16515
rect 12713 16459 12799 16515
rect 12855 16459 12941 16515
rect 12997 16459 13083 16515
rect 13139 16459 13225 16515
rect 13281 16459 13367 16515
rect 13423 16459 13509 16515
rect 13565 16459 13651 16515
rect 13707 16459 13793 16515
rect 13849 16459 13935 16515
rect 13991 16459 14077 16515
rect 14133 16459 14219 16515
rect 14275 16459 14361 16515
rect 14417 16459 14503 16515
rect 14559 16459 14645 16515
rect 14701 16459 14787 16515
rect 14843 16459 14853 16515
rect 151 16373 14853 16459
rect 151 16317 161 16373
rect 217 16317 303 16373
rect 359 16317 445 16373
rect 501 16317 587 16373
rect 643 16317 729 16373
rect 785 16317 871 16373
rect 927 16317 1013 16373
rect 1069 16317 1155 16373
rect 1211 16317 1297 16373
rect 1353 16317 1439 16373
rect 1495 16317 1581 16373
rect 1637 16317 1723 16373
rect 1779 16317 1865 16373
rect 1921 16317 2007 16373
rect 2063 16317 2149 16373
rect 2205 16317 2291 16373
rect 2347 16317 2433 16373
rect 2489 16317 2575 16373
rect 2631 16317 2717 16373
rect 2773 16317 2859 16373
rect 2915 16317 3001 16373
rect 3057 16317 3143 16373
rect 3199 16317 3285 16373
rect 3341 16317 3427 16373
rect 3483 16317 3569 16373
rect 3625 16317 3711 16373
rect 3767 16317 3853 16373
rect 3909 16317 3995 16373
rect 4051 16317 4137 16373
rect 4193 16317 4279 16373
rect 4335 16317 4421 16373
rect 4477 16317 4563 16373
rect 4619 16317 4705 16373
rect 4761 16317 4847 16373
rect 4903 16317 4989 16373
rect 5045 16317 5131 16373
rect 5187 16317 5273 16373
rect 5329 16317 5415 16373
rect 5471 16317 5557 16373
rect 5613 16317 5699 16373
rect 5755 16317 5841 16373
rect 5897 16317 5983 16373
rect 6039 16317 6125 16373
rect 6181 16317 6267 16373
rect 6323 16317 6409 16373
rect 6465 16317 6551 16373
rect 6607 16317 6693 16373
rect 6749 16317 6835 16373
rect 6891 16317 6977 16373
rect 7033 16317 7119 16373
rect 7175 16317 7261 16373
rect 7317 16317 7403 16373
rect 7459 16317 7545 16373
rect 7601 16317 7687 16373
rect 7743 16317 7829 16373
rect 7885 16317 7971 16373
rect 8027 16317 8113 16373
rect 8169 16317 8255 16373
rect 8311 16317 8397 16373
rect 8453 16317 8539 16373
rect 8595 16317 8681 16373
rect 8737 16317 8823 16373
rect 8879 16317 8965 16373
rect 9021 16317 9107 16373
rect 9163 16317 9249 16373
rect 9305 16317 9391 16373
rect 9447 16317 9533 16373
rect 9589 16317 9675 16373
rect 9731 16317 9817 16373
rect 9873 16317 9959 16373
rect 10015 16317 10101 16373
rect 10157 16317 10243 16373
rect 10299 16317 10385 16373
rect 10441 16317 10527 16373
rect 10583 16317 10669 16373
rect 10725 16317 10811 16373
rect 10867 16317 10953 16373
rect 11009 16317 11095 16373
rect 11151 16317 11237 16373
rect 11293 16317 11379 16373
rect 11435 16317 11521 16373
rect 11577 16317 11663 16373
rect 11719 16317 11805 16373
rect 11861 16317 11947 16373
rect 12003 16317 12089 16373
rect 12145 16317 12231 16373
rect 12287 16317 12373 16373
rect 12429 16317 12515 16373
rect 12571 16317 12657 16373
rect 12713 16317 12799 16373
rect 12855 16317 12941 16373
rect 12997 16317 13083 16373
rect 13139 16317 13225 16373
rect 13281 16317 13367 16373
rect 13423 16317 13509 16373
rect 13565 16317 13651 16373
rect 13707 16317 13793 16373
rect 13849 16317 13935 16373
rect 13991 16317 14077 16373
rect 14133 16317 14219 16373
rect 14275 16317 14361 16373
rect 14417 16317 14503 16373
rect 14559 16317 14645 16373
rect 14701 16317 14787 16373
rect 14843 16317 14853 16373
rect 151 16231 14853 16317
rect 151 16175 161 16231
rect 217 16175 303 16231
rect 359 16175 445 16231
rect 501 16175 587 16231
rect 643 16175 729 16231
rect 785 16175 871 16231
rect 927 16175 1013 16231
rect 1069 16175 1155 16231
rect 1211 16175 1297 16231
rect 1353 16175 1439 16231
rect 1495 16175 1581 16231
rect 1637 16175 1723 16231
rect 1779 16175 1865 16231
rect 1921 16175 2007 16231
rect 2063 16175 2149 16231
rect 2205 16175 2291 16231
rect 2347 16175 2433 16231
rect 2489 16175 2575 16231
rect 2631 16175 2717 16231
rect 2773 16175 2859 16231
rect 2915 16175 3001 16231
rect 3057 16175 3143 16231
rect 3199 16175 3285 16231
rect 3341 16175 3427 16231
rect 3483 16175 3569 16231
rect 3625 16175 3711 16231
rect 3767 16175 3853 16231
rect 3909 16175 3995 16231
rect 4051 16175 4137 16231
rect 4193 16175 4279 16231
rect 4335 16175 4421 16231
rect 4477 16175 4563 16231
rect 4619 16175 4705 16231
rect 4761 16175 4847 16231
rect 4903 16175 4989 16231
rect 5045 16175 5131 16231
rect 5187 16175 5273 16231
rect 5329 16175 5415 16231
rect 5471 16175 5557 16231
rect 5613 16175 5699 16231
rect 5755 16175 5841 16231
rect 5897 16175 5983 16231
rect 6039 16175 6125 16231
rect 6181 16175 6267 16231
rect 6323 16175 6409 16231
rect 6465 16175 6551 16231
rect 6607 16175 6693 16231
rect 6749 16175 6835 16231
rect 6891 16175 6977 16231
rect 7033 16175 7119 16231
rect 7175 16175 7261 16231
rect 7317 16175 7403 16231
rect 7459 16175 7545 16231
rect 7601 16175 7687 16231
rect 7743 16175 7829 16231
rect 7885 16175 7971 16231
rect 8027 16175 8113 16231
rect 8169 16175 8255 16231
rect 8311 16175 8397 16231
rect 8453 16175 8539 16231
rect 8595 16175 8681 16231
rect 8737 16175 8823 16231
rect 8879 16175 8965 16231
rect 9021 16175 9107 16231
rect 9163 16175 9249 16231
rect 9305 16175 9391 16231
rect 9447 16175 9533 16231
rect 9589 16175 9675 16231
rect 9731 16175 9817 16231
rect 9873 16175 9959 16231
rect 10015 16175 10101 16231
rect 10157 16175 10243 16231
rect 10299 16175 10385 16231
rect 10441 16175 10527 16231
rect 10583 16175 10669 16231
rect 10725 16175 10811 16231
rect 10867 16175 10953 16231
rect 11009 16175 11095 16231
rect 11151 16175 11237 16231
rect 11293 16175 11379 16231
rect 11435 16175 11521 16231
rect 11577 16175 11663 16231
rect 11719 16175 11805 16231
rect 11861 16175 11947 16231
rect 12003 16175 12089 16231
rect 12145 16175 12231 16231
rect 12287 16175 12373 16231
rect 12429 16175 12515 16231
rect 12571 16175 12657 16231
rect 12713 16175 12799 16231
rect 12855 16175 12941 16231
rect 12997 16175 13083 16231
rect 13139 16175 13225 16231
rect 13281 16175 13367 16231
rect 13423 16175 13509 16231
rect 13565 16175 13651 16231
rect 13707 16175 13793 16231
rect 13849 16175 13935 16231
rect 13991 16175 14077 16231
rect 14133 16175 14219 16231
rect 14275 16175 14361 16231
rect 14417 16175 14503 16231
rect 14559 16175 14645 16231
rect 14701 16175 14787 16231
rect 14843 16175 14853 16231
rect 151 16089 14853 16175
rect 151 16033 161 16089
rect 217 16033 303 16089
rect 359 16033 445 16089
rect 501 16033 587 16089
rect 643 16033 729 16089
rect 785 16033 871 16089
rect 927 16033 1013 16089
rect 1069 16033 1155 16089
rect 1211 16033 1297 16089
rect 1353 16033 1439 16089
rect 1495 16033 1581 16089
rect 1637 16033 1723 16089
rect 1779 16033 1865 16089
rect 1921 16033 2007 16089
rect 2063 16033 2149 16089
rect 2205 16033 2291 16089
rect 2347 16033 2433 16089
rect 2489 16033 2575 16089
rect 2631 16033 2717 16089
rect 2773 16033 2859 16089
rect 2915 16033 3001 16089
rect 3057 16033 3143 16089
rect 3199 16033 3285 16089
rect 3341 16033 3427 16089
rect 3483 16033 3569 16089
rect 3625 16033 3711 16089
rect 3767 16033 3853 16089
rect 3909 16033 3995 16089
rect 4051 16033 4137 16089
rect 4193 16033 4279 16089
rect 4335 16033 4421 16089
rect 4477 16033 4563 16089
rect 4619 16033 4705 16089
rect 4761 16033 4847 16089
rect 4903 16033 4989 16089
rect 5045 16033 5131 16089
rect 5187 16033 5273 16089
rect 5329 16033 5415 16089
rect 5471 16033 5557 16089
rect 5613 16033 5699 16089
rect 5755 16033 5841 16089
rect 5897 16033 5983 16089
rect 6039 16033 6125 16089
rect 6181 16033 6267 16089
rect 6323 16033 6409 16089
rect 6465 16033 6551 16089
rect 6607 16033 6693 16089
rect 6749 16033 6835 16089
rect 6891 16033 6977 16089
rect 7033 16033 7119 16089
rect 7175 16033 7261 16089
rect 7317 16033 7403 16089
rect 7459 16033 7545 16089
rect 7601 16033 7687 16089
rect 7743 16033 7829 16089
rect 7885 16033 7971 16089
rect 8027 16033 8113 16089
rect 8169 16033 8255 16089
rect 8311 16033 8397 16089
rect 8453 16033 8539 16089
rect 8595 16033 8681 16089
rect 8737 16033 8823 16089
rect 8879 16033 8965 16089
rect 9021 16033 9107 16089
rect 9163 16033 9249 16089
rect 9305 16033 9391 16089
rect 9447 16033 9533 16089
rect 9589 16033 9675 16089
rect 9731 16033 9817 16089
rect 9873 16033 9959 16089
rect 10015 16033 10101 16089
rect 10157 16033 10243 16089
rect 10299 16033 10385 16089
rect 10441 16033 10527 16089
rect 10583 16033 10669 16089
rect 10725 16033 10811 16089
rect 10867 16033 10953 16089
rect 11009 16033 11095 16089
rect 11151 16033 11237 16089
rect 11293 16033 11379 16089
rect 11435 16033 11521 16089
rect 11577 16033 11663 16089
rect 11719 16033 11805 16089
rect 11861 16033 11947 16089
rect 12003 16033 12089 16089
rect 12145 16033 12231 16089
rect 12287 16033 12373 16089
rect 12429 16033 12515 16089
rect 12571 16033 12657 16089
rect 12713 16033 12799 16089
rect 12855 16033 12941 16089
rect 12997 16033 13083 16089
rect 13139 16033 13225 16089
rect 13281 16033 13367 16089
rect 13423 16033 13509 16089
rect 13565 16033 13651 16089
rect 13707 16033 13793 16089
rect 13849 16033 13935 16089
rect 13991 16033 14077 16089
rect 14133 16033 14219 16089
rect 14275 16033 14361 16089
rect 14417 16033 14503 16089
rect 14559 16033 14645 16089
rect 14701 16033 14787 16089
rect 14843 16033 14853 16089
rect 151 15947 14853 16033
rect 151 15891 161 15947
rect 217 15891 303 15947
rect 359 15891 445 15947
rect 501 15891 587 15947
rect 643 15891 729 15947
rect 785 15891 871 15947
rect 927 15891 1013 15947
rect 1069 15891 1155 15947
rect 1211 15891 1297 15947
rect 1353 15891 1439 15947
rect 1495 15891 1581 15947
rect 1637 15891 1723 15947
rect 1779 15891 1865 15947
rect 1921 15891 2007 15947
rect 2063 15891 2149 15947
rect 2205 15891 2291 15947
rect 2347 15891 2433 15947
rect 2489 15891 2575 15947
rect 2631 15891 2717 15947
rect 2773 15891 2859 15947
rect 2915 15891 3001 15947
rect 3057 15891 3143 15947
rect 3199 15891 3285 15947
rect 3341 15891 3427 15947
rect 3483 15891 3569 15947
rect 3625 15891 3711 15947
rect 3767 15891 3853 15947
rect 3909 15891 3995 15947
rect 4051 15891 4137 15947
rect 4193 15891 4279 15947
rect 4335 15891 4421 15947
rect 4477 15891 4563 15947
rect 4619 15891 4705 15947
rect 4761 15891 4847 15947
rect 4903 15891 4989 15947
rect 5045 15891 5131 15947
rect 5187 15891 5273 15947
rect 5329 15891 5415 15947
rect 5471 15891 5557 15947
rect 5613 15891 5699 15947
rect 5755 15891 5841 15947
rect 5897 15891 5983 15947
rect 6039 15891 6125 15947
rect 6181 15891 6267 15947
rect 6323 15891 6409 15947
rect 6465 15891 6551 15947
rect 6607 15891 6693 15947
rect 6749 15891 6835 15947
rect 6891 15891 6977 15947
rect 7033 15891 7119 15947
rect 7175 15891 7261 15947
rect 7317 15891 7403 15947
rect 7459 15891 7545 15947
rect 7601 15891 7687 15947
rect 7743 15891 7829 15947
rect 7885 15891 7971 15947
rect 8027 15891 8113 15947
rect 8169 15891 8255 15947
rect 8311 15891 8397 15947
rect 8453 15891 8539 15947
rect 8595 15891 8681 15947
rect 8737 15891 8823 15947
rect 8879 15891 8965 15947
rect 9021 15891 9107 15947
rect 9163 15891 9249 15947
rect 9305 15891 9391 15947
rect 9447 15891 9533 15947
rect 9589 15891 9675 15947
rect 9731 15891 9817 15947
rect 9873 15891 9959 15947
rect 10015 15891 10101 15947
rect 10157 15891 10243 15947
rect 10299 15891 10385 15947
rect 10441 15891 10527 15947
rect 10583 15891 10669 15947
rect 10725 15891 10811 15947
rect 10867 15891 10953 15947
rect 11009 15891 11095 15947
rect 11151 15891 11237 15947
rect 11293 15891 11379 15947
rect 11435 15891 11521 15947
rect 11577 15891 11663 15947
rect 11719 15891 11805 15947
rect 11861 15891 11947 15947
rect 12003 15891 12089 15947
rect 12145 15891 12231 15947
rect 12287 15891 12373 15947
rect 12429 15891 12515 15947
rect 12571 15891 12657 15947
rect 12713 15891 12799 15947
rect 12855 15891 12941 15947
rect 12997 15891 13083 15947
rect 13139 15891 13225 15947
rect 13281 15891 13367 15947
rect 13423 15891 13509 15947
rect 13565 15891 13651 15947
rect 13707 15891 13793 15947
rect 13849 15891 13935 15947
rect 13991 15891 14077 15947
rect 14133 15891 14219 15947
rect 14275 15891 14361 15947
rect 14417 15891 14503 15947
rect 14559 15891 14645 15947
rect 14701 15891 14787 15947
rect 14843 15891 14853 15947
rect 151 15805 14853 15891
rect 151 15749 161 15805
rect 217 15749 303 15805
rect 359 15749 445 15805
rect 501 15749 587 15805
rect 643 15749 729 15805
rect 785 15749 871 15805
rect 927 15749 1013 15805
rect 1069 15749 1155 15805
rect 1211 15749 1297 15805
rect 1353 15749 1439 15805
rect 1495 15749 1581 15805
rect 1637 15749 1723 15805
rect 1779 15749 1865 15805
rect 1921 15749 2007 15805
rect 2063 15749 2149 15805
rect 2205 15749 2291 15805
rect 2347 15749 2433 15805
rect 2489 15749 2575 15805
rect 2631 15749 2717 15805
rect 2773 15749 2859 15805
rect 2915 15749 3001 15805
rect 3057 15749 3143 15805
rect 3199 15749 3285 15805
rect 3341 15749 3427 15805
rect 3483 15749 3569 15805
rect 3625 15749 3711 15805
rect 3767 15749 3853 15805
rect 3909 15749 3995 15805
rect 4051 15749 4137 15805
rect 4193 15749 4279 15805
rect 4335 15749 4421 15805
rect 4477 15749 4563 15805
rect 4619 15749 4705 15805
rect 4761 15749 4847 15805
rect 4903 15749 4989 15805
rect 5045 15749 5131 15805
rect 5187 15749 5273 15805
rect 5329 15749 5415 15805
rect 5471 15749 5557 15805
rect 5613 15749 5699 15805
rect 5755 15749 5841 15805
rect 5897 15749 5983 15805
rect 6039 15749 6125 15805
rect 6181 15749 6267 15805
rect 6323 15749 6409 15805
rect 6465 15749 6551 15805
rect 6607 15749 6693 15805
rect 6749 15749 6835 15805
rect 6891 15749 6977 15805
rect 7033 15749 7119 15805
rect 7175 15749 7261 15805
rect 7317 15749 7403 15805
rect 7459 15749 7545 15805
rect 7601 15749 7687 15805
rect 7743 15749 7829 15805
rect 7885 15749 7971 15805
rect 8027 15749 8113 15805
rect 8169 15749 8255 15805
rect 8311 15749 8397 15805
rect 8453 15749 8539 15805
rect 8595 15749 8681 15805
rect 8737 15749 8823 15805
rect 8879 15749 8965 15805
rect 9021 15749 9107 15805
rect 9163 15749 9249 15805
rect 9305 15749 9391 15805
rect 9447 15749 9533 15805
rect 9589 15749 9675 15805
rect 9731 15749 9817 15805
rect 9873 15749 9959 15805
rect 10015 15749 10101 15805
rect 10157 15749 10243 15805
rect 10299 15749 10385 15805
rect 10441 15749 10527 15805
rect 10583 15749 10669 15805
rect 10725 15749 10811 15805
rect 10867 15749 10953 15805
rect 11009 15749 11095 15805
rect 11151 15749 11237 15805
rect 11293 15749 11379 15805
rect 11435 15749 11521 15805
rect 11577 15749 11663 15805
rect 11719 15749 11805 15805
rect 11861 15749 11947 15805
rect 12003 15749 12089 15805
rect 12145 15749 12231 15805
rect 12287 15749 12373 15805
rect 12429 15749 12515 15805
rect 12571 15749 12657 15805
rect 12713 15749 12799 15805
rect 12855 15749 12941 15805
rect 12997 15749 13083 15805
rect 13139 15749 13225 15805
rect 13281 15749 13367 15805
rect 13423 15749 13509 15805
rect 13565 15749 13651 15805
rect 13707 15749 13793 15805
rect 13849 15749 13935 15805
rect 13991 15749 14077 15805
rect 14133 15749 14219 15805
rect 14275 15749 14361 15805
rect 14417 15749 14503 15805
rect 14559 15749 14645 15805
rect 14701 15749 14787 15805
rect 14843 15749 14853 15805
rect 151 15663 14853 15749
rect 151 15607 161 15663
rect 217 15607 303 15663
rect 359 15607 445 15663
rect 501 15607 587 15663
rect 643 15607 729 15663
rect 785 15607 871 15663
rect 927 15607 1013 15663
rect 1069 15607 1155 15663
rect 1211 15607 1297 15663
rect 1353 15607 1439 15663
rect 1495 15607 1581 15663
rect 1637 15607 1723 15663
rect 1779 15607 1865 15663
rect 1921 15607 2007 15663
rect 2063 15607 2149 15663
rect 2205 15607 2291 15663
rect 2347 15607 2433 15663
rect 2489 15607 2575 15663
rect 2631 15607 2717 15663
rect 2773 15607 2859 15663
rect 2915 15607 3001 15663
rect 3057 15607 3143 15663
rect 3199 15607 3285 15663
rect 3341 15607 3427 15663
rect 3483 15607 3569 15663
rect 3625 15607 3711 15663
rect 3767 15607 3853 15663
rect 3909 15607 3995 15663
rect 4051 15607 4137 15663
rect 4193 15607 4279 15663
rect 4335 15607 4421 15663
rect 4477 15607 4563 15663
rect 4619 15607 4705 15663
rect 4761 15607 4847 15663
rect 4903 15607 4989 15663
rect 5045 15607 5131 15663
rect 5187 15607 5273 15663
rect 5329 15607 5415 15663
rect 5471 15607 5557 15663
rect 5613 15607 5699 15663
rect 5755 15607 5841 15663
rect 5897 15607 5983 15663
rect 6039 15607 6125 15663
rect 6181 15607 6267 15663
rect 6323 15607 6409 15663
rect 6465 15607 6551 15663
rect 6607 15607 6693 15663
rect 6749 15607 6835 15663
rect 6891 15607 6977 15663
rect 7033 15607 7119 15663
rect 7175 15607 7261 15663
rect 7317 15607 7403 15663
rect 7459 15607 7545 15663
rect 7601 15607 7687 15663
rect 7743 15607 7829 15663
rect 7885 15607 7971 15663
rect 8027 15607 8113 15663
rect 8169 15607 8255 15663
rect 8311 15607 8397 15663
rect 8453 15607 8539 15663
rect 8595 15607 8681 15663
rect 8737 15607 8823 15663
rect 8879 15607 8965 15663
rect 9021 15607 9107 15663
rect 9163 15607 9249 15663
rect 9305 15607 9391 15663
rect 9447 15607 9533 15663
rect 9589 15607 9675 15663
rect 9731 15607 9817 15663
rect 9873 15607 9959 15663
rect 10015 15607 10101 15663
rect 10157 15607 10243 15663
rect 10299 15607 10385 15663
rect 10441 15607 10527 15663
rect 10583 15607 10669 15663
rect 10725 15607 10811 15663
rect 10867 15607 10953 15663
rect 11009 15607 11095 15663
rect 11151 15607 11237 15663
rect 11293 15607 11379 15663
rect 11435 15607 11521 15663
rect 11577 15607 11663 15663
rect 11719 15607 11805 15663
rect 11861 15607 11947 15663
rect 12003 15607 12089 15663
rect 12145 15607 12231 15663
rect 12287 15607 12373 15663
rect 12429 15607 12515 15663
rect 12571 15607 12657 15663
rect 12713 15607 12799 15663
rect 12855 15607 12941 15663
rect 12997 15607 13083 15663
rect 13139 15607 13225 15663
rect 13281 15607 13367 15663
rect 13423 15607 13509 15663
rect 13565 15607 13651 15663
rect 13707 15607 13793 15663
rect 13849 15607 13935 15663
rect 13991 15607 14077 15663
rect 14133 15607 14219 15663
rect 14275 15607 14361 15663
rect 14417 15607 14503 15663
rect 14559 15607 14645 15663
rect 14701 15607 14787 15663
rect 14843 15607 14853 15663
rect 151 15521 14853 15607
rect 151 15465 161 15521
rect 217 15465 303 15521
rect 359 15465 445 15521
rect 501 15465 587 15521
rect 643 15465 729 15521
rect 785 15465 871 15521
rect 927 15465 1013 15521
rect 1069 15465 1155 15521
rect 1211 15465 1297 15521
rect 1353 15465 1439 15521
rect 1495 15465 1581 15521
rect 1637 15465 1723 15521
rect 1779 15465 1865 15521
rect 1921 15465 2007 15521
rect 2063 15465 2149 15521
rect 2205 15465 2291 15521
rect 2347 15465 2433 15521
rect 2489 15465 2575 15521
rect 2631 15465 2717 15521
rect 2773 15465 2859 15521
rect 2915 15465 3001 15521
rect 3057 15465 3143 15521
rect 3199 15465 3285 15521
rect 3341 15465 3427 15521
rect 3483 15465 3569 15521
rect 3625 15465 3711 15521
rect 3767 15465 3853 15521
rect 3909 15465 3995 15521
rect 4051 15465 4137 15521
rect 4193 15465 4279 15521
rect 4335 15465 4421 15521
rect 4477 15465 4563 15521
rect 4619 15465 4705 15521
rect 4761 15465 4847 15521
rect 4903 15465 4989 15521
rect 5045 15465 5131 15521
rect 5187 15465 5273 15521
rect 5329 15465 5415 15521
rect 5471 15465 5557 15521
rect 5613 15465 5699 15521
rect 5755 15465 5841 15521
rect 5897 15465 5983 15521
rect 6039 15465 6125 15521
rect 6181 15465 6267 15521
rect 6323 15465 6409 15521
rect 6465 15465 6551 15521
rect 6607 15465 6693 15521
rect 6749 15465 6835 15521
rect 6891 15465 6977 15521
rect 7033 15465 7119 15521
rect 7175 15465 7261 15521
rect 7317 15465 7403 15521
rect 7459 15465 7545 15521
rect 7601 15465 7687 15521
rect 7743 15465 7829 15521
rect 7885 15465 7971 15521
rect 8027 15465 8113 15521
rect 8169 15465 8255 15521
rect 8311 15465 8397 15521
rect 8453 15465 8539 15521
rect 8595 15465 8681 15521
rect 8737 15465 8823 15521
rect 8879 15465 8965 15521
rect 9021 15465 9107 15521
rect 9163 15465 9249 15521
rect 9305 15465 9391 15521
rect 9447 15465 9533 15521
rect 9589 15465 9675 15521
rect 9731 15465 9817 15521
rect 9873 15465 9959 15521
rect 10015 15465 10101 15521
rect 10157 15465 10243 15521
rect 10299 15465 10385 15521
rect 10441 15465 10527 15521
rect 10583 15465 10669 15521
rect 10725 15465 10811 15521
rect 10867 15465 10953 15521
rect 11009 15465 11095 15521
rect 11151 15465 11237 15521
rect 11293 15465 11379 15521
rect 11435 15465 11521 15521
rect 11577 15465 11663 15521
rect 11719 15465 11805 15521
rect 11861 15465 11947 15521
rect 12003 15465 12089 15521
rect 12145 15465 12231 15521
rect 12287 15465 12373 15521
rect 12429 15465 12515 15521
rect 12571 15465 12657 15521
rect 12713 15465 12799 15521
rect 12855 15465 12941 15521
rect 12997 15465 13083 15521
rect 13139 15465 13225 15521
rect 13281 15465 13367 15521
rect 13423 15465 13509 15521
rect 13565 15465 13651 15521
rect 13707 15465 13793 15521
rect 13849 15465 13935 15521
rect 13991 15465 14077 15521
rect 14133 15465 14219 15521
rect 14275 15465 14361 15521
rect 14417 15465 14503 15521
rect 14559 15465 14645 15521
rect 14701 15465 14787 15521
rect 14843 15465 14853 15521
rect 151 15379 14853 15465
rect 151 15323 161 15379
rect 217 15323 303 15379
rect 359 15323 445 15379
rect 501 15323 587 15379
rect 643 15323 729 15379
rect 785 15323 871 15379
rect 927 15323 1013 15379
rect 1069 15323 1155 15379
rect 1211 15323 1297 15379
rect 1353 15323 1439 15379
rect 1495 15323 1581 15379
rect 1637 15323 1723 15379
rect 1779 15323 1865 15379
rect 1921 15323 2007 15379
rect 2063 15323 2149 15379
rect 2205 15323 2291 15379
rect 2347 15323 2433 15379
rect 2489 15323 2575 15379
rect 2631 15323 2717 15379
rect 2773 15323 2859 15379
rect 2915 15323 3001 15379
rect 3057 15323 3143 15379
rect 3199 15323 3285 15379
rect 3341 15323 3427 15379
rect 3483 15323 3569 15379
rect 3625 15323 3711 15379
rect 3767 15323 3853 15379
rect 3909 15323 3995 15379
rect 4051 15323 4137 15379
rect 4193 15323 4279 15379
rect 4335 15323 4421 15379
rect 4477 15323 4563 15379
rect 4619 15323 4705 15379
rect 4761 15323 4847 15379
rect 4903 15323 4989 15379
rect 5045 15323 5131 15379
rect 5187 15323 5273 15379
rect 5329 15323 5415 15379
rect 5471 15323 5557 15379
rect 5613 15323 5699 15379
rect 5755 15323 5841 15379
rect 5897 15323 5983 15379
rect 6039 15323 6125 15379
rect 6181 15323 6267 15379
rect 6323 15323 6409 15379
rect 6465 15323 6551 15379
rect 6607 15323 6693 15379
rect 6749 15323 6835 15379
rect 6891 15323 6977 15379
rect 7033 15323 7119 15379
rect 7175 15323 7261 15379
rect 7317 15323 7403 15379
rect 7459 15323 7545 15379
rect 7601 15323 7687 15379
rect 7743 15323 7829 15379
rect 7885 15323 7971 15379
rect 8027 15323 8113 15379
rect 8169 15323 8255 15379
rect 8311 15323 8397 15379
rect 8453 15323 8539 15379
rect 8595 15323 8681 15379
rect 8737 15323 8823 15379
rect 8879 15323 8965 15379
rect 9021 15323 9107 15379
rect 9163 15323 9249 15379
rect 9305 15323 9391 15379
rect 9447 15323 9533 15379
rect 9589 15323 9675 15379
rect 9731 15323 9817 15379
rect 9873 15323 9959 15379
rect 10015 15323 10101 15379
rect 10157 15323 10243 15379
rect 10299 15323 10385 15379
rect 10441 15323 10527 15379
rect 10583 15323 10669 15379
rect 10725 15323 10811 15379
rect 10867 15323 10953 15379
rect 11009 15323 11095 15379
rect 11151 15323 11237 15379
rect 11293 15323 11379 15379
rect 11435 15323 11521 15379
rect 11577 15323 11663 15379
rect 11719 15323 11805 15379
rect 11861 15323 11947 15379
rect 12003 15323 12089 15379
rect 12145 15323 12231 15379
rect 12287 15323 12373 15379
rect 12429 15323 12515 15379
rect 12571 15323 12657 15379
rect 12713 15323 12799 15379
rect 12855 15323 12941 15379
rect 12997 15323 13083 15379
rect 13139 15323 13225 15379
rect 13281 15323 13367 15379
rect 13423 15323 13509 15379
rect 13565 15323 13651 15379
rect 13707 15323 13793 15379
rect 13849 15323 13935 15379
rect 13991 15323 14077 15379
rect 14133 15323 14219 15379
rect 14275 15323 14361 15379
rect 14417 15323 14503 15379
rect 14559 15323 14645 15379
rect 14701 15323 14787 15379
rect 14843 15323 14853 15379
rect 151 15237 14853 15323
rect 151 15181 161 15237
rect 217 15181 303 15237
rect 359 15181 445 15237
rect 501 15181 587 15237
rect 643 15181 729 15237
rect 785 15181 871 15237
rect 927 15181 1013 15237
rect 1069 15181 1155 15237
rect 1211 15181 1297 15237
rect 1353 15181 1439 15237
rect 1495 15181 1581 15237
rect 1637 15181 1723 15237
rect 1779 15181 1865 15237
rect 1921 15181 2007 15237
rect 2063 15181 2149 15237
rect 2205 15181 2291 15237
rect 2347 15181 2433 15237
rect 2489 15181 2575 15237
rect 2631 15181 2717 15237
rect 2773 15181 2859 15237
rect 2915 15181 3001 15237
rect 3057 15181 3143 15237
rect 3199 15181 3285 15237
rect 3341 15181 3427 15237
rect 3483 15181 3569 15237
rect 3625 15181 3711 15237
rect 3767 15181 3853 15237
rect 3909 15181 3995 15237
rect 4051 15181 4137 15237
rect 4193 15181 4279 15237
rect 4335 15181 4421 15237
rect 4477 15181 4563 15237
rect 4619 15181 4705 15237
rect 4761 15181 4847 15237
rect 4903 15181 4989 15237
rect 5045 15181 5131 15237
rect 5187 15181 5273 15237
rect 5329 15181 5415 15237
rect 5471 15181 5557 15237
rect 5613 15181 5699 15237
rect 5755 15181 5841 15237
rect 5897 15181 5983 15237
rect 6039 15181 6125 15237
rect 6181 15181 6267 15237
rect 6323 15181 6409 15237
rect 6465 15181 6551 15237
rect 6607 15181 6693 15237
rect 6749 15181 6835 15237
rect 6891 15181 6977 15237
rect 7033 15181 7119 15237
rect 7175 15181 7261 15237
rect 7317 15181 7403 15237
rect 7459 15181 7545 15237
rect 7601 15181 7687 15237
rect 7743 15181 7829 15237
rect 7885 15181 7971 15237
rect 8027 15181 8113 15237
rect 8169 15181 8255 15237
rect 8311 15181 8397 15237
rect 8453 15181 8539 15237
rect 8595 15181 8681 15237
rect 8737 15181 8823 15237
rect 8879 15181 8965 15237
rect 9021 15181 9107 15237
rect 9163 15181 9249 15237
rect 9305 15181 9391 15237
rect 9447 15181 9533 15237
rect 9589 15181 9675 15237
rect 9731 15181 9817 15237
rect 9873 15181 9959 15237
rect 10015 15181 10101 15237
rect 10157 15181 10243 15237
rect 10299 15181 10385 15237
rect 10441 15181 10527 15237
rect 10583 15181 10669 15237
rect 10725 15181 10811 15237
rect 10867 15181 10953 15237
rect 11009 15181 11095 15237
rect 11151 15181 11237 15237
rect 11293 15181 11379 15237
rect 11435 15181 11521 15237
rect 11577 15181 11663 15237
rect 11719 15181 11805 15237
rect 11861 15181 11947 15237
rect 12003 15181 12089 15237
rect 12145 15181 12231 15237
rect 12287 15181 12373 15237
rect 12429 15181 12515 15237
rect 12571 15181 12657 15237
rect 12713 15181 12799 15237
rect 12855 15181 12941 15237
rect 12997 15181 13083 15237
rect 13139 15181 13225 15237
rect 13281 15181 13367 15237
rect 13423 15181 13509 15237
rect 13565 15181 13651 15237
rect 13707 15181 13793 15237
rect 13849 15181 13935 15237
rect 13991 15181 14077 15237
rect 14133 15181 14219 15237
rect 14275 15181 14361 15237
rect 14417 15181 14503 15237
rect 14559 15181 14645 15237
rect 14701 15181 14787 15237
rect 14843 15181 14853 15237
rect 151 15095 14853 15181
rect 151 15039 161 15095
rect 217 15039 303 15095
rect 359 15039 445 15095
rect 501 15039 587 15095
rect 643 15039 729 15095
rect 785 15039 871 15095
rect 927 15039 1013 15095
rect 1069 15039 1155 15095
rect 1211 15039 1297 15095
rect 1353 15039 1439 15095
rect 1495 15039 1581 15095
rect 1637 15039 1723 15095
rect 1779 15039 1865 15095
rect 1921 15039 2007 15095
rect 2063 15039 2149 15095
rect 2205 15039 2291 15095
rect 2347 15039 2433 15095
rect 2489 15039 2575 15095
rect 2631 15039 2717 15095
rect 2773 15039 2859 15095
rect 2915 15039 3001 15095
rect 3057 15039 3143 15095
rect 3199 15039 3285 15095
rect 3341 15039 3427 15095
rect 3483 15039 3569 15095
rect 3625 15039 3711 15095
rect 3767 15039 3853 15095
rect 3909 15039 3995 15095
rect 4051 15039 4137 15095
rect 4193 15039 4279 15095
rect 4335 15039 4421 15095
rect 4477 15039 4563 15095
rect 4619 15039 4705 15095
rect 4761 15039 4847 15095
rect 4903 15039 4989 15095
rect 5045 15039 5131 15095
rect 5187 15039 5273 15095
rect 5329 15039 5415 15095
rect 5471 15039 5557 15095
rect 5613 15039 5699 15095
rect 5755 15039 5841 15095
rect 5897 15039 5983 15095
rect 6039 15039 6125 15095
rect 6181 15039 6267 15095
rect 6323 15039 6409 15095
rect 6465 15039 6551 15095
rect 6607 15039 6693 15095
rect 6749 15039 6835 15095
rect 6891 15039 6977 15095
rect 7033 15039 7119 15095
rect 7175 15039 7261 15095
rect 7317 15039 7403 15095
rect 7459 15039 7545 15095
rect 7601 15039 7687 15095
rect 7743 15039 7829 15095
rect 7885 15039 7971 15095
rect 8027 15039 8113 15095
rect 8169 15039 8255 15095
rect 8311 15039 8397 15095
rect 8453 15039 8539 15095
rect 8595 15039 8681 15095
rect 8737 15039 8823 15095
rect 8879 15039 8965 15095
rect 9021 15039 9107 15095
rect 9163 15039 9249 15095
rect 9305 15039 9391 15095
rect 9447 15039 9533 15095
rect 9589 15039 9675 15095
rect 9731 15039 9817 15095
rect 9873 15039 9959 15095
rect 10015 15039 10101 15095
rect 10157 15039 10243 15095
rect 10299 15039 10385 15095
rect 10441 15039 10527 15095
rect 10583 15039 10669 15095
rect 10725 15039 10811 15095
rect 10867 15039 10953 15095
rect 11009 15039 11095 15095
rect 11151 15039 11237 15095
rect 11293 15039 11379 15095
rect 11435 15039 11521 15095
rect 11577 15039 11663 15095
rect 11719 15039 11805 15095
rect 11861 15039 11947 15095
rect 12003 15039 12089 15095
rect 12145 15039 12231 15095
rect 12287 15039 12373 15095
rect 12429 15039 12515 15095
rect 12571 15039 12657 15095
rect 12713 15039 12799 15095
rect 12855 15039 12941 15095
rect 12997 15039 13083 15095
rect 13139 15039 13225 15095
rect 13281 15039 13367 15095
rect 13423 15039 13509 15095
rect 13565 15039 13651 15095
rect 13707 15039 13793 15095
rect 13849 15039 13935 15095
rect 13991 15039 14077 15095
rect 14133 15039 14219 15095
rect 14275 15039 14361 15095
rect 14417 15039 14503 15095
rect 14559 15039 14645 15095
rect 14701 15039 14787 15095
rect 14843 15039 14853 15095
rect 151 14953 14853 15039
rect 151 14897 161 14953
rect 217 14897 303 14953
rect 359 14897 445 14953
rect 501 14897 587 14953
rect 643 14897 729 14953
rect 785 14897 871 14953
rect 927 14897 1013 14953
rect 1069 14897 1155 14953
rect 1211 14897 1297 14953
rect 1353 14897 1439 14953
rect 1495 14897 1581 14953
rect 1637 14897 1723 14953
rect 1779 14897 1865 14953
rect 1921 14897 2007 14953
rect 2063 14897 2149 14953
rect 2205 14897 2291 14953
rect 2347 14897 2433 14953
rect 2489 14897 2575 14953
rect 2631 14897 2717 14953
rect 2773 14897 2859 14953
rect 2915 14897 3001 14953
rect 3057 14897 3143 14953
rect 3199 14897 3285 14953
rect 3341 14897 3427 14953
rect 3483 14897 3569 14953
rect 3625 14897 3711 14953
rect 3767 14897 3853 14953
rect 3909 14897 3995 14953
rect 4051 14897 4137 14953
rect 4193 14897 4279 14953
rect 4335 14897 4421 14953
rect 4477 14897 4563 14953
rect 4619 14897 4705 14953
rect 4761 14897 4847 14953
rect 4903 14897 4989 14953
rect 5045 14897 5131 14953
rect 5187 14897 5273 14953
rect 5329 14897 5415 14953
rect 5471 14897 5557 14953
rect 5613 14897 5699 14953
rect 5755 14897 5841 14953
rect 5897 14897 5983 14953
rect 6039 14897 6125 14953
rect 6181 14897 6267 14953
rect 6323 14897 6409 14953
rect 6465 14897 6551 14953
rect 6607 14897 6693 14953
rect 6749 14897 6835 14953
rect 6891 14897 6977 14953
rect 7033 14897 7119 14953
rect 7175 14897 7261 14953
rect 7317 14897 7403 14953
rect 7459 14897 7545 14953
rect 7601 14897 7687 14953
rect 7743 14897 7829 14953
rect 7885 14897 7971 14953
rect 8027 14897 8113 14953
rect 8169 14897 8255 14953
rect 8311 14897 8397 14953
rect 8453 14897 8539 14953
rect 8595 14897 8681 14953
rect 8737 14897 8823 14953
rect 8879 14897 8965 14953
rect 9021 14897 9107 14953
rect 9163 14897 9249 14953
rect 9305 14897 9391 14953
rect 9447 14897 9533 14953
rect 9589 14897 9675 14953
rect 9731 14897 9817 14953
rect 9873 14897 9959 14953
rect 10015 14897 10101 14953
rect 10157 14897 10243 14953
rect 10299 14897 10385 14953
rect 10441 14897 10527 14953
rect 10583 14897 10669 14953
rect 10725 14897 10811 14953
rect 10867 14897 10953 14953
rect 11009 14897 11095 14953
rect 11151 14897 11237 14953
rect 11293 14897 11379 14953
rect 11435 14897 11521 14953
rect 11577 14897 11663 14953
rect 11719 14897 11805 14953
rect 11861 14897 11947 14953
rect 12003 14897 12089 14953
rect 12145 14897 12231 14953
rect 12287 14897 12373 14953
rect 12429 14897 12515 14953
rect 12571 14897 12657 14953
rect 12713 14897 12799 14953
rect 12855 14897 12941 14953
rect 12997 14897 13083 14953
rect 13139 14897 13225 14953
rect 13281 14897 13367 14953
rect 13423 14897 13509 14953
rect 13565 14897 13651 14953
rect 13707 14897 13793 14953
rect 13849 14897 13935 14953
rect 13991 14897 14077 14953
rect 14133 14897 14219 14953
rect 14275 14897 14361 14953
rect 14417 14897 14503 14953
rect 14559 14897 14645 14953
rect 14701 14897 14787 14953
rect 14843 14897 14853 14953
rect 151 14811 14853 14897
rect 151 14755 161 14811
rect 217 14755 303 14811
rect 359 14755 445 14811
rect 501 14755 587 14811
rect 643 14755 729 14811
rect 785 14755 871 14811
rect 927 14755 1013 14811
rect 1069 14755 1155 14811
rect 1211 14755 1297 14811
rect 1353 14755 1439 14811
rect 1495 14755 1581 14811
rect 1637 14755 1723 14811
rect 1779 14755 1865 14811
rect 1921 14755 2007 14811
rect 2063 14755 2149 14811
rect 2205 14755 2291 14811
rect 2347 14755 2433 14811
rect 2489 14755 2575 14811
rect 2631 14755 2717 14811
rect 2773 14755 2859 14811
rect 2915 14755 3001 14811
rect 3057 14755 3143 14811
rect 3199 14755 3285 14811
rect 3341 14755 3427 14811
rect 3483 14755 3569 14811
rect 3625 14755 3711 14811
rect 3767 14755 3853 14811
rect 3909 14755 3995 14811
rect 4051 14755 4137 14811
rect 4193 14755 4279 14811
rect 4335 14755 4421 14811
rect 4477 14755 4563 14811
rect 4619 14755 4705 14811
rect 4761 14755 4847 14811
rect 4903 14755 4989 14811
rect 5045 14755 5131 14811
rect 5187 14755 5273 14811
rect 5329 14755 5415 14811
rect 5471 14755 5557 14811
rect 5613 14755 5699 14811
rect 5755 14755 5841 14811
rect 5897 14755 5983 14811
rect 6039 14755 6125 14811
rect 6181 14755 6267 14811
rect 6323 14755 6409 14811
rect 6465 14755 6551 14811
rect 6607 14755 6693 14811
rect 6749 14755 6835 14811
rect 6891 14755 6977 14811
rect 7033 14755 7119 14811
rect 7175 14755 7261 14811
rect 7317 14755 7403 14811
rect 7459 14755 7545 14811
rect 7601 14755 7687 14811
rect 7743 14755 7829 14811
rect 7885 14755 7971 14811
rect 8027 14755 8113 14811
rect 8169 14755 8255 14811
rect 8311 14755 8397 14811
rect 8453 14755 8539 14811
rect 8595 14755 8681 14811
rect 8737 14755 8823 14811
rect 8879 14755 8965 14811
rect 9021 14755 9107 14811
rect 9163 14755 9249 14811
rect 9305 14755 9391 14811
rect 9447 14755 9533 14811
rect 9589 14755 9675 14811
rect 9731 14755 9817 14811
rect 9873 14755 9959 14811
rect 10015 14755 10101 14811
rect 10157 14755 10243 14811
rect 10299 14755 10385 14811
rect 10441 14755 10527 14811
rect 10583 14755 10669 14811
rect 10725 14755 10811 14811
rect 10867 14755 10953 14811
rect 11009 14755 11095 14811
rect 11151 14755 11237 14811
rect 11293 14755 11379 14811
rect 11435 14755 11521 14811
rect 11577 14755 11663 14811
rect 11719 14755 11805 14811
rect 11861 14755 11947 14811
rect 12003 14755 12089 14811
rect 12145 14755 12231 14811
rect 12287 14755 12373 14811
rect 12429 14755 12515 14811
rect 12571 14755 12657 14811
rect 12713 14755 12799 14811
rect 12855 14755 12941 14811
rect 12997 14755 13083 14811
rect 13139 14755 13225 14811
rect 13281 14755 13367 14811
rect 13423 14755 13509 14811
rect 13565 14755 13651 14811
rect 13707 14755 13793 14811
rect 13849 14755 13935 14811
rect 13991 14755 14077 14811
rect 14133 14755 14219 14811
rect 14275 14755 14361 14811
rect 14417 14755 14503 14811
rect 14559 14755 14645 14811
rect 14701 14755 14787 14811
rect 14843 14755 14853 14811
rect 151 14669 14853 14755
rect 151 14613 161 14669
rect 217 14613 303 14669
rect 359 14613 445 14669
rect 501 14613 587 14669
rect 643 14613 729 14669
rect 785 14613 871 14669
rect 927 14613 1013 14669
rect 1069 14613 1155 14669
rect 1211 14613 1297 14669
rect 1353 14613 1439 14669
rect 1495 14613 1581 14669
rect 1637 14613 1723 14669
rect 1779 14613 1865 14669
rect 1921 14613 2007 14669
rect 2063 14613 2149 14669
rect 2205 14613 2291 14669
rect 2347 14613 2433 14669
rect 2489 14613 2575 14669
rect 2631 14613 2717 14669
rect 2773 14613 2859 14669
rect 2915 14613 3001 14669
rect 3057 14613 3143 14669
rect 3199 14613 3285 14669
rect 3341 14613 3427 14669
rect 3483 14613 3569 14669
rect 3625 14613 3711 14669
rect 3767 14613 3853 14669
rect 3909 14613 3995 14669
rect 4051 14613 4137 14669
rect 4193 14613 4279 14669
rect 4335 14613 4421 14669
rect 4477 14613 4563 14669
rect 4619 14613 4705 14669
rect 4761 14613 4847 14669
rect 4903 14613 4989 14669
rect 5045 14613 5131 14669
rect 5187 14613 5273 14669
rect 5329 14613 5415 14669
rect 5471 14613 5557 14669
rect 5613 14613 5699 14669
rect 5755 14613 5841 14669
rect 5897 14613 5983 14669
rect 6039 14613 6125 14669
rect 6181 14613 6267 14669
rect 6323 14613 6409 14669
rect 6465 14613 6551 14669
rect 6607 14613 6693 14669
rect 6749 14613 6835 14669
rect 6891 14613 6977 14669
rect 7033 14613 7119 14669
rect 7175 14613 7261 14669
rect 7317 14613 7403 14669
rect 7459 14613 7545 14669
rect 7601 14613 7687 14669
rect 7743 14613 7829 14669
rect 7885 14613 7971 14669
rect 8027 14613 8113 14669
rect 8169 14613 8255 14669
rect 8311 14613 8397 14669
rect 8453 14613 8539 14669
rect 8595 14613 8681 14669
rect 8737 14613 8823 14669
rect 8879 14613 8965 14669
rect 9021 14613 9107 14669
rect 9163 14613 9249 14669
rect 9305 14613 9391 14669
rect 9447 14613 9533 14669
rect 9589 14613 9675 14669
rect 9731 14613 9817 14669
rect 9873 14613 9959 14669
rect 10015 14613 10101 14669
rect 10157 14613 10243 14669
rect 10299 14613 10385 14669
rect 10441 14613 10527 14669
rect 10583 14613 10669 14669
rect 10725 14613 10811 14669
rect 10867 14613 10953 14669
rect 11009 14613 11095 14669
rect 11151 14613 11237 14669
rect 11293 14613 11379 14669
rect 11435 14613 11521 14669
rect 11577 14613 11663 14669
rect 11719 14613 11805 14669
rect 11861 14613 11947 14669
rect 12003 14613 12089 14669
rect 12145 14613 12231 14669
rect 12287 14613 12373 14669
rect 12429 14613 12515 14669
rect 12571 14613 12657 14669
rect 12713 14613 12799 14669
rect 12855 14613 12941 14669
rect 12997 14613 13083 14669
rect 13139 14613 13225 14669
rect 13281 14613 13367 14669
rect 13423 14613 13509 14669
rect 13565 14613 13651 14669
rect 13707 14613 13793 14669
rect 13849 14613 13935 14669
rect 13991 14613 14077 14669
rect 14133 14613 14219 14669
rect 14275 14613 14361 14669
rect 14417 14613 14503 14669
rect 14559 14613 14645 14669
rect 14701 14613 14787 14669
rect 14843 14613 14853 14669
rect 151 14527 14853 14613
rect 151 14471 161 14527
rect 217 14471 303 14527
rect 359 14471 445 14527
rect 501 14471 587 14527
rect 643 14471 729 14527
rect 785 14471 871 14527
rect 927 14471 1013 14527
rect 1069 14471 1155 14527
rect 1211 14471 1297 14527
rect 1353 14471 1439 14527
rect 1495 14471 1581 14527
rect 1637 14471 1723 14527
rect 1779 14471 1865 14527
rect 1921 14471 2007 14527
rect 2063 14471 2149 14527
rect 2205 14471 2291 14527
rect 2347 14471 2433 14527
rect 2489 14471 2575 14527
rect 2631 14471 2717 14527
rect 2773 14471 2859 14527
rect 2915 14471 3001 14527
rect 3057 14471 3143 14527
rect 3199 14471 3285 14527
rect 3341 14471 3427 14527
rect 3483 14471 3569 14527
rect 3625 14471 3711 14527
rect 3767 14471 3853 14527
rect 3909 14471 3995 14527
rect 4051 14471 4137 14527
rect 4193 14471 4279 14527
rect 4335 14471 4421 14527
rect 4477 14471 4563 14527
rect 4619 14471 4705 14527
rect 4761 14471 4847 14527
rect 4903 14471 4989 14527
rect 5045 14471 5131 14527
rect 5187 14471 5273 14527
rect 5329 14471 5415 14527
rect 5471 14471 5557 14527
rect 5613 14471 5699 14527
rect 5755 14471 5841 14527
rect 5897 14471 5983 14527
rect 6039 14471 6125 14527
rect 6181 14471 6267 14527
rect 6323 14471 6409 14527
rect 6465 14471 6551 14527
rect 6607 14471 6693 14527
rect 6749 14471 6835 14527
rect 6891 14471 6977 14527
rect 7033 14471 7119 14527
rect 7175 14471 7261 14527
rect 7317 14471 7403 14527
rect 7459 14471 7545 14527
rect 7601 14471 7687 14527
rect 7743 14471 7829 14527
rect 7885 14471 7971 14527
rect 8027 14471 8113 14527
rect 8169 14471 8255 14527
rect 8311 14471 8397 14527
rect 8453 14471 8539 14527
rect 8595 14471 8681 14527
rect 8737 14471 8823 14527
rect 8879 14471 8965 14527
rect 9021 14471 9107 14527
rect 9163 14471 9249 14527
rect 9305 14471 9391 14527
rect 9447 14471 9533 14527
rect 9589 14471 9675 14527
rect 9731 14471 9817 14527
rect 9873 14471 9959 14527
rect 10015 14471 10101 14527
rect 10157 14471 10243 14527
rect 10299 14471 10385 14527
rect 10441 14471 10527 14527
rect 10583 14471 10669 14527
rect 10725 14471 10811 14527
rect 10867 14471 10953 14527
rect 11009 14471 11095 14527
rect 11151 14471 11237 14527
rect 11293 14471 11379 14527
rect 11435 14471 11521 14527
rect 11577 14471 11663 14527
rect 11719 14471 11805 14527
rect 11861 14471 11947 14527
rect 12003 14471 12089 14527
rect 12145 14471 12231 14527
rect 12287 14471 12373 14527
rect 12429 14471 12515 14527
rect 12571 14471 12657 14527
rect 12713 14471 12799 14527
rect 12855 14471 12941 14527
rect 12997 14471 13083 14527
rect 13139 14471 13225 14527
rect 13281 14471 13367 14527
rect 13423 14471 13509 14527
rect 13565 14471 13651 14527
rect 13707 14471 13793 14527
rect 13849 14471 13935 14527
rect 13991 14471 14077 14527
rect 14133 14471 14219 14527
rect 14275 14471 14361 14527
rect 14417 14471 14503 14527
rect 14559 14471 14645 14527
rect 14701 14471 14787 14527
rect 14843 14471 14853 14527
rect 151 14385 14853 14471
rect 151 14329 161 14385
rect 217 14329 303 14385
rect 359 14329 445 14385
rect 501 14329 587 14385
rect 643 14329 729 14385
rect 785 14329 871 14385
rect 927 14329 1013 14385
rect 1069 14329 1155 14385
rect 1211 14329 1297 14385
rect 1353 14329 1439 14385
rect 1495 14329 1581 14385
rect 1637 14329 1723 14385
rect 1779 14329 1865 14385
rect 1921 14329 2007 14385
rect 2063 14329 2149 14385
rect 2205 14329 2291 14385
rect 2347 14329 2433 14385
rect 2489 14329 2575 14385
rect 2631 14329 2717 14385
rect 2773 14329 2859 14385
rect 2915 14329 3001 14385
rect 3057 14329 3143 14385
rect 3199 14329 3285 14385
rect 3341 14329 3427 14385
rect 3483 14329 3569 14385
rect 3625 14329 3711 14385
rect 3767 14329 3853 14385
rect 3909 14329 3995 14385
rect 4051 14329 4137 14385
rect 4193 14329 4279 14385
rect 4335 14329 4421 14385
rect 4477 14329 4563 14385
rect 4619 14329 4705 14385
rect 4761 14329 4847 14385
rect 4903 14329 4989 14385
rect 5045 14329 5131 14385
rect 5187 14329 5273 14385
rect 5329 14329 5415 14385
rect 5471 14329 5557 14385
rect 5613 14329 5699 14385
rect 5755 14329 5841 14385
rect 5897 14329 5983 14385
rect 6039 14329 6125 14385
rect 6181 14329 6267 14385
rect 6323 14329 6409 14385
rect 6465 14329 6551 14385
rect 6607 14329 6693 14385
rect 6749 14329 6835 14385
rect 6891 14329 6977 14385
rect 7033 14329 7119 14385
rect 7175 14329 7261 14385
rect 7317 14329 7403 14385
rect 7459 14329 7545 14385
rect 7601 14329 7687 14385
rect 7743 14329 7829 14385
rect 7885 14329 7971 14385
rect 8027 14329 8113 14385
rect 8169 14329 8255 14385
rect 8311 14329 8397 14385
rect 8453 14329 8539 14385
rect 8595 14329 8681 14385
rect 8737 14329 8823 14385
rect 8879 14329 8965 14385
rect 9021 14329 9107 14385
rect 9163 14329 9249 14385
rect 9305 14329 9391 14385
rect 9447 14329 9533 14385
rect 9589 14329 9675 14385
rect 9731 14329 9817 14385
rect 9873 14329 9959 14385
rect 10015 14329 10101 14385
rect 10157 14329 10243 14385
rect 10299 14329 10385 14385
rect 10441 14329 10527 14385
rect 10583 14329 10669 14385
rect 10725 14329 10811 14385
rect 10867 14329 10953 14385
rect 11009 14329 11095 14385
rect 11151 14329 11237 14385
rect 11293 14329 11379 14385
rect 11435 14329 11521 14385
rect 11577 14329 11663 14385
rect 11719 14329 11805 14385
rect 11861 14329 11947 14385
rect 12003 14329 12089 14385
rect 12145 14329 12231 14385
rect 12287 14329 12373 14385
rect 12429 14329 12515 14385
rect 12571 14329 12657 14385
rect 12713 14329 12799 14385
rect 12855 14329 12941 14385
rect 12997 14329 13083 14385
rect 13139 14329 13225 14385
rect 13281 14329 13367 14385
rect 13423 14329 13509 14385
rect 13565 14329 13651 14385
rect 13707 14329 13793 14385
rect 13849 14329 13935 14385
rect 13991 14329 14077 14385
rect 14133 14329 14219 14385
rect 14275 14329 14361 14385
rect 14417 14329 14503 14385
rect 14559 14329 14645 14385
rect 14701 14329 14787 14385
rect 14843 14329 14853 14385
rect 151 14243 14853 14329
rect 151 14187 161 14243
rect 217 14187 303 14243
rect 359 14187 445 14243
rect 501 14187 587 14243
rect 643 14187 729 14243
rect 785 14187 871 14243
rect 927 14187 1013 14243
rect 1069 14187 1155 14243
rect 1211 14187 1297 14243
rect 1353 14187 1439 14243
rect 1495 14187 1581 14243
rect 1637 14187 1723 14243
rect 1779 14187 1865 14243
rect 1921 14187 2007 14243
rect 2063 14187 2149 14243
rect 2205 14187 2291 14243
rect 2347 14187 2433 14243
rect 2489 14187 2575 14243
rect 2631 14187 2717 14243
rect 2773 14187 2859 14243
rect 2915 14187 3001 14243
rect 3057 14187 3143 14243
rect 3199 14187 3285 14243
rect 3341 14187 3427 14243
rect 3483 14187 3569 14243
rect 3625 14187 3711 14243
rect 3767 14187 3853 14243
rect 3909 14187 3995 14243
rect 4051 14187 4137 14243
rect 4193 14187 4279 14243
rect 4335 14187 4421 14243
rect 4477 14187 4563 14243
rect 4619 14187 4705 14243
rect 4761 14187 4847 14243
rect 4903 14187 4989 14243
rect 5045 14187 5131 14243
rect 5187 14187 5273 14243
rect 5329 14187 5415 14243
rect 5471 14187 5557 14243
rect 5613 14187 5699 14243
rect 5755 14187 5841 14243
rect 5897 14187 5983 14243
rect 6039 14187 6125 14243
rect 6181 14187 6267 14243
rect 6323 14187 6409 14243
rect 6465 14187 6551 14243
rect 6607 14187 6693 14243
rect 6749 14187 6835 14243
rect 6891 14187 6977 14243
rect 7033 14187 7119 14243
rect 7175 14187 7261 14243
rect 7317 14187 7403 14243
rect 7459 14187 7545 14243
rect 7601 14187 7687 14243
rect 7743 14187 7829 14243
rect 7885 14187 7971 14243
rect 8027 14187 8113 14243
rect 8169 14187 8255 14243
rect 8311 14187 8397 14243
rect 8453 14187 8539 14243
rect 8595 14187 8681 14243
rect 8737 14187 8823 14243
rect 8879 14187 8965 14243
rect 9021 14187 9107 14243
rect 9163 14187 9249 14243
rect 9305 14187 9391 14243
rect 9447 14187 9533 14243
rect 9589 14187 9675 14243
rect 9731 14187 9817 14243
rect 9873 14187 9959 14243
rect 10015 14187 10101 14243
rect 10157 14187 10243 14243
rect 10299 14187 10385 14243
rect 10441 14187 10527 14243
rect 10583 14187 10669 14243
rect 10725 14187 10811 14243
rect 10867 14187 10953 14243
rect 11009 14187 11095 14243
rect 11151 14187 11237 14243
rect 11293 14187 11379 14243
rect 11435 14187 11521 14243
rect 11577 14187 11663 14243
rect 11719 14187 11805 14243
rect 11861 14187 11947 14243
rect 12003 14187 12089 14243
rect 12145 14187 12231 14243
rect 12287 14187 12373 14243
rect 12429 14187 12515 14243
rect 12571 14187 12657 14243
rect 12713 14187 12799 14243
rect 12855 14187 12941 14243
rect 12997 14187 13083 14243
rect 13139 14187 13225 14243
rect 13281 14187 13367 14243
rect 13423 14187 13509 14243
rect 13565 14187 13651 14243
rect 13707 14187 13793 14243
rect 13849 14187 13935 14243
rect 13991 14187 14077 14243
rect 14133 14187 14219 14243
rect 14275 14187 14361 14243
rect 14417 14187 14503 14243
rect 14559 14187 14645 14243
rect 14701 14187 14787 14243
rect 14843 14187 14853 14243
rect 151 14101 14853 14187
rect 151 14045 161 14101
rect 217 14045 303 14101
rect 359 14045 445 14101
rect 501 14045 587 14101
rect 643 14045 729 14101
rect 785 14045 871 14101
rect 927 14045 1013 14101
rect 1069 14045 1155 14101
rect 1211 14045 1297 14101
rect 1353 14045 1439 14101
rect 1495 14045 1581 14101
rect 1637 14045 1723 14101
rect 1779 14045 1865 14101
rect 1921 14045 2007 14101
rect 2063 14045 2149 14101
rect 2205 14045 2291 14101
rect 2347 14045 2433 14101
rect 2489 14045 2575 14101
rect 2631 14045 2717 14101
rect 2773 14045 2859 14101
rect 2915 14045 3001 14101
rect 3057 14045 3143 14101
rect 3199 14045 3285 14101
rect 3341 14045 3427 14101
rect 3483 14045 3569 14101
rect 3625 14045 3711 14101
rect 3767 14045 3853 14101
rect 3909 14045 3995 14101
rect 4051 14045 4137 14101
rect 4193 14045 4279 14101
rect 4335 14045 4421 14101
rect 4477 14045 4563 14101
rect 4619 14045 4705 14101
rect 4761 14045 4847 14101
rect 4903 14045 4989 14101
rect 5045 14045 5131 14101
rect 5187 14045 5273 14101
rect 5329 14045 5415 14101
rect 5471 14045 5557 14101
rect 5613 14045 5699 14101
rect 5755 14045 5841 14101
rect 5897 14045 5983 14101
rect 6039 14045 6125 14101
rect 6181 14045 6267 14101
rect 6323 14045 6409 14101
rect 6465 14045 6551 14101
rect 6607 14045 6693 14101
rect 6749 14045 6835 14101
rect 6891 14045 6977 14101
rect 7033 14045 7119 14101
rect 7175 14045 7261 14101
rect 7317 14045 7403 14101
rect 7459 14045 7545 14101
rect 7601 14045 7687 14101
rect 7743 14045 7829 14101
rect 7885 14045 7971 14101
rect 8027 14045 8113 14101
rect 8169 14045 8255 14101
rect 8311 14045 8397 14101
rect 8453 14045 8539 14101
rect 8595 14045 8681 14101
rect 8737 14045 8823 14101
rect 8879 14045 8965 14101
rect 9021 14045 9107 14101
rect 9163 14045 9249 14101
rect 9305 14045 9391 14101
rect 9447 14045 9533 14101
rect 9589 14045 9675 14101
rect 9731 14045 9817 14101
rect 9873 14045 9959 14101
rect 10015 14045 10101 14101
rect 10157 14045 10243 14101
rect 10299 14045 10385 14101
rect 10441 14045 10527 14101
rect 10583 14045 10669 14101
rect 10725 14045 10811 14101
rect 10867 14045 10953 14101
rect 11009 14045 11095 14101
rect 11151 14045 11237 14101
rect 11293 14045 11379 14101
rect 11435 14045 11521 14101
rect 11577 14045 11663 14101
rect 11719 14045 11805 14101
rect 11861 14045 11947 14101
rect 12003 14045 12089 14101
rect 12145 14045 12231 14101
rect 12287 14045 12373 14101
rect 12429 14045 12515 14101
rect 12571 14045 12657 14101
rect 12713 14045 12799 14101
rect 12855 14045 12941 14101
rect 12997 14045 13083 14101
rect 13139 14045 13225 14101
rect 13281 14045 13367 14101
rect 13423 14045 13509 14101
rect 13565 14045 13651 14101
rect 13707 14045 13793 14101
rect 13849 14045 13935 14101
rect 13991 14045 14077 14101
rect 14133 14045 14219 14101
rect 14275 14045 14361 14101
rect 14417 14045 14503 14101
rect 14559 14045 14645 14101
rect 14701 14045 14787 14101
rect 14843 14045 14853 14101
rect 151 14035 14853 14045
<< via3 >>
rect 161 69581 217 69637
rect 303 69581 359 69637
rect 445 69581 501 69637
rect 587 69581 643 69637
rect 729 69581 785 69637
rect 871 69581 927 69637
rect 1013 69581 1069 69637
rect 1155 69581 1211 69637
rect 1297 69581 1353 69637
rect 1439 69581 1495 69637
rect 1581 69581 1637 69637
rect 1723 69581 1779 69637
rect 1865 69581 1921 69637
rect 2007 69581 2063 69637
rect 2149 69581 2205 69637
rect 2291 69581 2347 69637
rect 2433 69581 2489 69637
rect 2575 69581 2631 69637
rect 2717 69581 2773 69637
rect 2859 69581 2915 69637
rect 3001 69581 3057 69637
rect 3143 69581 3199 69637
rect 3285 69581 3341 69637
rect 3427 69581 3483 69637
rect 3569 69581 3625 69637
rect 3711 69581 3767 69637
rect 3853 69581 3909 69637
rect 3995 69581 4051 69637
rect 4137 69581 4193 69637
rect 4279 69581 4335 69637
rect 4421 69581 4477 69637
rect 4563 69581 4619 69637
rect 4705 69581 4761 69637
rect 4847 69581 4903 69637
rect 4989 69581 5045 69637
rect 5131 69581 5187 69637
rect 5273 69581 5329 69637
rect 5415 69581 5471 69637
rect 5557 69581 5613 69637
rect 5699 69581 5755 69637
rect 5841 69581 5897 69637
rect 5983 69581 6039 69637
rect 6125 69581 6181 69637
rect 6267 69581 6323 69637
rect 6409 69581 6465 69637
rect 6551 69581 6607 69637
rect 6693 69581 6749 69637
rect 6835 69581 6891 69637
rect 6977 69581 7033 69637
rect 7119 69581 7175 69637
rect 7261 69581 7317 69637
rect 7403 69581 7459 69637
rect 7545 69581 7601 69637
rect 7687 69581 7743 69637
rect 7829 69581 7885 69637
rect 7971 69581 8027 69637
rect 8113 69581 8169 69637
rect 8255 69581 8311 69637
rect 8397 69581 8453 69637
rect 8539 69581 8595 69637
rect 8681 69581 8737 69637
rect 8823 69581 8879 69637
rect 8965 69581 9021 69637
rect 9107 69581 9163 69637
rect 9249 69581 9305 69637
rect 9391 69581 9447 69637
rect 9533 69581 9589 69637
rect 9675 69581 9731 69637
rect 9817 69581 9873 69637
rect 9959 69581 10015 69637
rect 10101 69581 10157 69637
rect 10243 69581 10299 69637
rect 10385 69581 10441 69637
rect 10527 69581 10583 69637
rect 10669 69581 10725 69637
rect 10811 69581 10867 69637
rect 10953 69581 11009 69637
rect 11095 69581 11151 69637
rect 11237 69581 11293 69637
rect 11379 69581 11435 69637
rect 11521 69581 11577 69637
rect 11663 69581 11719 69637
rect 11805 69581 11861 69637
rect 11947 69581 12003 69637
rect 12089 69581 12145 69637
rect 12231 69581 12287 69637
rect 12373 69581 12429 69637
rect 12515 69581 12571 69637
rect 12657 69581 12713 69637
rect 12799 69581 12855 69637
rect 12941 69581 12997 69637
rect 13083 69581 13139 69637
rect 13225 69581 13281 69637
rect 13367 69581 13423 69637
rect 13509 69581 13565 69637
rect 13651 69581 13707 69637
rect 13793 69581 13849 69637
rect 13935 69581 13991 69637
rect 14077 69581 14133 69637
rect 14219 69581 14275 69637
rect 14361 69581 14417 69637
rect 14503 69581 14559 69637
rect 14645 69581 14701 69637
rect 14787 69581 14843 69637
rect 161 69439 217 69495
rect 303 69439 359 69495
rect 445 69439 501 69495
rect 587 69439 643 69495
rect 729 69439 785 69495
rect 871 69439 927 69495
rect 1013 69439 1069 69495
rect 1155 69439 1211 69495
rect 1297 69439 1353 69495
rect 1439 69439 1495 69495
rect 1581 69439 1637 69495
rect 1723 69439 1779 69495
rect 1865 69439 1921 69495
rect 2007 69439 2063 69495
rect 2149 69439 2205 69495
rect 2291 69439 2347 69495
rect 2433 69439 2489 69495
rect 2575 69439 2631 69495
rect 2717 69439 2773 69495
rect 2859 69439 2915 69495
rect 3001 69439 3057 69495
rect 3143 69439 3199 69495
rect 3285 69439 3341 69495
rect 3427 69439 3483 69495
rect 3569 69439 3625 69495
rect 3711 69439 3767 69495
rect 3853 69439 3909 69495
rect 3995 69439 4051 69495
rect 4137 69439 4193 69495
rect 4279 69439 4335 69495
rect 4421 69439 4477 69495
rect 4563 69439 4619 69495
rect 4705 69439 4761 69495
rect 4847 69439 4903 69495
rect 4989 69439 5045 69495
rect 5131 69439 5187 69495
rect 5273 69439 5329 69495
rect 5415 69439 5471 69495
rect 5557 69439 5613 69495
rect 5699 69439 5755 69495
rect 5841 69439 5897 69495
rect 5983 69439 6039 69495
rect 6125 69439 6181 69495
rect 6267 69439 6323 69495
rect 6409 69439 6465 69495
rect 6551 69439 6607 69495
rect 6693 69439 6749 69495
rect 6835 69439 6891 69495
rect 6977 69439 7033 69495
rect 7119 69439 7175 69495
rect 7261 69439 7317 69495
rect 7403 69439 7459 69495
rect 7545 69439 7601 69495
rect 7687 69439 7743 69495
rect 7829 69439 7885 69495
rect 7971 69439 8027 69495
rect 8113 69439 8169 69495
rect 8255 69439 8311 69495
rect 8397 69439 8453 69495
rect 8539 69439 8595 69495
rect 8681 69439 8737 69495
rect 8823 69439 8879 69495
rect 8965 69439 9021 69495
rect 9107 69439 9163 69495
rect 9249 69439 9305 69495
rect 9391 69439 9447 69495
rect 9533 69439 9589 69495
rect 9675 69439 9731 69495
rect 9817 69439 9873 69495
rect 9959 69439 10015 69495
rect 10101 69439 10157 69495
rect 10243 69439 10299 69495
rect 10385 69439 10441 69495
rect 10527 69439 10583 69495
rect 10669 69439 10725 69495
rect 10811 69439 10867 69495
rect 10953 69439 11009 69495
rect 11095 69439 11151 69495
rect 11237 69439 11293 69495
rect 11379 69439 11435 69495
rect 11521 69439 11577 69495
rect 11663 69439 11719 69495
rect 11805 69439 11861 69495
rect 11947 69439 12003 69495
rect 12089 69439 12145 69495
rect 12231 69439 12287 69495
rect 12373 69439 12429 69495
rect 12515 69439 12571 69495
rect 12657 69439 12713 69495
rect 12799 69439 12855 69495
rect 12941 69439 12997 69495
rect 13083 69439 13139 69495
rect 13225 69439 13281 69495
rect 13367 69439 13423 69495
rect 13509 69439 13565 69495
rect 13651 69439 13707 69495
rect 13793 69439 13849 69495
rect 13935 69439 13991 69495
rect 14077 69439 14133 69495
rect 14219 69439 14275 69495
rect 14361 69439 14417 69495
rect 14503 69439 14559 69495
rect 14645 69439 14701 69495
rect 14787 69439 14843 69495
rect 161 69297 217 69353
rect 303 69297 359 69353
rect 445 69297 501 69353
rect 587 69297 643 69353
rect 729 69297 785 69353
rect 871 69297 927 69353
rect 1013 69297 1069 69353
rect 1155 69297 1211 69353
rect 1297 69297 1353 69353
rect 1439 69297 1495 69353
rect 1581 69297 1637 69353
rect 1723 69297 1779 69353
rect 1865 69297 1921 69353
rect 2007 69297 2063 69353
rect 2149 69297 2205 69353
rect 2291 69297 2347 69353
rect 2433 69297 2489 69353
rect 2575 69297 2631 69353
rect 2717 69297 2773 69353
rect 2859 69297 2915 69353
rect 3001 69297 3057 69353
rect 3143 69297 3199 69353
rect 3285 69297 3341 69353
rect 3427 69297 3483 69353
rect 3569 69297 3625 69353
rect 3711 69297 3767 69353
rect 3853 69297 3909 69353
rect 3995 69297 4051 69353
rect 4137 69297 4193 69353
rect 4279 69297 4335 69353
rect 4421 69297 4477 69353
rect 4563 69297 4619 69353
rect 4705 69297 4761 69353
rect 4847 69297 4903 69353
rect 4989 69297 5045 69353
rect 5131 69297 5187 69353
rect 5273 69297 5329 69353
rect 5415 69297 5471 69353
rect 5557 69297 5613 69353
rect 5699 69297 5755 69353
rect 5841 69297 5897 69353
rect 5983 69297 6039 69353
rect 6125 69297 6181 69353
rect 6267 69297 6323 69353
rect 6409 69297 6465 69353
rect 6551 69297 6607 69353
rect 6693 69297 6749 69353
rect 6835 69297 6891 69353
rect 6977 69297 7033 69353
rect 7119 69297 7175 69353
rect 7261 69297 7317 69353
rect 7403 69297 7459 69353
rect 7545 69297 7601 69353
rect 7687 69297 7743 69353
rect 7829 69297 7885 69353
rect 7971 69297 8027 69353
rect 8113 69297 8169 69353
rect 8255 69297 8311 69353
rect 8397 69297 8453 69353
rect 8539 69297 8595 69353
rect 8681 69297 8737 69353
rect 8823 69297 8879 69353
rect 8965 69297 9021 69353
rect 9107 69297 9163 69353
rect 9249 69297 9305 69353
rect 9391 69297 9447 69353
rect 9533 69297 9589 69353
rect 9675 69297 9731 69353
rect 9817 69297 9873 69353
rect 9959 69297 10015 69353
rect 10101 69297 10157 69353
rect 10243 69297 10299 69353
rect 10385 69297 10441 69353
rect 10527 69297 10583 69353
rect 10669 69297 10725 69353
rect 10811 69297 10867 69353
rect 10953 69297 11009 69353
rect 11095 69297 11151 69353
rect 11237 69297 11293 69353
rect 11379 69297 11435 69353
rect 11521 69297 11577 69353
rect 11663 69297 11719 69353
rect 11805 69297 11861 69353
rect 11947 69297 12003 69353
rect 12089 69297 12145 69353
rect 12231 69297 12287 69353
rect 12373 69297 12429 69353
rect 12515 69297 12571 69353
rect 12657 69297 12713 69353
rect 12799 69297 12855 69353
rect 12941 69297 12997 69353
rect 13083 69297 13139 69353
rect 13225 69297 13281 69353
rect 13367 69297 13423 69353
rect 13509 69297 13565 69353
rect 13651 69297 13707 69353
rect 13793 69297 13849 69353
rect 13935 69297 13991 69353
rect 14077 69297 14133 69353
rect 14219 69297 14275 69353
rect 14361 69297 14417 69353
rect 14503 69297 14559 69353
rect 14645 69297 14701 69353
rect 14787 69297 14843 69353
rect 161 69155 217 69211
rect 303 69155 359 69211
rect 445 69155 501 69211
rect 587 69155 643 69211
rect 729 69155 785 69211
rect 871 69155 927 69211
rect 1013 69155 1069 69211
rect 1155 69155 1211 69211
rect 1297 69155 1353 69211
rect 1439 69155 1495 69211
rect 1581 69155 1637 69211
rect 1723 69155 1779 69211
rect 1865 69155 1921 69211
rect 2007 69155 2063 69211
rect 2149 69155 2205 69211
rect 2291 69155 2347 69211
rect 2433 69155 2489 69211
rect 2575 69155 2631 69211
rect 2717 69155 2773 69211
rect 2859 69155 2915 69211
rect 3001 69155 3057 69211
rect 3143 69155 3199 69211
rect 3285 69155 3341 69211
rect 3427 69155 3483 69211
rect 3569 69155 3625 69211
rect 3711 69155 3767 69211
rect 3853 69155 3909 69211
rect 3995 69155 4051 69211
rect 4137 69155 4193 69211
rect 4279 69155 4335 69211
rect 4421 69155 4477 69211
rect 4563 69155 4619 69211
rect 4705 69155 4761 69211
rect 4847 69155 4903 69211
rect 4989 69155 5045 69211
rect 5131 69155 5187 69211
rect 5273 69155 5329 69211
rect 5415 69155 5471 69211
rect 5557 69155 5613 69211
rect 5699 69155 5755 69211
rect 5841 69155 5897 69211
rect 5983 69155 6039 69211
rect 6125 69155 6181 69211
rect 6267 69155 6323 69211
rect 6409 69155 6465 69211
rect 6551 69155 6607 69211
rect 6693 69155 6749 69211
rect 6835 69155 6891 69211
rect 6977 69155 7033 69211
rect 7119 69155 7175 69211
rect 7261 69155 7317 69211
rect 7403 69155 7459 69211
rect 7545 69155 7601 69211
rect 7687 69155 7743 69211
rect 7829 69155 7885 69211
rect 7971 69155 8027 69211
rect 8113 69155 8169 69211
rect 8255 69155 8311 69211
rect 8397 69155 8453 69211
rect 8539 69155 8595 69211
rect 8681 69155 8737 69211
rect 8823 69155 8879 69211
rect 8965 69155 9021 69211
rect 9107 69155 9163 69211
rect 9249 69155 9305 69211
rect 9391 69155 9447 69211
rect 9533 69155 9589 69211
rect 9675 69155 9731 69211
rect 9817 69155 9873 69211
rect 9959 69155 10015 69211
rect 10101 69155 10157 69211
rect 10243 69155 10299 69211
rect 10385 69155 10441 69211
rect 10527 69155 10583 69211
rect 10669 69155 10725 69211
rect 10811 69155 10867 69211
rect 10953 69155 11009 69211
rect 11095 69155 11151 69211
rect 11237 69155 11293 69211
rect 11379 69155 11435 69211
rect 11521 69155 11577 69211
rect 11663 69155 11719 69211
rect 11805 69155 11861 69211
rect 11947 69155 12003 69211
rect 12089 69155 12145 69211
rect 12231 69155 12287 69211
rect 12373 69155 12429 69211
rect 12515 69155 12571 69211
rect 12657 69155 12713 69211
rect 12799 69155 12855 69211
rect 12941 69155 12997 69211
rect 13083 69155 13139 69211
rect 13225 69155 13281 69211
rect 13367 69155 13423 69211
rect 13509 69155 13565 69211
rect 13651 69155 13707 69211
rect 13793 69155 13849 69211
rect 13935 69155 13991 69211
rect 14077 69155 14133 69211
rect 14219 69155 14275 69211
rect 14361 69155 14417 69211
rect 14503 69155 14559 69211
rect 14645 69155 14701 69211
rect 14787 69155 14843 69211
rect 161 69013 217 69069
rect 303 69013 359 69069
rect 445 69013 501 69069
rect 587 69013 643 69069
rect 729 69013 785 69069
rect 871 69013 927 69069
rect 1013 69013 1069 69069
rect 1155 69013 1211 69069
rect 1297 69013 1353 69069
rect 1439 69013 1495 69069
rect 1581 69013 1637 69069
rect 1723 69013 1779 69069
rect 1865 69013 1921 69069
rect 2007 69013 2063 69069
rect 2149 69013 2205 69069
rect 2291 69013 2347 69069
rect 2433 69013 2489 69069
rect 2575 69013 2631 69069
rect 2717 69013 2773 69069
rect 2859 69013 2915 69069
rect 3001 69013 3057 69069
rect 3143 69013 3199 69069
rect 3285 69013 3341 69069
rect 3427 69013 3483 69069
rect 3569 69013 3625 69069
rect 3711 69013 3767 69069
rect 3853 69013 3909 69069
rect 3995 69013 4051 69069
rect 4137 69013 4193 69069
rect 4279 69013 4335 69069
rect 4421 69013 4477 69069
rect 4563 69013 4619 69069
rect 4705 69013 4761 69069
rect 4847 69013 4903 69069
rect 4989 69013 5045 69069
rect 5131 69013 5187 69069
rect 5273 69013 5329 69069
rect 5415 69013 5471 69069
rect 5557 69013 5613 69069
rect 5699 69013 5755 69069
rect 5841 69013 5897 69069
rect 5983 69013 6039 69069
rect 6125 69013 6181 69069
rect 6267 69013 6323 69069
rect 6409 69013 6465 69069
rect 6551 69013 6607 69069
rect 6693 69013 6749 69069
rect 6835 69013 6891 69069
rect 6977 69013 7033 69069
rect 7119 69013 7175 69069
rect 7261 69013 7317 69069
rect 7403 69013 7459 69069
rect 7545 69013 7601 69069
rect 7687 69013 7743 69069
rect 7829 69013 7885 69069
rect 7971 69013 8027 69069
rect 8113 69013 8169 69069
rect 8255 69013 8311 69069
rect 8397 69013 8453 69069
rect 8539 69013 8595 69069
rect 8681 69013 8737 69069
rect 8823 69013 8879 69069
rect 8965 69013 9021 69069
rect 9107 69013 9163 69069
rect 9249 69013 9305 69069
rect 9391 69013 9447 69069
rect 9533 69013 9589 69069
rect 9675 69013 9731 69069
rect 9817 69013 9873 69069
rect 9959 69013 10015 69069
rect 10101 69013 10157 69069
rect 10243 69013 10299 69069
rect 10385 69013 10441 69069
rect 10527 69013 10583 69069
rect 10669 69013 10725 69069
rect 10811 69013 10867 69069
rect 10953 69013 11009 69069
rect 11095 69013 11151 69069
rect 11237 69013 11293 69069
rect 11379 69013 11435 69069
rect 11521 69013 11577 69069
rect 11663 69013 11719 69069
rect 11805 69013 11861 69069
rect 11947 69013 12003 69069
rect 12089 69013 12145 69069
rect 12231 69013 12287 69069
rect 12373 69013 12429 69069
rect 12515 69013 12571 69069
rect 12657 69013 12713 69069
rect 12799 69013 12855 69069
rect 12941 69013 12997 69069
rect 13083 69013 13139 69069
rect 13225 69013 13281 69069
rect 13367 69013 13423 69069
rect 13509 69013 13565 69069
rect 13651 69013 13707 69069
rect 13793 69013 13849 69069
rect 13935 69013 13991 69069
rect 14077 69013 14133 69069
rect 14219 69013 14275 69069
rect 14361 69013 14417 69069
rect 14503 69013 14559 69069
rect 14645 69013 14701 69069
rect 14787 69013 14843 69069
rect 161 68871 217 68927
rect 303 68871 359 68927
rect 445 68871 501 68927
rect 587 68871 643 68927
rect 729 68871 785 68927
rect 871 68871 927 68927
rect 1013 68871 1069 68927
rect 1155 68871 1211 68927
rect 1297 68871 1353 68927
rect 1439 68871 1495 68927
rect 1581 68871 1637 68927
rect 1723 68871 1779 68927
rect 1865 68871 1921 68927
rect 2007 68871 2063 68927
rect 2149 68871 2205 68927
rect 2291 68871 2347 68927
rect 2433 68871 2489 68927
rect 2575 68871 2631 68927
rect 2717 68871 2773 68927
rect 2859 68871 2915 68927
rect 3001 68871 3057 68927
rect 3143 68871 3199 68927
rect 3285 68871 3341 68927
rect 3427 68871 3483 68927
rect 3569 68871 3625 68927
rect 3711 68871 3767 68927
rect 3853 68871 3909 68927
rect 3995 68871 4051 68927
rect 4137 68871 4193 68927
rect 4279 68871 4335 68927
rect 4421 68871 4477 68927
rect 4563 68871 4619 68927
rect 4705 68871 4761 68927
rect 4847 68871 4903 68927
rect 4989 68871 5045 68927
rect 5131 68871 5187 68927
rect 5273 68871 5329 68927
rect 5415 68871 5471 68927
rect 5557 68871 5613 68927
rect 5699 68871 5755 68927
rect 5841 68871 5897 68927
rect 5983 68871 6039 68927
rect 6125 68871 6181 68927
rect 6267 68871 6323 68927
rect 6409 68871 6465 68927
rect 6551 68871 6607 68927
rect 6693 68871 6749 68927
rect 6835 68871 6891 68927
rect 6977 68871 7033 68927
rect 7119 68871 7175 68927
rect 7261 68871 7317 68927
rect 7403 68871 7459 68927
rect 7545 68871 7601 68927
rect 7687 68871 7743 68927
rect 7829 68871 7885 68927
rect 7971 68871 8027 68927
rect 8113 68871 8169 68927
rect 8255 68871 8311 68927
rect 8397 68871 8453 68927
rect 8539 68871 8595 68927
rect 8681 68871 8737 68927
rect 8823 68871 8879 68927
rect 8965 68871 9021 68927
rect 9107 68871 9163 68927
rect 9249 68871 9305 68927
rect 9391 68871 9447 68927
rect 9533 68871 9589 68927
rect 9675 68871 9731 68927
rect 9817 68871 9873 68927
rect 9959 68871 10015 68927
rect 10101 68871 10157 68927
rect 10243 68871 10299 68927
rect 10385 68871 10441 68927
rect 10527 68871 10583 68927
rect 10669 68871 10725 68927
rect 10811 68871 10867 68927
rect 10953 68871 11009 68927
rect 11095 68871 11151 68927
rect 11237 68871 11293 68927
rect 11379 68871 11435 68927
rect 11521 68871 11577 68927
rect 11663 68871 11719 68927
rect 11805 68871 11861 68927
rect 11947 68871 12003 68927
rect 12089 68871 12145 68927
rect 12231 68871 12287 68927
rect 12373 68871 12429 68927
rect 12515 68871 12571 68927
rect 12657 68871 12713 68927
rect 12799 68871 12855 68927
rect 12941 68871 12997 68927
rect 13083 68871 13139 68927
rect 13225 68871 13281 68927
rect 13367 68871 13423 68927
rect 13509 68871 13565 68927
rect 13651 68871 13707 68927
rect 13793 68871 13849 68927
rect 13935 68871 13991 68927
rect 14077 68871 14133 68927
rect 14219 68871 14275 68927
rect 14361 68871 14417 68927
rect 14503 68871 14559 68927
rect 14645 68871 14701 68927
rect 14787 68871 14843 68927
rect 161 68729 217 68785
rect 303 68729 359 68785
rect 445 68729 501 68785
rect 587 68729 643 68785
rect 729 68729 785 68785
rect 871 68729 927 68785
rect 1013 68729 1069 68785
rect 1155 68729 1211 68785
rect 1297 68729 1353 68785
rect 1439 68729 1495 68785
rect 1581 68729 1637 68785
rect 1723 68729 1779 68785
rect 1865 68729 1921 68785
rect 2007 68729 2063 68785
rect 2149 68729 2205 68785
rect 2291 68729 2347 68785
rect 2433 68729 2489 68785
rect 2575 68729 2631 68785
rect 2717 68729 2773 68785
rect 2859 68729 2915 68785
rect 3001 68729 3057 68785
rect 3143 68729 3199 68785
rect 3285 68729 3341 68785
rect 3427 68729 3483 68785
rect 3569 68729 3625 68785
rect 3711 68729 3767 68785
rect 3853 68729 3909 68785
rect 3995 68729 4051 68785
rect 4137 68729 4193 68785
rect 4279 68729 4335 68785
rect 4421 68729 4477 68785
rect 4563 68729 4619 68785
rect 4705 68729 4761 68785
rect 4847 68729 4903 68785
rect 4989 68729 5045 68785
rect 5131 68729 5187 68785
rect 5273 68729 5329 68785
rect 5415 68729 5471 68785
rect 5557 68729 5613 68785
rect 5699 68729 5755 68785
rect 5841 68729 5897 68785
rect 5983 68729 6039 68785
rect 6125 68729 6181 68785
rect 6267 68729 6323 68785
rect 6409 68729 6465 68785
rect 6551 68729 6607 68785
rect 6693 68729 6749 68785
rect 6835 68729 6891 68785
rect 6977 68729 7033 68785
rect 7119 68729 7175 68785
rect 7261 68729 7317 68785
rect 7403 68729 7459 68785
rect 7545 68729 7601 68785
rect 7687 68729 7743 68785
rect 7829 68729 7885 68785
rect 7971 68729 8027 68785
rect 8113 68729 8169 68785
rect 8255 68729 8311 68785
rect 8397 68729 8453 68785
rect 8539 68729 8595 68785
rect 8681 68729 8737 68785
rect 8823 68729 8879 68785
rect 8965 68729 9021 68785
rect 9107 68729 9163 68785
rect 9249 68729 9305 68785
rect 9391 68729 9447 68785
rect 9533 68729 9589 68785
rect 9675 68729 9731 68785
rect 9817 68729 9873 68785
rect 9959 68729 10015 68785
rect 10101 68729 10157 68785
rect 10243 68729 10299 68785
rect 10385 68729 10441 68785
rect 10527 68729 10583 68785
rect 10669 68729 10725 68785
rect 10811 68729 10867 68785
rect 10953 68729 11009 68785
rect 11095 68729 11151 68785
rect 11237 68729 11293 68785
rect 11379 68729 11435 68785
rect 11521 68729 11577 68785
rect 11663 68729 11719 68785
rect 11805 68729 11861 68785
rect 11947 68729 12003 68785
rect 12089 68729 12145 68785
rect 12231 68729 12287 68785
rect 12373 68729 12429 68785
rect 12515 68729 12571 68785
rect 12657 68729 12713 68785
rect 12799 68729 12855 68785
rect 12941 68729 12997 68785
rect 13083 68729 13139 68785
rect 13225 68729 13281 68785
rect 13367 68729 13423 68785
rect 13509 68729 13565 68785
rect 13651 68729 13707 68785
rect 13793 68729 13849 68785
rect 13935 68729 13991 68785
rect 14077 68729 14133 68785
rect 14219 68729 14275 68785
rect 14361 68729 14417 68785
rect 14503 68729 14559 68785
rect 14645 68729 14701 68785
rect 14787 68729 14843 68785
rect 161 68587 217 68643
rect 303 68587 359 68643
rect 445 68587 501 68643
rect 587 68587 643 68643
rect 729 68587 785 68643
rect 871 68587 927 68643
rect 1013 68587 1069 68643
rect 1155 68587 1211 68643
rect 1297 68587 1353 68643
rect 1439 68587 1495 68643
rect 1581 68587 1637 68643
rect 1723 68587 1779 68643
rect 1865 68587 1921 68643
rect 2007 68587 2063 68643
rect 2149 68587 2205 68643
rect 2291 68587 2347 68643
rect 2433 68587 2489 68643
rect 2575 68587 2631 68643
rect 2717 68587 2773 68643
rect 2859 68587 2915 68643
rect 3001 68587 3057 68643
rect 3143 68587 3199 68643
rect 3285 68587 3341 68643
rect 3427 68587 3483 68643
rect 3569 68587 3625 68643
rect 3711 68587 3767 68643
rect 3853 68587 3909 68643
rect 3995 68587 4051 68643
rect 4137 68587 4193 68643
rect 4279 68587 4335 68643
rect 4421 68587 4477 68643
rect 4563 68587 4619 68643
rect 4705 68587 4761 68643
rect 4847 68587 4903 68643
rect 4989 68587 5045 68643
rect 5131 68587 5187 68643
rect 5273 68587 5329 68643
rect 5415 68587 5471 68643
rect 5557 68587 5613 68643
rect 5699 68587 5755 68643
rect 5841 68587 5897 68643
rect 5983 68587 6039 68643
rect 6125 68587 6181 68643
rect 6267 68587 6323 68643
rect 6409 68587 6465 68643
rect 6551 68587 6607 68643
rect 6693 68587 6749 68643
rect 6835 68587 6891 68643
rect 6977 68587 7033 68643
rect 7119 68587 7175 68643
rect 7261 68587 7317 68643
rect 7403 68587 7459 68643
rect 7545 68587 7601 68643
rect 7687 68587 7743 68643
rect 7829 68587 7885 68643
rect 7971 68587 8027 68643
rect 8113 68587 8169 68643
rect 8255 68587 8311 68643
rect 8397 68587 8453 68643
rect 8539 68587 8595 68643
rect 8681 68587 8737 68643
rect 8823 68587 8879 68643
rect 8965 68587 9021 68643
rect 9107 68587 9163 68643
rect 9249 68587 9305 68643
rect 9391 68587 9447 68643
rect 9533 68587 9589 68643
rect 9675 68587 9731 68643
rect 9817 68587 9873 68643
rect 9959 68587 10015 68643
rect 10101 68587 10157 68643
rect 10243 68587 10299 68643
rect 10385 68587 10441 68643
rect 10527 68587 10583 68643
rect 10669 68587 10725 68643
rect 10811 68587 10867 68643
rect 10953 68587 11009 68643
rect 11095 68587 11151 68643
rect 11237 68587 11293 68643
rect 11379 68587 11435 68643
rect 11521 68587 11577 68643
rect 11663 68587 11719 68643
rect 11805 68587 11861 68643
rect 11947 68587 12003 68643
rect 12089 68587 12145 68643
rect 12231 68587 12287 68643
rect 12373 68587 12429 68643
rect 12515 68587 12571 68643
rect 12657 68587 12713 68643
rect 12799 68587 12855 68643
rect 12941 68587 12997 68643
rect 13083 68587 13139 68643
rect 13225 68587 13281 68643
rect 13367 68587 13423 68643
rect 13509 68587 13565 68643
rect 13651 68587 13707 68643
rect 13793 68587 13849 68643
rect 13935 68587 13991 68643
rect 14077 68587 14133 68643
rect 14219 68587 14275 68643
rect 14361 68587 14417 68643
rect 14503 68587 14559 68643
rect 14645 68587 14701 68643
rect 14787 68587 14843 68643
rect 161 68445 217 68501
rect 303 68445 359 68501
rect 445 68445 501 68501
rect 587 68445 643 68501
rect 729 68445 785 68501
rect 871 68445 927 68501
rect 1013 68445 1069 68501
rect 1155 68445 1211 68501
rect 1297 68445 1353 68501
rect 1439 68445 1495 68501
rect 1581 68445 1637 68501
rect 1723 68445 1779 68501
rect 1865 68445 1921 68501
rect 2007 68445 2063 68501
rect 2149 68445 2205 68501
rect 2291 68445 2347 68501
rect 2433 68445 2489 68501
rect 2575 68445 2631 68501
rect 2717 68445 2773 68501
rect 2859 68445 2915 68501
rect 3001 68445 3057 68501
rect 3143 68445 3199 68501
rect 3285 68445 3341 68501
rect 3427 68445 3483 68501
rect 3569 68445 3625 68501
rect 3711 68445 3767 68501
rect 3853 68445 3909 68501
rect 3995 68445 4051 68501
rect 4137 68445 4193 68501
rect 4279 68445 4335 68501
rect 4421 68445 4477 68501
rect 4563 68445 4619 68501
rect 4705 68445 4761 68501
rect 4847 68445 4903 68501
rect 4989 68445 5045 68501
rect 5131 68445 5187 68501
rect 5273 68445 5329 68501
rect 5415 68445 5471 68501
rect 5557 68445 5613 68501
rect 5699 68445 5755 68501
rect 5841 68445 5897 68501
rect 5983 68445 6039 68501
rect 6125 68445 6181 68501
rect 6267 68445 6323 68501
rect 6409 68445 6465 68501
rect 6551 68445 6607 68501
rect 6693 68445 6749 68501
rect 6835 68445 6891 68501
rect 6977 68445 7033 68501
rect 7119 68445 7175 68501
rect 7261 68445 7317 68501
rect 7403 68445 7459 68501
rect 7545 68445 7601 68501
rect 7687 68445 7743 68501
rect 7829 68445 7885 68501
rect 7971 68445 8027 68501
rect 8113 68445 8169 68501
rect 8255 68445 8311 68501
rect 8397 68445 8453 68501
rect 8539 68445 8595 68501
rect 8681 68445 8737 68501
rect 8823 68445 8879 68501
rect 8965 68445 9021 68501
rect 9107 68445 9163 68501
rect 9249 68445 9305 68501
rect 9391 68445 9447 68501
rect 9533 68445 9589 68501
rect 9675 68445 9731 68501
rect 9817 68445 9873 68501
rect 9959 68445 10015 68501
rect 10101 68445 10157 68501
rect 10243 68445 10299 68501
rect 10385 68445 10441 68501
rect 10527 68445 10583 68501
rect 10669 68445 10725 68501
rect 10811 68445 10867 68501
rect 10953 68445 11009 68501
rect 11095 68445 11151 68501
rect 11237 68445 11293 68501
rect 11379 68445 11435 68501
rect 11521 68445 11577 68501
rect 11663 68445 11719 68501
rect 11805 68445 11861 68501
rect 11947 68445 12003 68501
rect 12089 68445 12145 68501
rect 12231 68445 12287 68501
rect 12373 68445 12429 68501
rect 12515 68445 12571 68501
rect 12657 68445 12713 68501
rect 12799 68445 12855 68501
rect 12941 68445 12997 68501
rect 13083 68445 13139 68501
rect 13225 68445 13281 68501
rect 13367 68445 13423 68501
rect 13509 68445 13565 68501
rect 13651 68445 13707 68501
rect 13793 68445 13849 68501
rect 13935 68445 13991 68501
rect 14077 68445 14133 68501
rect 14219 68445 14275 68501
rect 14361 68445 14417 68501
rect 14503 68445 14559 68501
rect 14645 68445 14701 68501
rect 14787 68445 14843 68501
rect 161 68115 217 68171
rect 303 68115 359 68171
rect 445 68115 501 68171
rect 587 68115 643 68171
rect 729 68115 785 68171
rect 871 68115 927 68171
rect 1013 68115 1069 68171
rect 1155 68115 1211 68171
rect 1297 68115 1353 68171
rect 1439 68115 1495 68171
rect 1581 68115 1637 68171
rect 1723 68115 1779 68171
rect 1865 68115 1921 68171
rect 2007 68115 2063 68171
rect 2149 68115 2205 68171
rect 2291 68115 2347 68171
rect 2433 68115 2489 68171
rect 2575 68115 2631 68171
rect 2717 68115 2773 68171
rect 2859 68115 2915 68171
rect 3001 68115 3057 68171
rect 3143 68115 3199 68171
rect 3285 68115 3341 68171
rect 3427 68115 3483 68171
rect 3569 68115 3625 68171
rect 3711 68115 3767 68171
rect 3853 68115 3909 68171
rect 3995 68115 4051 68171
rect 4137 68115 4193 68171
rect 4279 68115 4335 68171
rect 4421 68115 4477 68171
rect 4563 68115 4619 68171
rect 4705 68115 4761 68171
rect 4847 68115 4903 68171
rect 4989 68115 5045 68171
rect 5131 68115 5187 68171
rect 5273 68115 5329 68171
rect 5415 68115 5471 68171
rect 5557 68115 5613 68171
rect 5699 68115 5755 68171
rect 5841 68115 5897 68171
rect 5983 68115 6039 68171
rect 6125 68115 6181 68171
rect 6267 68115 6323 68171
rect 6409 68115 6465 68171
rect 6551 68115 6607 68171
rect 6693 68115 6749 68171
rect 6835 68115 6891 68171
rect 6977 68115 7033 68171
rect 7119 68115 7175 68171
rect 7261 68115 7317 68171
rect 7403 68115 7459 68171
rect 7545 68115 7601 68171
rect 7687 68115 7743 68171
rect 7829 68115 7885 68171
rect 7971 68115 8027 68171
rect 8113 68115 8169 68171
rect 8255 68115 8311 68171
rect 8397 68115 8453 68171
rect 8539 68115 8595 68171
rect 8681 68115 8737 68171
rect 8823 68115 8879 68171
rect 8965 68115 9021 68171
rect 9107 68115 9163 68171
rect 9249 68115 9305 68171
rect 9391 68115 9447 68171
rect 9533 68115 9589 68171
rect 9675 68115 9731 68171
rect 9817 68115 9873 68171
rect 9959 68115 10015 68171
rect 10101 68115 10157 68171
rect 10243 68115 10299 68171
rect 10385 68115 10441 68171
rect 10527 68115 10583 68171
rect 10669 68115 10725 68171
rect 10811 68115 10867 68171
rect 10953 68115 11009 68171
rect 11095 68115 11151 68171
rect 11237 68115 11293 68171
rect 11379 68115 11435 68171
rect 11521 68115 11577 68171
rect 11663 68115 11719 68171
rect 11805 68115 11861 68171
rect 11947 68115 12003 68171
rect 12089 68115 12145 68171
rect 12231 68115 12287 68171
rect 12373 68115 12429 68171
rect 12515 68115 12571 68171
rect 12657 68115 12713 68171
rect 12799 68115 12855 68171
rect 12941 68115 12997 68171
rect 13083 68115 13139 68171
rect 13225 68115 13281 68171
rect 13367 68115 13423 68171
rect 13509 68115 13565 68171
rect 13651 68115 13707 68171
rect 13793 68115 13849 68171
rect 13935 68115 13991 68171
rect 14077 68115 14133 68171
rect 14219 68115 14275 68171
rect 14361 68115 14417 68171
rect 14503 68115 14559 68171
rect 14645 68115 14701 68171
rect 14787 68115 14843 68171
rect 161 67973 217 68029
rect 303 67973 359 68029
rect 445 67973 501 68029
rect 587 67973 643 68029
rect 729 67973 785 68029
rect 871 67973 927 68029
rect 1013 67973 1069 68029
rect 1155 67973 1211 68029
rect 1297 67973 1353 68029
rect 1439 67973 1495 68029
rect 1581 67973 1637 68029
rect 1723 67973 1779 68029
rect 1865 67973 1921 68029
rect 2007 67973 2063 68029
rect 2149 67973 2205 68029
rect 2291 67973 2347 68029
rect 2433 67973 2489 68029
rect 2575 67973 2631 68029
rect 2717 67973 2773 68029
rect 2859 67973 2915 68029
rect 3001 67973 3057 68029
rect 3143 67973 3199 68029
rect 3285 67973 3341 68029
rect 3427 67973 3483 68029
rect 3569 67973 3625 68029
rect 3711 67973 3767 68029
rect 3853 67973 3909 68029
rect 3995 67973 4051 68029
rect 4137 67973 4193 68029
rect 4279 67973 4335 68029
rect 4421 67973 4477 68029
rect 4563 67973 4619 68029
rect 4705 67973 4761 68029
rect 4847 67973 4903 68029
rect 4989 67973 5045 68029
rect 5131 67973 5187 68029
rect 5273 67973 5329 68029
rect 5415 67973 5471 68029
rect 5557 67973 5613 68029
rect 5699 67973 5755 68029
rect 5841 67973 5897 68029
rect 5983 67973 6039 68029
rect 6125 67973 6181 68029
rect 6267 67973 6323 68029
rect 6409 67973 6465 68029
rect 6551 67973 6607 68029
rect 6693 67973 6749 68029
rect 6835 67973 6891 68029
rect 6977 67973 7033 68029
rect 7119 67973 7175 68029
rect 7261 67973 7317 68029
rect 7403 67973 7459 68029
rect 7545 67973 7601 68029
rect 7687 67973 7743 68029
rect 7829 67973 7885 68029
rect 7971 67973 8027 68029
rect 8113 67973 8169 68029
rect 8255 67973 8311 68029
rect 8397 67973 8453 68029
rect 8539 67973 8595 68029
rect 8681 67973 8737 68029
rect 8823 67973 8879 68029
rect 8965 67973 9021 68029
rect 9107 67973 9163 68029
rect 9249 67973 9305 68029
rect 9391 67973 9447 68029
rect 9533 67973 9589 68029
rect 9675 67973 9731 68029
rect 9817 67973 9873 68029
rect 9959 67973 10015 68029
rect 10101 67973 10157 68029
rect 10243 67973 10299 68029
rect 10385 67973 10441 68029
rect 10527 67973 10583 68029
rect 10669 67973 10725 68029
rect 10811 67973 10867 68029
rect 10953 67973 11009 68029
rect 11095 67973 11151 68029
rect 11237 67973 11293 68029
rect 11379 67973 11435 68029
rect 11521 67973 11577 68029
rect 11663 67973 11719 68029
rect 11805 67973 11861 68029
rect 11947 67973 12003 68029
rect 12089 67973 12145 68029
rect 12231 67973 12287 68029
rect 12373 67973 12429 68029
rect 12515 67973 12571 68029
rect 12657 67973 12713 68029
rect 12799 67973 12855 68029
rect 12941 67973 12997 68029
rect 13083 67973 13139 68029
rect 13225 67973 13281 68029
rect 13367 67973 13423 68029
rect 13509 67973 13565 68029
rect 13651 67973 13707 68029
rect 13793 67973 13849 68029
rect 13935 67973 13991 68029
rect 14077 67973 14133 68029
rect 14219 67973 14275 68029
rect 14361 67973 14417 68029
rect 14503 67973 14559 68029
rect 14645 67973 14701 68029
rect 14787 67973 14843 68029
rect 161 67831 217 67887
rect 303 67831 359 67887
rect 445 67831 501 67887
rect 587 67831 643 67887
rect 729 67831 785 67887
rect 871 67831 927 67887
rect 1013 67831 1069 67887
rect 1155 67831 1211 67887
rect 1297 67831 1353 67887
rect 1439 67831 1495 67887
rect 1581 67831 1637 67887
rect 1723 67831 1779 67887
rect 1865 67831 1921 67887
rect 2007 67831 2063 67887
rect 2149 67831 2205 67887
rect 2291 67831 2347 67887
rect 2433 67831 2489 67887
rect 2575 67831 2631 67887
rect 2717 67831 2773 67887
rect 2859 67831 2915 67887
rect 3001 67831 3057 67887
rect 3143 67831 3199 67887
rect 3285 67831 3341 67887
rect 3427 67831 3483 67887
rect 3569 67831 3625 67887
rect 3711 67831 3767 67887
rect 3853 67831 3909 67887
rect 3995 67831 4051 67887
rect 4137 67831 4193 67887
rect 4279 67831 4335 67887
rect 4421 67831 4477 67887
rect 4563 67831 4619 67887
rect 4705 67831 4761 67887
rect 4847 67831 4903 67887
rect 4989 67831 5045 67887
rect 5131 67831 5187 67887
rect 5273 67831 5329 67887
rect 5415 67831 5471 67887
rect 5557 67831 5613 67887
rect 5699 67831 5755 67887
rect 5841 67831 5897 67887
rect 5983 67831 6039 67887
rect 6125 67831 6181 67887
rect 6267 67831 6323 67887
rect 6409 67831 6465 67887
rect 6551 67831 6607 67887
rect 6693 67831 6749 67887
rect 6835 67831 6891 67887
rect 6977 67831 7033 67887
rect 7119 67831 7175 67887
rect 7261 67831 7317 67887
rect 7403 67831 7459 67887
rect 7545 67831 7601 67887
rect 7687 67831 7743 67887
rect 7829 67831 7885 67887
rect 7971 67831 8027 67887
rect 8113 67831 8169 67887
rect 8255 67831 8311 67887
rect 8397 67831 8453 67887
rect 8539 67831 8595 67887
rect 8681 67831 8737 67887
rect 8823 67831 8879 67887
rect 8965 67831 9021 67887
rect 9107 67831 9163 67887
rect 9249 67831 9305 67887
rect 9391 67831 9447 67887
rect 9533 67831 9589 67887
rect 9675 67831 9731 67887
rect 9817 67831 9873 67887
rect 9959 67831 10015 67887
rect 10101 67831 10157 67887
rect 10243 67831 10299 67887
rect 10385 67831 10441 67887
rect 10527 67831 10583 67887
rect 10669 67831 10725 67887
rect 10811 67831 10867 67887
rect 10953 67831 11009 67887
rect 11095 67831 11151 67887
rect 11237 67831 11293 67887
rect 11379 67831 11435 67887
rect 11521 67831 11577 67887
rect 11663 67831 11719 67887
rect 11805 67831 11861 67887
rect 11947 67831 12003 67887
rect 12089 67831 12145 67887
rect 12231 67831 12287 67887
rect 12373 67831 12429 67887
rect 12515 67831 12571 67887
rect 12657 67831 12713 67887
rect 12799 67831 12855 67887
rect 12941 67831 12997 67887
rect 13083 67831 13139 67887
rect 13225 67831 13281 67887
rect 13367 67831 13423 67887
rect 13509 67831 13565 67887
rect 13651 67831 13707 67887
rect 13793 67831 13849 67887
rect 13935 67831 13991 67887
rect 14077 67831 14133 67887
rect 14219 67831 14275 67887
rect 14361 67831 14417 67887
rect 14503 67831 14559 67887
rect 14645 67831 14701 67887
rect 14787 67831 14843 67887
rect 161 67689 217 67745
rect 303 67689 359 67745
rect 445 67689 501 67745
rect 587 67689 643 67745
rect 729 67689 785 67745
rect 871 67689 927 67745
rect 1013 67689 1069 67745
rect 1155 67689 1211 67745
rect 1297 67689 1353 67745
rect 1439 67689 1495 67745
rect 1581 67689 1637 67745
rect 1723 67689 1779 67745
rect 1865 67689 1921 67745
rect 2007 67689 2063 67745
rect 2149 67689 2205 67745
rect 2291 67689 2347 67745
rect 2433 67689 2489 67745
rect 2575 67689 2631 67745
rect 2717 67689 2773 67745
rect 2859 67689 2915 67745
rect 3001 67689 3057 67745
rect 3143 67689 3199 67745
rect 3285 67689 3341 67745
rect 3427 67689 3483 67745
rect 3569 67689 3625 67745
rect 3711 67689 3767 67745
rect 3853 67689 3909 67745
rect 3995 67689 4051 67745
rect 4137 67689 4193 67745
rect 4279 67689 4335 67745
rect 4421 67689 4477 67745
rect 4563 67689 4619 67745
rect 4705 67689 4761 67745
rect 4847 67689 4903 67745
rect 4989 67689 5045 67745
rect 5131 67689 5187 67745
rect 5273 67689 5329 67745
rect 5415 67689 5471 67745
rect 5557 67689 5613 67745
rect 5699 67689 5755 67745
rect 5841 67689 5897 67745
rect 5983 67689 6039 67745
rect 6125 67689 6181 67745
rect 6267 67689 6323 67745
rect 6409 67689 6465 67745
rect 6551 67689 6607 67745
rect 6693 67689 6749 67745
rect 6835 67689 6891 67745
rect 6977 67689 7033 67745
rect 7119 67689 7175 67745
rect 7261 67689 7317 67745
rect 7403 67689 7459 67745
rect 7545 67689 7601 67745
rect 7687 67689 7743 67745
rect 7829 67689 7885 67745
rect 7971 67689 8027 67745
rect 8113 67689 8169 67745
rect 8255 67689 8311 67745
rect 8397 67689 8453 67745
rect 8539 67689 8595 67745
rect 8681 67689 8737 67745
rect 8823 67689 8879 67745
rect 8965 67689 9021 67745
rect 9107 67689 9163 67745
rect 9249 67689 9305 67745
rect 9391 67689 9447 67745
rect 9533 67689 9589 67745
rect 9675 67689 9731 67745
rect 9817 67689 9873 67745
rect 9959 67689 10015 67745
rect 10101 67689 10157 67745
rect 10243 67689 10299 67745
rect 10385 67689 10441 67745
rect 10527 67689 10583 67745
rect 10669 67689 10725 67745
rect 10811 67689 10867 67745
rect 10953 67689 11009 67745
rect 11095 67689 11151 67745
rect 11237 67689 11293 67745
rect 11379 67689 11435 67745
rect 11521 67689 11577 67745
rect 11663 67689 11719 67745
rect 11805 67689 11861 67745
rect 11947 67689 12003 67745
rect 12089 67689 12145 67745
rect 12231 67689 12287 67745
rect 12373 67689 12429 67745
rect 12515 67689 12571 67745
rect 12657 67689 12713 67745
rect 12799 67689 12855 67745
rect 12941 67689 12997 67745
rect 13083 67689 13139 67745
rect 13225 67689 13281 67745
rect 13367 67689 13423 67745
rect 13509 67689 13565 67745
rect 13651 67689 13707 67745
rect 13793 67689 13849 67745
rect 13935 67689 13991 67745
rect 14077 67689 14133 67745
rect 14219 67689 14275 67745
rect 14361 67689 14417 67745
rect 14503 67689 14559 67745
rect 14645 67689 14701 67745
rect 14787 67689 14843 67745
rect 161 67547 217 67603
rect 303 67547 359 67603
rect 445 67547 501 67603
rect 587 67547 643 67603
rect 729 67547 785 67603
rect 871 67547 927 67603
rect 1013 67547 1069 67603
rect 1155 67547 1211 67603
rect 1297 67547 1353 67603
rect 1439 67547 1495 67603
rect 1581 67547 1637 67603
rect 1723 67547 1779 67603
rect 1865 67547 1921 67603
rect 2007 67547 2063 67603
rect 2149 67547 2205 67603
rect 2291 67547 2347 67603
rect 2433 67547 2489 67603
rect 2575 67547 2631 67603
rect 2717 67547 2773 67603
rect 2859 67547 2915 67603
rect 3001 67547 3057 67603
rect 3143 67547 3199 67603
rect 3285 67547 3341 67603
rect 3427 67547 3483 67603
rect 3569 67547 3625 67603
rect 3711 67547 3767 67603
rect 3853 67547 3909 67603
rect 3995 67547 4051 67603
rect 4137 67547 4193 67603
rect 4279 67547 4335 67603
rect 4421 67547 4477 67603
rect 4563 67547 4619 67603
rect 4705 67547 4761 67603
rect 4847 67547 4903 67603
rect 4989 67547 5045 67603
rect 5131 67547 5187 67603
rect 5273 67547 5329 67603
rect 5415 67547 5471 67603
rect 5557 67547 5613 67603
rect 5699 67547 5755 67603
rect 5841 67547 5897 67603
rect 5983 67547 6039 67603
rect 6125 67547 6181 67603
rect 6267 67547 6323 67603
rect 6409 67547 6465 67603
rect 6551 67547 6607 67603
rect 6693 67547 6749 67603
rect 6835 67547 6891 67603
rect 6977 67547 7033 67603
rect 7119 67547 7175 67603
rect 7261 67547 7317 67603
rect 7403 67547 7459 67603
rect 7545 67547 7601 67603
rect 7687 67547 7743 67603
rect 7829 67547 7885 67603
rect 7971 67547 8027 67603
rect 8113 67547 8169 67603
rect 8255 67547 8311 67603
rect 8397 67547 8453 67603
rect 8539 67547 8595 67603
rect 8681 67547 8737 67603
rect 8823 67547 8879 67603
rect 8965 67547 9021 67603
rect 9107 67547 9163 67603
rect 9249 67547 9305 67603
rect 9391 67547 9447 67603
rect 9533 67547 9589 67603
rect 9675 67547 9731 67603
rect 9817 67547 9873 67603
rect 9959 67547 10015 67603
rect 10101 67547 10157 67603
rect 10243 67547 10299 67603
rect 10385 67547 10441 67603
rect 10527 67547 10583 67603
rect 10669 67547 10725 67603
rect 10811 67547 10867 67603
rect 10953 67547 11009 67603
rect 11095 67547 11151 67603
rect 11237 67547 11293 67603
rect 11379 67547 11435 67603
rect 11521 67547 11577 67603
rect 11663 67547 11719 67603
rect 11805 67547 11861 67603
rect 11947 67547 12003 67603
rect 12089 67547 12145 67603
rect 12231 67547 12287 67603
rect 12373 67547 12429 67603
rect 12515 67547 12571 67603
rect 12657 67547 12713 67603
rect 12799 67547 12855 67603
rect 12941 67547 12997 67603
rect 13083 67547 13139 67603
rect 13225 67547 13281 67603
rect 13367 67547 13423 67603
rect 13509 67547 13565 67603
rect 13651 67547 13707 67603
rect 13793 67547 13849 67603
rect 13935 67547 13991 67603
rect 14077 67547 14133 67603
rect 14219 67547 14275 67603
rect 14361 67547 14417 67603
rect 14503 67547 14559 67603
rect 14645 67547 14701 67603
rect 14787 67547 14843 67603
rect 161 67405 217 67461
rect 303 67405 359 67461
rect 445 67405 501 67461
rect 587 67405 643 67461
rect 729 67405 785 67461
rect 871 67405 927 67461
rect 1013 67405 1069 67461
rect 1155 67405 1211 67461
rect 1297 67405 1353 67461
rect 1439 67405 1495 67461
rect 1581 67405 1637 67461
rect 1723 67405 1779 67461
rect 1865 67405 1921 67461
rect 2007 67405 2063 67461
rect 2149 67405 2205 67461
rect 2291 67405 2347 67461
rect 2433 67405 2489 67461
rect 2575 67405 2631 67461
rect 2717 67405 2773 67461
rect 2859 67405 2915 67461
rect 3001 67405 3057 67461
rect 3143 67405 3199 67461
rect 3285 67405 3341 67461
rect 3427 67405 3483 67461
rect 3569 67405 3625 67461
rect 3711 67405 3767 67461
rect 3853 67405 3909 67461
rect 3995 67405 4051 67461
rect 4137 67405 4193 67461
rect 4279 67405 4335 67461
rect 4421 67405 4477 67461
rect 4563 67405 4619 67461
rect 4705 67405 4761 67461
rect 4847 67405 4903 67461
rect 4989 67405 5045 67461
rect 5131 67405 5187 67461
rect 5273 67405 5329 67461
rect 5415 67405 5471 67461
rect 5557 67405 5613 67461
rect 5699 67405 5755 67461
rect 5841 67405 5897 67461
rect 5983 67405 6039 67461
rect 6125 67405 6181 67461
rect 6267 67405 6323 67461
rect 6409 67405 6465 67461
rect 6551 67405 6607 67461
rect 6693 67405 6749 67461
rect 6835 67405 6891 67461
rect 6977 67405 7033 67461
rect 7119 67405 7175 67461
rect 7261 67405 7317 67461
rect 7403 67405 7459 67461
rect 7545 67405 7601 67461
rect 7687 67405 7743 67461
rect 7829 67405 7885 67461
rect 7971 67405 8027 67461
rect 8113 67405 8169 67461
rect 8255 67405 8311 67461
rect 8397 67405 8453 67461
rect 8539 67405 8595 67461
rect 8681 67405 8737 67461
rect 8823 67405 8879 67461
rect 8965 67405 9021 67461
rect 9107 67405 9163 67461
rect 9249 67405 9305 67461
rect 9391 67405 9447 67461
rect 9533 67405 9589 67461
rect 9675 67405 9731 67461
rect 9817 67405 9873 67461
rect 9959 67405 10015 67461
rect 10101 67405 10157 67461
rect 10243 67405 10299 67461
rect 10385 67405 10441 67461
rect 10527 67405 10583 67461
rect 10669 67405 10725 67461
rect 10811 67405 10867 67461
rect 10953 67405 11009 67461
rect 11095 67405 11151 67461
rect 11237 67405 11293 67461
rect 11379 67405 11435 67461
rect 11521 67405 11577 67461
rect 11663 67405 11719 67461
rect 11805 67405 11861 67461
rect 11947 67405 12003 67461
rect 12089 67405 12145 67461
rect 12231 67405 12287 67461
rect 12373 67405 12429 67461
rect 12515 67405 12571 67461
rect 12657 67405 12713 67461
rect 12799 67405 12855 67461
rect 12941 67405 12997 67461
rect 13083 67405 13139 67461
rect 13225 67405 13281 67461
rect 13367 67405 13423 67461
rect 13509 67405 13565 67461
rect 13651 67405 13707 67461
rect 13793 67405 13849 67461
rect 13935 67405 13991 67461
rect 14077 67405 14133 67461
rect 14219 67405 14275 67461
rect 14361 67405 14417 67461
rect 14503 67405 14559 67461
rect 14645 67405 14701 67461
rect 14787 67405 14843 67461
rect 161 67263 217 67319
rect 303 67263 359 67319
rect 445 67263 501 67319
rect 587 67263 643 67319
rect 729 67263 785 67319
rect 871 67263 927 67319
rect 1013 67263 1069 67319
rect 1155 67263 1211 67319
rect 1297 67263 1353 67319
rect 1439 67263 1495 67319
rect 1581 67263 1637 67319
rect 1723 67263 1779 67319
rect 1865 67263 1921 67319
rect 2007 67263 2063 67319
rect 2149 67263 2205 67319
rect 2291 67263 2347 67319
rect 2433 67263 2489 67319
rect 2575 67263 2631 67319
rect 2717 67263 2773 67319
rect 2859 67263 2915 67319
rect 3001 67263 3057 67319
rect 3143 67263 3199 67319
rect 3285 67263 3341 67319
rect 3427 67263 3483 67319
rect 3569 67263 3625 67319
rect 3711 67263 3767 67319
rect 3853 67263 3909 67319
rect 3995 67263 4051 67319
rect 4137 67263 4193 67319
rect 4279 67263 4335 67319
rect 4421 67263 4477 67319
rect 4563 67263 4619 67319
rect 4705 67263 4761 67319
rect 4847 67263 4903 67319
rect 4989 67263 5045 67319
rect 5131 67263 5187 67319
rect 5273 67263 5329 67319
rect 5415 67263 5471 67319
rect 5557 67263 5613 67319
rect 5699 67263 5755 67319
rect 5841 67263 5897 67319
rect 5983 67263 6039 67319
rect 6125 67263 6181 67319
rect 6267 67263 6323 67319
rect 6409 67263 6465 67319
rect 6551 67263 6607 67319
rect 6693 67263 6749 67319
rect 6835 67263 6891 67319
rect 6977 67263 7033 67319
rect 7119 67263 7175 67319
rect 7261 67263 7317 67319
rect 7403 67263 7459 67319
rect 7545 67263 7601 67319
rect 7687 67263 7743 67319
rect 7829 67263 7885 67319
rect 7971 67263 8027 67319
rect 8113 67263 8169 67319
rect 8255 67263 8311 67319
rect 8397 67263 8453 67319
rect 8539 67263 8595 67319
rect 8681 67263 8737 67319
rect 8823 67263 8879 67319
rect 8965 67263 9021 67319
rect 9107 67263 9163 67319
rect 9249 67263 9305 67319
rect 9391 67263 9447 67319
rect 9533 67263 9589 67319
rect 9675 67263 9731 67319
rect 9817 67263 9873 67319
rect 9959 67263 10015 67319
rect 10101 67263 10157 67319
rect 10243 67263 10299 67319
rect 10385 67263 10441 67319
rect 10527 67263 10583 67319
rect 10669 67263 10725 67319
rect 10811 67263 10867 67319
rect 10953 67263 11009 67319
rect 11095 67263 11151 67319
rect 11237 67263 11293 67319
rect 11379 67263 11435 67319
rect 11521 67263 11577 67319
rect 11663 67263 11719 67319
rect 11805 67263 11861 67319
rect 11947 67263 12003 67319
rect 12089 67263 12145 67319
rect 12231 67263 12287 67319
rect 12373 67263 12429 67319
rect 12515 67263 12571 67319
rect 12657 67263 12713 67319
rect 12799 67263 12855 67319
rect 12941 67263 12997 67319
rect 13083 67263 13139 67319
rect 13225 67263 13281 67319
rect 13367 67263 13423 67319
rect 13509 67263 13565 67319
rect 13651 67263 13707 67319
rect 13793 67263 13849 67319
rect 13935 67263 13991 67319
rect 14077 67263 14133 67319
rect 14219 67263 14275 67319
rect 14361 67263 14417 67319
rect 14503 67263 14559 67319
rect 14645 67263 14701 67319
rect 14787 67263 14843 67319
rect 161 67121 217 67177
rect 303 67121 359 67177
rect 445 67121 501 67177
rect 587 67121 643 67177
rect 729 67121 785 67177
rect 871 67121 927 67177
rect 1013 67121 1069 67177
rect 1155 67121 1211 67177
rect 1297 67121 1353 67177
rect 1439 67121 1495 67177
rect 1581 67121 1637 67177
rect 1723 67121 1779 67177
rect 1865 67121 1921 67177
rect 2007 67121 2063 67177
rect 2149 67121 2205 67177
rect 2291 67121 2347 67177
rect 2433 67121 2489 67177
rect 2575 67121 2631 67177
rect 2717 67121 2773 67177
rect 2859 67121 2915 67177
rect 3001 67121 3057 67177
rect 3143 67121 3199 67177
rect 3285 67121 3341 67177
rect 3427 67121 3483 67177
rect 3569 67121 3625 67177
rect 3711 67121 3767 67177
rect 3853 67121 3909 67177
rect 3995 67121 4051 67177
rect 4137 67121 4193 67177
rect 4279 67121 4335 67177
rect 4421 67121 4477 67177
rect 4563 67121 4619 67177
rect 4705 67121 4761 67177
rect 4847 67121 4903 67177
rect 4989 67121 5045 67177
rect 5131 67121 5187 67177
rect 5273 67121 5329 67177
rect 5415 67121 5471 67177
rect 5557 67121 5613 67177
rect 5699 67121 5755 67177
rect 5841 67121 5897 67177
rect 5983 67121 6039 67177
rect 6125 67121 6181 67177
rect 6267 67121 6323 67177
rect 6409 67121 6465 67177
rect 6551 67121 6607 67177
rect 6693 67121 6749 67177
rect 6835 67121 6891 67177
rect 6977 67121 7033 67177
rect 7119 67121 7175 67177
rect 7261 67121 7317 67177
rect 7403 67121 7459 67177
rect 7545 67121 7601 67177
rect 7687 67121 7743 67177
rect 7829 67121 7885 67177
rect 7971 67121 8027 67177
rect 8113 67121 8169 67177
rect 8255 67121 8311 67177
rect 8397 67121 8453 67177
rect 8539 67121 8595 67177
rect 8681 67121 8737 67177
rect 8823 67121 8879 67177
rect 8965 67121 9021 67177
rect 9107 67121 9163 67177
rect 9249 67121 9305 67177
rect 9391 67121 9447 67177
rect 9533 67121 9589 67177
rect 9675 67121 9731 67177
rect 9817 67121 9873 67177
rect 9959 67121 10015 67177
rect 10101 67121 10157 67177
rect 10243 67121 10299 67177
rect 10385 67121 10441 67177
rect 10527 67121 10583 67177
rect 10669 67121 10725 67177
rect 10811 67121 10867 67177
rect 10953 67121 11009 67177
rect 11095 67121 11151 67177
rect 11237 67121 11293 67177
rect 11379 67121 11435 67177
rect 11521 67121 11577 67177
rect 11663 67121 11719 67177
rect 11805 67121 11861 67177
rect 11947 67121 12003 67177
rect 12089 67121 12145 67177
rect 12231 67121 12287 67177
rect 12373 67121 12429 67177
rect 12515 67121 12571 67177
rect 12657 67121 12713 67177
rect 12799 67121 12855 67177
rect 12941 67121 12997 67177
rect 13083 67121 13139 67177
rect 13225 67121 13281 67177
rect 13367 67121 13423 67177
rect 13509 67121 13565 67177
rect 13651 67121 13707 67177
rect 13793 67121 13849 67177
rect 13935 67121 13991 67177
rect 14077 67121 14133 67177
rect 14219 67121 14275 67177
rect 14361 67121 14417 67177
rect 14503 67121 14559 67177
rect 14645 67121 14701 67177
rect 14787 67121 14843 67177
rect 161 66979 217 67035
rect 303 66979 359 67035
rect 445 66979 501 67035
rect 587 66979 643 67035
rect 729 66979 785 67035
rect 871 66979 927 67035
rect 1013 66979 1069 67035
rect 1155 66979 1211 67035
rect 1297 66979 1353 67035
rect 1439 66979 1495 67035
rect 1581 66979 1637 67035
rect 1723 66979 1779 67035
rect 1865 66979 1921 67035
rect 2007 66979 2063 67035
rect 2149 66979 2205 67035
rect 2291 66979 2347 67035
rect 2433 66979 2489 67035
rect 2575 66979 2631 67035
rect 2717 66979 2773 67035
rect 2859 66979 2915 67035
rect 3001 66979 3057 67035
rect 3143 66979 3199 67035
rect 3285 66979 3341 67035
rect 3427 66979 3483 67035
rect 3569 66979 3625 67035
rect 3711 66979 3767 67035
rect 3853 66979 3909 67035
rect 3995 66979 4051 67035
rect 4137 66979 4193 67035
rect 4279 66979 4335 67035
rect 4421 66979 4477 67035
rect 4563 66979 4619 67035
rect 4705 66979 4761 67035
rect 4847 66979 4903 67035
rect 4989 66979 5045 67035
rect 5131 66979 5187 67035
rect 5273 66979 5329 67035
rect 5415 66979 5471 67035
rect 5557 66979 5613 67035
rect 5699 66979 5755 67035
rect 5841 66979 5897 67035
rect 5983 66979 6039 67035
rect 6125 66979 6181 67035
rect 6267 66979 6323 67035
rect 6409 66979 6465 67035
rect 6551 66979 6607 67035
rect 6693 66979 6749 67035
rect 6835 66979 6891 67035
rect 6977 66979 7033 67035
rect 7119 66979 7175 67035
rect 7261 66979 7317 67035
rect 7403 66979 7459 67035
rect 7545 66979 7601 67035
rect 7687 66979 7743 67035
rect 7829 66979 7885 67035
rect 7971 66979 8027 67035
rect 8113 66979 8169 67035
rect 8255 66979 8311 67035
rect 8397 66979 8453 67035
rect 8539 66979 8595 67035
rect 8681 66979 8737 67035
rect 8823 66979 8879 67035
rect 8965 66979 9021 67035
rect 9107 66979 9163 67035
rect 9249 66979 9305 67035
rect 9391 66979 9447 67035
rect 9533 66979 9589 67035
rect 9675 66979 9731 67035
rect 9817 66979 9873 67035
rect 9959 66979 10015 67035
rect 10101 66979 10157 67035
rect 10243 66979 10299 67035
rect 10385 66979 10441 67035
rect 10527 66979 10583 67035
rect 10669 66979 10725 67035
rect 10811 66979 10867 67035
rect 10953 66979 11009 67035
rect 11095 66979 11151 67035
rect 11237 66979 11293 67035
rect 11379 66979 11435 67035
rect 11521 66979 11577 67035
rect 11663 66979 11719 67035
rect 11805 66979 11861 67035
rect 11947 66979 12003 67035
rect 12089 66979 12145 67035
rect 12231 66979 12287 67035
rect 12373 66979 12429 67035
rect 12515 66979 12571 67035
rect 12657 66979 12713 67035
rect 12799 66979 12855 67035
rect 12941 66979 12997 67035
rect 13083 66979 13139 67035
rect 13225 66979 13281 67035
rect 13367 66979 13423 67035
rect 13509 66979 13565 67035
rect 13651 66979 13707 67035
rect 13793 66979 13849 67035
rect 13935 66979 13991 67035
rect 14077 66979 14133 67035
rect 14219 66979 14275 67035
rect 14361 66979 14417 67035
rect 14503 66979 14559 67035
rect 14645 66979 14701 67035
rect 14787 66979 14843 67035
rect 161 66837 217 66893
rect 303 66837 359 66893
rect 445 66837 501 66893
rect 587 66837 643 66893
rect 729 66837 785 66893
rect 871 66837 927 66893
rect 1013 66837 1069 66893
rect 1155 66837 1211 66893
rect 1297 66837 1353 66893
rect 1439 66837 1495 66893
rect 1581 66837 1637 66893
rect 1723 66837 1779 66893
rect 1865 66837 1921 66893
rect 2007 66837 2063 66893
rect 2149 66837 2205 66893
rect 2291 66837 2347 66893
rect 2433 66837 2489 66893
rect 2575 66837 2631 66893
rect 2717 66837 2773 66893
rect 2859 66837 2915 66893
rect 3001 66837 3057 66893
rect 3143 66837 3199 66893
rect 3285 66837 3341 66893
rect 3427 66837 3483 66893
rect 3569 66837 3625 66893
rect 3711 66837 3767 66893
rect 3853 66837 3909 66893
rect 3995 66837 4051 66893
rect 4137 66837 4193 66893
rect 4279 66837 4335 66893
rect 4421 66837 4477 66893
rect 4563 66837 4619 66893
rect 4705 66837 4761 66893
rect 4847 66837 4903 66893
rect 4989 66837 5045 66893
rect 5131 66837 5187 66893
rect 5273 66837 5329 66893
rect 5415 66837 5471 66893
rect 5557 66837 5613 66893
rect 5699 66837 5755 66893
rect 5841 66837 5897 66893
rect 5983 66837 6039 66893
rect 6125 66837 6181 66893
rect 6267 66837 6323 66893
rect 6409 66837 6465 66893
rect 6551 66837 6607 66893
rect 6693 66837 6749 66893
rect 6835 66837 6891 66893
rect 6977 66837 7033 66893
rect 7119 66837 7175 66893
rect 7261 66837 7317 66893
rect 7403 66837 7459 66893
rect 7545 66837 7601 66893
rect 7687 66837 7743 66893
rect 7829 66837 7885 66893
rect 7971 66837 8027 66893
rect 8113 66837 8169 66893
rect 8255 66837 8311 66893
rect 8397 66837 8453 66893
rect 8539 66837 8595 66893
rect 8681 66837 8737 66893
rect 8823 66837 8879 66893
rect 8965 66837 9021 66893
rect 9107 66837 9163 66893
rect 9249 66837 9305 66893
rect 9391 66837 9447 66893
rect 9533 66837 9589 66893
rect 9675 66837 9731 66893
rect 9817 66837 9873 66893
rect 9959 66837 10015 66893
rect 10101 66837 10157 66893
rect 10243 66837 10299 66893
rect 10385 66837 10441 66893
rect 10527 66837 10583 66893
rect 10669 66837 10725 66893
rect 10811 66837 10867 66893
rect 10953 66837 11009 66893
rect 11095 66837 11151 66893
rect 11237 66837 11293 66893
rect 11379 66837 11435 66893
rect 11521 66837 11577 66893
rect 11663 66837 11719 66893
rect 11805 66837 11861 66893
rect 11947 66837 12003 66893
rect 12089 66837 12145 66893
rect 12231 66837 12287 66893
rect 12373 66837 12429 66893
rect 12515 66837 12571 66893
rect 12657 66837 12713 66893
rect 12799 66837 12855 66893
rect 12941 66837 12997 66893
rect 13083 66837 13139 66893
rect 13225 66837 13281 66893
rect 13367 66837 13423 66893
rect 13509 66837 13565 66893
rect 13651 66837 13707 66893
rect 13793 66837 13849 66893
rect 13935 66837 13991 66893
rect 14077 66837 14133 66893
rect 14219 66837 14275 66893
rect 14361 66837 14417 66893
rect 14503 66837 14559 66893
rect 14645 66837 14701 66893
rect 14787 66837 14843 66893
rect 161 66515 217 66571
rect 303 66515 359 66571
rect 445 66515 501 66571
rect 587 66515 643 66571
rect 729 66515 785 66571
rect 871 66515 927 66571
rect 1013 66515 1069 66571
rect 1155 66515 1211 66571
rect 1297 66515 1353 66571
rect 1439 66515 1495 66571
rect 1581 66515 1637 66571
rect 1723 66515 1779 66571
rect 1865 66515 1921 66571
rect 2007 66515 2063 66571
rect 2149 66515 2205 66571
rect 2291 66515 2347 66571
rect 2433 66515 2489 66571
rect 2575 66515 2631 66571
rect 2717 66515 2773 66571
rect 2859 66515 2915 66571
rect 3001 66515 3057 66571
rect 3143 66515 3199 66571
rect 3285 66515 3341 66571
rect 3427 66515 3483 66571
rect 3569 66515 3625 66571
rect 3711 66515 3767 66571
rect 3853 66515 3909 66571
rect 3995 66515 4051 66571
rect 4137 66515 4193 66571
rect 4279 66515 4335 66571
rect 4421 66515 4477 66571
rect 4563 66515 4619 66571
rect 4705 66515 4761 66571
rect 4847 66515 4903 66571
rect 4989 66515 5045 66571
rect 5131 66515 5187 66571
rect 5273 66515 5329 66571
rect 5415 66515 5471 66571
rect 5557 66515 5613 66571
rect 5699 66515 5755 66571
rect 5841 66515 5897 66571
rect 5983 66515 6039 66571
rect 6125 66515 6181 66571
rect 6267 66515 6323 66571
rect 6409 66515 6465 66571
rect 6551 66515 6607 66571
rect 6693 66515 6749 66571
rect 6835 66515 6891 66571
rect 6977 66515 7033 66571
rect 7119 66515 7175 66571
rect 7261 66515 7317 66571
rect 7403 66515 7459 66571
rect 7545 66515 7601 66571
rect 7687 66515 7743 66571
rect 7829 66515 7885 66571
rect 7971 66515 8027 66571
rect 8113 66515 8169 66571
rect 8255 66515 8311 66571
rect 8397 66515 8453 66571
rect 8539 66515 8595 66571
rect 8681 66515 8737 66571
rect 8823 66515 8879 66571
rect 8965 66515 9021 66571
rect 9107 66515 9163 66571
rect 9249 66515 9305 66571
rect 9391 66515 9447 66571
rect 9533 66515 9589 66571
rect 9675 66515 9731 66571
rect 9817 66515 9873 66571
rect 9959 66515 10015 66571
rect 10101 66515 10157 66571
rect 10243 66515 10299 66571
rect 10385 66515 10441 66571
rect 10527 66515 10583 66571
rect 10669 66515 10725 66571
rect 10811 66515 10867 66571
rect 10953 66515 11009 66571
rect 11095 66515 11151 66571
rect 11237 66515 11293 66571
rect 11379 66515 11435 66571
rect 11521 66515 11577 66571
rect 11663 66515 11719 66571
rect 11805 66515 11861 66571
rect 11947 66515 12003 66571
rect 12089 66515 12145 66571
rect 12231 66515 12287 66571
rect 12373 66515 12429 66571
rect 12515 66515 12571 66571
rect 12657 66515 12713 66571
rect 12799 66515 12855 66571
rect 12941 66515 12997 66571
rect 13083 66515 13139 66571
rect 13225 66515 13281 66571
rect 13367 66515 13423 66571
rect 13509 66515 13565 66571
rect 13651 66515 13707 66571
rect 13793 66515 13849 66571
rect 13935 66515 13991 66571
rect 14077 66515 14133 66571
rect 14219 66515 14275 66571
rect 14361 66515 14417 66571
rect 14503 66515 14559 66571
rect 14645 66515 14701 66571
rect 14787 66515 14843 66571
rect 161 66373 217 66429
rect 303 66373 359 66429
rect 445 66373 501 66429
rect 587 66373 643 66429
rect 729 66373 785 66429
rect 871 66373 927 66429
rect 1013 66373 1069 66429
rect 1155 66373 1211 66429
rect 1297 66373 1353 66429
rect 1439 66373 1495 66429
rect 1581 66373 1637 66429
rect 1723 66373 1779 66429
rect 1865 66373 1921 66429
rect 2007 66373 2063 66429
rect 2149 66373 2205 66429
rect 2291 66373 2347 66429
rect 2433 66373 2489 66429
rect 2575 66373 2631 66429
rect 2717 66373 2773 66429
rect 2859 66373 2915 66429
rect 3001 66373 3057 66429
rect 3143 66373 3199 66429
rect 3285 66373 3341 66429
rect 3427 66373 3483 66429
rect 3569 66373 3625 66429
rect 3711 66373 3767 66429
rect 3853 66373 3909 66429
rect 3995 66373 4051 66429
rect 4137 66373 4193 66429
rect 4279 66373 4335 66429
rect 4421 66373 4477 66429
rect 4563 66373 4619 66429
rect 4705 66373 4761 66429
rect 4847 66373 4903 66429
rect 4989 66373 5045 66429
rect 5131 66373 5187 66429
rect 5273 66373 5329 66429
rect 5415 66373 5471 66429
rect 5557 66373 5613 66429
rect 5699 66373 5755 66429
rect 5841 66373 5897 66429
rect 5983 66373 6039 66429
rect 6125 66373 6181 66429
rect 6267 66373 6323 66429
rect 6409 66373 6465 66429
rect 6551 66373 6607 66429
rect 6693 66373 6749 66429
rect 6835 66373 6891 66429
rect 6977 66373 7033 66429
rect 7119 66373 7175 66429
rect 7261 66373 7317 66429
rect 7403 66373 7459 66429
rect 7545 66373 7601 66429
rect 7687 66373 7743 66429
rect 7829 66373 7885 66429
rect 7971 66373 8027 66429
rect 8113 66373 8169 66429
rect 8255 66373 8311 66429
rect 8397 66373 8453 66429
rect 8539 66373 8595 66429
rect 8681 66373 8737 66429
rect 8823 66373 8879 66429
rect 8965 66373 9021 66429
rect 9107 66373 9163 66429
rect 9249 66373 9305 66429
rect 9391 66373 9447 66429
rect 9533 66373 9589 66429
rect 9675 66373 9731 66429
rect 9817 66373 9873 66429
rect 9959 66373 10015 66429
rect 10101 66373 10157 66429
rect 10243 66373 10299 66429
rect 10385 66373 10441 66429
rect 10527 66373 10583 66429
rect 10669 66373 10725 66429
rect 10811 66373 10867 66429
rect 10953 66373 11009 66429
rect 11095 66373 11151 66429
rect 11237 66373 11293 66429
rect 11379 66373 11435 66429
rect 11521 66373 11577 66429
rect 11663 66373 11719 66429
rect 11805 66373 11861 66429
rect 11947 66373 12003 66429
rect 12089 66373 12145 66429
rect 12231 66373 12287 66429
rect 12373 66373 12429 66429
rect 12515 66373 12571 66429
rect 12657 66373 12713 66429
rect 12799 66373 12855 66429
rect 12941 66373 12997 66429
rect 13083 66373 13139 66429
rect 13225 66373 13281 66429
rect 13367 66373 13423 66429
rect 13509 66373 13565 66429
rect 13651 66373 13707 66429
rect 13793 66373 13849 66429
rect 13935 66373 13991 66429
rect 14077 66373 14133 66429
rect 14219 66373 14275 66429
rect 14361 66373 14417 66429
rect 14503 66373 14559 66429
rect 14645 66373 14701 66429
rect 14787 66373 14843 66429
rect 161 66231 217 66287
rect 303 66231 359 66287
rect 445 66231 501 66287
rect 587 66231 643 66287
rect 729 66231 785 66287
rect 871 66231 927 66287
rect 1013 66231 1069 66287
rect 1155 66231 1211 66287
rect 1297 66231 1353 66287
rect 1439 66231 1495 66287
rect 1581 66231 1637 66287
rect 1723 66231 1779 66287
rect 1865 66231 1921 66287
rect 2007 66231 2063 66287
rect 2149 66231 2205 66287
rect 2291 66231 2347 66287
rect 2433 66231 2489 66287
rect 2575 66231 2631 66287
rect 2717 66231 2773 66287
rect 2859 66231 2915 66287
rect 3001 66231 3057 66287
rect 3143 66231 3199 66287
rect 3285 66231 3341 66287
rect 3427 66231 3483 66287
rect 3569 66231 3625 66287
rect 3711 66231 3767 66287
rect 3853 66231 3909 66287
rect 3995 66231 4051 66287
rect 4137 66231 4193 66287
rect 4279 66231 4335 66287
rect 4421 66231 4477 66287
rect 4563 66231 4619 66287
rect 4705 66231 4761 66287
rect 4847 66231 4903 66287
rect 4989 66231 5045 66287
rect 5131 66231 5187 66287
rect 5273 66231 5329 66287
rect 5415 66231 5471 66287
rect 5557 66231 5613 66287
rect 5699 66231 5755 66287
rect 5841 66231 5897 66287
rect 5983 66231 6039 66287
rect 6125 66231 6181 66287
rect 6267 66231 6323 66287
rect 6409 66231 6465 66287
rect 6551 66231 6607 66287
rect 6693 66231 6749 66287
rect 6835 66231 6891 66287
rect 6977 66231 7033 66287
rect 7119 66231 7175 66287
rect 7261 66231 7317 66287
rect 7403 66231 7459 66287
rect 7545 66231 7601 66287
rect 7687 66231 7743 66287
rect 7829 66231 7885 66287
rect 7971 66231 8027 66287
rect 8113 66231 8169 66287
rect 8255 66231 8311 66287
rect 8397 66231 8453 66287
rect 8539 66231 8595 66287
rect 8681 66231 8737 66287
rect 8823 66231 8879 66287
rect 8965 66231 9021 66287
rect 9107 66231 9163 66287
rect 9249 66231 9305 66287
rect 9391 66231 9447 66287
rect 9533 66231 9589 66287
rect 9675 66231 9731 66287
rect 9817 66231 9873 66287
rect 9959 66231 10015 66287
rect 10101 66231 10157 66287
rect 10243 66231 10299 66287
rect 10385 66231 10441 66287
rect 10527 66231 10583 66287
rect 10669 66231 10725 66287
rect 10811 66231 10867 66287
rect 10953 66231 11009 66287
rect 11095 66231 11151 66287
rect 11237 66231 11293 66287
rect 11379 66231 11435 66287
rect 11521 66231 11577 66287
rect 11663 66231 11719 66287
rect 11805 66231 11861 66287
rect 11947 66231 12003 66287
rect 12089 66231 12145 66287
rect 12231 66231 12287 66287
rect 12373 66231 12429 66287
rect 12515 66231 12571 66287
rect 12657 66231 12713 66287
rect 12799 66231 12855 66287
rect 12941 66231 12997 66287
rect 13083 66231 13139 66287
rect 13225 66231 13281 66287
rect 13367 66231 13423 66287
rect 13509 66231 13565 66287
rect 13651 66231 13707 66287
rect 13793 66231 13849 66287
rect 13935 66231 13991 66287
rect 14077 66231 14133 66287
rect 14219 66231 14275 66287
rect 14361 66231 14417 66287
rect 14503 66231 14559 66287
rect 14645 66231 14701 66287
rect 14787 66231 14843 66287
rect 161 66089 217 66145
rect 303 66089 359 66145
rect 445 66089 501 66145
rect 587 66089 643 66145
rect 729 66089 785 66145
rect 871 66089 927 66145
rect 1013 66089 1069 66145
rect 1155 66089 1211 66145
rect 1297 66089 1353 66145
rect 1439 66089 1495 66145
rect 1581 66089 1637 66145
rect 1723 66089 1779 66145
rect 1865 66089 1921 66145
rect 2007 66089 2063 66145
rect 2149 66089 2205 66145
rect 2291 66089 2347 66145
rect 2433 66089 2489 66145
rect 2575 66089 2631 66145
rect 2717 66089 2773 66145
rect 2859 66089 2915 66145
rect 3001 66089 3057 66145
rect 3143 66089 3199 66145
rect 3285 66089 3341 66145
rect 3427 66089 3483 66145
rect 3569 66089 3625 66145
rect 3711 66089 3767 66145
rect 3853 66089 3909 66145
rect 3995 66089 4051 66145
rect 4137 66089 4193 66145
rect 4279 66089 4335 66145
rect 4421 66089 4477 66145
rect 4563 66089 4619 66145
rect 4705 66089 4761 66145
rect 4847 66089 4903 66145
rect 4989 66089 5045 66145
rect 5131 66089 5187 66145
rect 5273 66089 5329 66145
rect 5415 66089 5471 66145
rect 5557 66089 5613 66145
rect 5699 66089 5755 66145
rect 5841 66089 5897 66145
rect 5983 66089 6039 66145
rect 6125 66089 6181 66145
rect 6267 66089 6323 66145
rect 6409 66089 6465 66145
rect 6551 66089 6607 66145
rect 6693 66089 6749 66145
rect 6835 66089 6891 66145
rect 6977 66089 7033 66145
rect 7119 66089 7175 66145
rect 7261 66089 7317 66145
rect 7403 66089 7459 66145
rect 7545 66089 7601 66145
rect 7687 66089 7743 66145
rect 7829 66089 7885 66145
rect 7971 66089 8027 66145
rect 8113 66089 8169 66145
rect 8255 66089 8311 66145
rect 8397 66089 8453 66145
rect 8539 66089 8595 66145
rect 8681 66089 8737 66145
rect 8823 66089 8879 66145
rect 8965 66089 9021 66145
rect 9107 66089 9163 66145
rect 9249 66089 9305 66145
rect 9391 66089 9447 66145
rect 9533 66089 9589 66145
rect 9675 66089 9731 66145
rect 9817 66089 9873 66145
rect 9959 66089 10015 66145
rect 10101 66089 10157 66145
rect 10243 66089 10299 66145
rect 10385 66089 10441 66145
rect 10527 66089 10583 66145
rect 10669 66089 10725 66145
rect 10811 66089 10867 66145
rect 10953 66089 11009 66145
rect 11095 66089 11151 66145
rect 11237 66089 11293 66145
rect 11379 66089 11435 66145
rect 11521 66089 11577 66145
rect 11663 66089 11719 66145
rect 11805 66089 11861 66145
rect 11947 66089 12003 66145
rect 12089 66089 12145 66145
rect 12231 66089 12287 66145
rect 12373 66089 12429 66145
rect 12515 66089 12571 66145
rect 12657 66089 12713 66145
rect 12799 66089 12855 66145
rect 12941 66089 12997 66145
rect 13083 66089 13139 66145
rect 13225 66089 13281 66145
rect 13367 66089 13423 66145
rect 13509 66089 13565 66145
rect 13651 66089 13707 66145
rect 13793 66089 13849 66145
rect 13935 66089 13991 66145
rect 14077 66089 14133 66145
rect 14219 66089 14275 66145
rect 14361 66089 14417 66145
rect 14503 66089 14559 66145
rect 14645 66089 14701 66145
rect 14787 66089 14843 66145
rect 161 65947 217 66003
rect 303 65947 359 66003
rect 445 65947 501 66003
rect 587 65947 643 66003
rect 729 65947 785 66003
rect 871 65947 927 66003
rect 1013 65947 1069 66003
rect 1155 65947 1211 66003
rect 1297 65947 1353 66003
rect 1439 65947 1495 66003
rect 1581 65947 1637 66003
rect 1723 65947 1779 66003
rect 1865 65947 1921 66003
rect 2007 65947 2063 66003
rect 2149 65947 2205 66003
rect 2291 65947 2347 66003
rect 2433 65947 2489 66003
rect 2575 65947 2631 66003
rect 2717 65947 2773 66003
rect 2859 65947 2915 66003
rect 3001 65947 3057 66003
rect 3143 65947 3199 66003
rect 3285 65947 3341 66003
rect 3427 65947 3483 66003
rect 3569 65947 3625 66003
rect 3711 65947 3767 66003
rect 3853 65947 3909 66003
rect 3995 65947 4051 66003
rect 4137 65947 4193 66003
rect 4279 65947 4335 66003
rect 4421 65947 4477 66003
rect 4563 65947 4619 66003
rect 4705 65947 4761 66003
rect 4847 65947 4903 66003
rect 4989 65947 5045 66003
rect 5131 65947 5187 66003
rect 5273 65947 5329 66003
rect 5415 65947 5471 66003
rect 5557 65947 5613 66003
rect 5699 65947 5755 66003
rect 5841 65947 5897 66003
rect 5983 65947 6039 66003
rect 6125 65947 6181 66003
rect 6267 65947 6323 66003
rect 6409 65947 6465 66003
rect 6551 65947 6607 66003
rect 6693 65947 6749 66003
rect 6835 65947 6891 66003
rect 6977 65947 7033 66003
rect 7119 65947 7175 66003
rect 7261 65947 7317 66003
rect 7403 65947 7459 66003
rect 7545 65947 7601 66003
rect 7687 65947 7743 66003
rect 7829 65947 7885 66003
rect 7971 65947 8027 66003
rect 8113 65947 8169 66003
rect 8255 65947 8311 66003
rect 8397 65947 8453 66003
rect 8539 65947 8595 66003
rect 8681 65947 8737 66003
rect 8823 65947 8879 66003
rect 8965 65947 9021 66003
rect 9107 65947 9163 66003
rect 9249 65947 9305 66003
rect 9391 65947 9447 66003
rect 9533 65947 9589 66003
rect 9675 65947 9731 66003
rect 9817 65947 9873 66003
rect 9959 65947 10015 66003
rect 10101 65947 10157 66003
rect 10243 65947 10299 66003
rect 10385 65947 10441 66003
rect 10527 65947 10583 66003
rect 10669 65947 10725 66003
rect 10811 65947 10867 66003
rect 10953 65947 11009 66003
rect 11095 65947 11151 66003
rect 11237 65947 11293 66003
rect 11379 65947 11435 66003
rect 11521 65947 11577 66003
rect 11663 65947 11719 66003
rect 11805 65947 11861 66003
rect 11947 65947 12003 66003
rect 12089 65947 12145 66003
rect 12231 65947 12287 66003
rect 12373 65947 12429 66003
rect 12515 65947 12571 66003
rect 12657 65947 12713 66003
rect 12799 65947 12855 66003
rect 12941 65947 12997 66003
rect 13083 65947 13139 66003
rect 13225 65947 13281 66003
rect 13367 65947 13423 66003
rect 13509 65947 13565 66003
rect 13651 65947 13707 66003
rect 13793 65947 13849 66003
rect 13935 65947 13991 66003
rect 14077 65947 14133 66003
rect 14219 65947 14275 66003
rect 14361 65947 14417 66003
rect 14503 65947 14559 66003
rect 14645 65947 14701 66003
rect 14787 65947 14843 66003
rect 161 65805 217 65861
rect 303 65805 359 65861
rect 445 65805 501 65861
rect 587 65805 643 65861
rect 729 65805 785 65861
rect 871 65805 927 65861
rect 1013 65805 1069 65861
rect 1155 65805 1211 65861
rect 1297 65805 1353 65861
rect 1439 65805 1495 65861
rect 1581 65805 1637 65861
rect 1723 65805 1779 65861
rect 1865 65805 1921 65861
rect 2007 65805 2063 65861
rect 2149 65805 2205 65861
rect 2291 65805 2347 65861
rect 2433 65805 2489 65861
rect 2575 65805 2631 65861
rect 2717 65805 2773 65861
rect 2859 65805 2915 65861
rect 3001 65805 3057 65861
rect 3143 65805 3199 65861
rect 3285 65805 3341 65861
rect 3427 65805 3483 65861
rect 3569 65805 3625 65861
rect 3711 65805 3767 65861
rect 3853 65805 3909 65861
rect 3995 65805 4051 65861
rect 4137 65805 4193 65861
rect 4279 65805 4335 65861
rect 4421 65805 4477 65861
rect 4563 65805 4619 65861
rect 4705 65805 4761 65861
rect 4847 65805 4903 65861
rect 4989 65805 5045 65861
rect 5131 65805 5187 65861
rect 5273 65805 5329 65861
rect 5415 65805 5471 65861
rect 5557 65805 5613 65861
rect 5699 65805 5755 65861
rect 5841 65805 5897 65861
rect 5983 65805 6039 65861
rect 6125 65805 6181 65861
rect 6267 65805 6323 65861
rect 6409 65805 6465 65861
rect 6551 65805 6607 65861
rect 6693 65805 6749 65861
rect 6835 65805 6891 65861
rect 6977 65805 7033 65861
rect 7119 65805 7175 65861
rect 7261 65805 7317 65861
rect 7403 65805 7459 65861
rect 7545 65805 7601 65861
rect 7687 65805 7743 65861
rect 7829 65805 7885 65861
rect 7971 65805 8027 65861
rect 8113 65805 8169 65861
rect 8255 65805 8311 65861
rect 8397 65805 8453 65861
rect 8539 65805 8595 65861
rect 8681 65805 8737 65861
rect 8823 65805 8879 65861
rect 8965 65805 9021 65861
rect 9107 65805 9163 65861
rect 9249 65805 9305 65861
rect 9391 65805 9447 65861
rect 9533 65805 9589 65861
rect 9675 65805 9731 65861
rect 9817 65805 9873 65861
rect 9959 65805 10015 65861
rect 10101 65805 10157 65861
rect 10243 65805 10299 65861
rect 10385 65805 10441 65861
rect 10527 65805 10583 65861
rect 10669 65805 10725 65861
rect 10811 65805 10867 65861
rect 10953 65805 11009 65861
rect 11095 65805 11151 65861
rect 11237 65805 11293 65861
rect 11379 65805 11435 65861
rect 11521 65805 11577 65861
rect 11663 65805 11719 65861
rect 11805 65805 11861 65861
rect 11947 65805 12003 65861
rect 12089 65805 12145 65861
rect 12231 65805 12287 65861
rect 12373 65805 12429 65861
rect 12515 65805 12571 65861
rect 12657 65805 12713 65861
rect 12799 65805 12855 65861
rect 12941 65805 12997 65861
rect 13083 65805 13139 65861
rect 13225 65805 13281 65861
rect 13367 65805 13423 65861
rect 13509 65805 13565 65861
rect 13651 65805 13707 65861
rect 13793 65805 13849 65861
rect 13935 65805 13991 65861
rect 14077 65805 14133 65861
rect 14219 65805 14275 65861
rect 14361 65805 14417 65861
rect 14503 65805 14559 65861
rect 14645 65805 14701 65861
rect 14787 65805 14843 65861
rect 161 65663 217 65719
rect 303 65663 359 65719
rect 445 65663 501 65719
rect 587 65663 643 65719
rect 729 65663 785 65719
rect 871 65663 927 65719
rect 1013 65663 1069 65719
rect 1155 65663 1211 65719
rect 1297 65663 1353 65719
rect 1439 65663 1495 65719
rect 1581 65663 1637 65719
rect 1723 65663 1779 65719
rect 1865 65663 1921 65719
rect 2007 65663 2063 65719
rect 2149 65663 2205 65719
rect 2291 65663 2347 65719
rect 2433 65663 2489 65719
rect 2575 65663 2631 65719
rect 2717 65663 2773 65719
rect 2859 65663 2915 65719
rect 3001 65663 3057 65719
rect 3143 65663 3199 65719
rect 3285 65663 3341 65719
rect 3427 65663 3483 65719
rect 3569 65663 3625 65719
rect 3711 65663 3767 65719
rect 3853 65663 3909 65719
rect 3995 65663 4051 65719
rect 4137 65663 4193 65719
rect 4279 65663 4335 65719
rect 4421 65663 4477 65719
rect 4563 65663 4619 65719
rect 4705 65663 4761 65719
rect 4847 65663 4903 65719
rect 4989 65663 5045 65719
rect 5131 65663 5187 65719
rect 5273 65663 5329 65719
rect 5415 65663 5471 65719
rect 5557 65663 5613 65719
rect 5699 65663 5755 65719
rect 5841 65663 5897 65719
rect 5983 65663 6039 65719
rect 6125 65663 6181 65719
rect 6267 65663 6323 65719
rect 6409 65663 6465 65719
rect 6551 65663 6607 65719
rect 6693 65663 6749 65719
rect 6835 65663 6891 65719
rect 6977 65663 7033 65719
rect 7119 65663 7175 65719
rect 7261 65663 7317 65719
rect 7403 65663 7459 65719
rect 7545 65663 7601 65719
rect 7687 65663 7743 65719
rect 7829 65663 7885 65719
rect 7971 65663 8027 65719
rect 8113 65663 8169 65719
rect 8255 65663 8311 65719
rect 8397 65663 8453 65719
rect 8539 65663 8595 65719
rect 8681 65663 8737 65719
rect 8823 65663 8879 65719
rect 8965 65663 9021 65719
rect 9107 65663 9163 65719
rect 9249 65663 9305 65719
rect 9391 65663 9447 65719
rect 9533 65663 9589 65719
rect 9675 65663 9731 65719
rect 9817 65663 9873 65719
rect 9959 65663 10015 65719
rect 10101 65663 10157 65719
rect 10243 65663 10299 65719
rect 10385 65663 10441 65719
rect 10527 65663 10583 65719
rect 10669 65663 10725 65719
rect 10811 65663 10867 65719
rect 10953 65663 11009 65719
rect 11095 65663 11151 65719
rect 11237 65663 11293 65719
rect 11379 65663 11435 65719
rect 11521 65663 11577 65719
rect 11663 65663 11719 65719
rect 11805 65663 11861 65719
rect 11947 65663 12003 65719
rect 12089 65663 12145 65719
rect 12231 65663 12287 65719
rect 12373 65663 12429 65719
rect 12515 65663 12571 65719
rect 12657 65663 12713 65719
rect 12799 65663 12855 65719
rect 12941 65663 12997 65719
rect 13083 65663 13139 65719
rect 13225 65663 13281 65719
rect 13367 65663 13423 65719
rect 13509 65663 13565 65719
rect 13651 65663 13707 65719
rect 13793 65663 13849 65719
rect 13935 65663 13991 65719
rect 14077 65663 14133 65719
rect 14219 65663 14275 65719
rect 14361 65663 14417 65719
rect 14503 65663 14559 65719
rect 14645 65663 14701 65719
rect 14787 65663 14843 65719
rect 161 65521 217 65577
rect 303 65521 359 65577
rect 445 65521 501 65577
rect 587 65521 643 65577
rect 729 65521 785 65577
rect 871 65521 927 65577
rect 1013 65521 1069 65577
rect 1155 65521 1211 65577
rect 1297 65521 1353 65577
rect 1439 65521 1495 65577
rect 1581 65521 1637 65577
rect 1723 65521 1779 65577
rect 1865 65521 1921 65577
rect 2007 65521 2063 65577
rect 2149 65521 2205 65577
rect 2291 65521 2347 65577
rect 2433 65521 2489 65577
rect 2575 65521 2631 65577
rect 2717 65521 2773 65577
rect 2859 65521 2915 65577
rect 3001 65521 3057 65577
rect 3143 65521 3199 65577
rect 3285 65521 3341 65577
rect 3427 65521 3483 65577
rect 3569 65521 3625 65577
rect 3711 65521 3767 65577
rect 3853 65521 3909 65577
rect 3995 65521 4051 65577
rect 4137 65521 4193 65577
rect 4279 65521 4335 65577
rect 4421 65521 4477 65577
rect 4563 65521 4619 65577
rect 4705 65521 4761 65577
rect 4847 65521 4903 65577
rect 4989 65521 5045 65577
rect 5131 65521 5187 65577
rect 5273 65521 5329 65577
rect 5415 65521 5471 65577
rect 5557 65521 5613 65577
rect 5699 65521 5755 65577
rect 5841 65521 5897 65577
rect 5983 65521 6039 65577
rect 6125 65521 6181 65577
rect 6267 65521 6323 65577
rect 6409 65521 6465 65577
rect 6551 65521 6607 65577
rect 6693 65521 6749 65577
rect 6835 65521 6891 65577
rect 6977 65521 7033 65577
rect 7119 65521 7175 65577
rect 7261 65521 7317 65577
rect 7403 65521 7459 65577
rect 7545 65521 7601 65577
rect 7687 65521 7743 65577
rect 7829 65521 7885 65577
rect 7971 65521 8027 65577
rect 8113 65521 8169 65577
rect 8255 65521 8311 65577
rect 8397 65521 8453 65577
rect 8539 65521 8595 65577
rect 8681 65521 8737 65577
rect 8823 65521 8879 65577
rect 8965 65521 9021 65577
rect 9107 65521 9163 65577
rect 9249 65521 9305 65577
rect 9391 65521 9447 65577
rect 9533 65521 9589 65577
rect 9675 65521 9731 65577
rect 9817 65521 9873 65577
rect 9959 65521 10015 65577
rect 10101 65521 10157 65577
rect 10243 65521 10299 65577
rect 10385 65521 10441 65577
rect 10527 65521 10583 65577
rect 10669 65521 10725 65577
rect 10811 65521 10867 65577
rect 10953 65521 11009 65577
rect 11095 65521 11151 65577
rect 11237 65521 11293 65577
rect 11379 65521 11435 65577
rect 11521 65521 11577 65577
rect 11663 65521 11719 65577
rect 11805 65521 11861 65577
rect 11947 65521 12003 65577
rect 12089 65521 12145 65577
rect 12231 65521 12287 65577
rect 12373 65521 12429 65577
rect 12515 65521 12571 65577
rect 12657 65521 12713 65577
rect 12799 65521 12855 65577
rect 12941 65521 12997 65577
rect 13083 65521 13139 65577
rect 13225 65521 13281 65577
rect 13367 65521 13423 65577
rect 13509 65521 13565 65577
rect 13651 65521 13707 65577
rect 13793 65521 13849 65577
rect 13935 65521 13991 65577
rect 14077 65521 14133 65577
rect 14219 65521 14275 65577
rect 14361 65521 14417 65577
rect 14503 65521 14559 65577
rect 14645 65521 14701 65577
rect 14787 65521 14843 65577
rect 161 65379 217 65435
rect 303 65379 359 65435
rect 445 65379 501 65435
rect 587 65379 643 65435
rect 729 65379 785 65435
rect 871 65379 927 65435
rect 1013 65379 1069 65435
rect 1155 65379 1211 65435
rect 1297 65379 1353 65435
rect 1439 65379 1495 65435
rect 1581 65379 1637 65435
rect 1723 65379 1779 65435
rect 1865 65379 1921 65435
rect 2007 65379 2063 65435
rect 2149 65379 2205 65435
rect 2291 65379 2347 65435
rect 2433 65379 2489 65435
rect 2575 65379 2631 65435
rect 2717 65379 2773 65435
rect 2859 65379 2915 65435
rect 3001 65379 3057 65435
rect 3143 65379 3199 65435
rect 3285 65379 3341 65435
rect 3427 65379 3483 65435
rect 3569 65379 3625 65435
rect 3711 65379 3767 65435
rect 3853 65379 3909 65435
rect 3995 65379 4051 65435
rect 4137 65379 4193 65435
rect 4279 65379 4335 65435
rect 4421 65379 4477 65435
rect 4563 65379 4619 65435
rect 4705 65379 4761 65435
rect 4847 65379 4903 65435
rect 4989 65379 5045 65435
rect 5131 65379 5187 65435
rect 5273 65379 5329 65435
rect 5415 65379 5471 65435
rect 5557 65379 5613 65435
rect 5699 65379 5755 65435
rect 5841 65379 5897 65435
rect 5983 65379 6039 65435
rect 6125 65379 6181 65435
rect 6267 65379 6323 65435
rect 6409 65379 6465 65435
rect 6551 65379 6607 65435
rect 6693 65379 6749 65435
rect 6835 65379 6891 65435
rect 6977 65379 7033 65435
rect 7119 65379 7175 65435
rect 7261 65379 7317 65435
rect 7403 65379 7459 65435
rect 7545 65379 7601 65435
rect 7687 65379 7743 65435
rect 7829 65379 7885 65435
rect 7971 65379 8027 65435
rect 8113 65379 8169 65435
rect 8255 65379 8311 65435
rect 8397 65379 8453 65435
rect 8539 65379 8595 65435
rect 8681 65379 8737 65435
rect 8823 65379 8879 65435
rect 8965 65379 9021 65435
rect 9107 65379 9163 65435
rect 9249 65379 9305 65435
rect 9391 65379 9447 65435
rect 9533 65379 9589 65435
rect 9675 65379 9731 65435
rect 9817 65379 9873 65435
rect 9959 65379 10015 65435
rect 10101 65379 10157 65435
rect 10243 65379 10299 65435
rect 10385 65379 10441 65435
rect 10527 65379 10583 65435
rect 10669 65379 10725 65435
rect 10811 65379 10867 65435
rect 10953 65379 11009 65435
rect 11095 65379 11151 65435
rect 11237 65379 11293 65435
rect 11379 65379 11435 65435
rect 11521 65379 11577 65435
rect 11663 65379 11719 65435
rect 11805 65379 11861 65435
rect 11947 65379 12003 65435
rect 12089 65379 12145 65435
rect 12231 65379 12287 65435
rect 12373 65379 12429 65435
rect 12515 65379 12571 65435
rect 12657 65379 12713 65435
rect 12799 65379 12855 65435
rect 12941 65379 12997 65435
rect 13083 65379 13139 65435
rect 13225 65379 13281 65435
rect 13367 65379 13423 65435
rect 13509 65379 13565 65435
rect 13651 65379 13707 65435
rect 13793 65379 13849 65435
rect 13935 65379 13991 65435
rect 14077 65379 14133 65435
rect 14219 65379 14275 65435
rect 14361 65379 14417 65435
rect 14503 65379 14559 65435
rect 14645 65379 14701 65435
rect 14787 65379 14843 65435
rect 161 65237 217 65293
rect 303 65237 359 65293
rect 445 65237 501 65293
rect 587 65237 643 65293
rect 729 65237 785 65293
rect 871 65237 927 65293
rect 1013 65237 1069 65293
rect 1155 65237 1211 65293
rect 1297 65237 1353 65293
rect 1439 65237 1495 65293
rect 1581 65237 1637 65293
rect 1723 65237 1779 65293
rect 1865 65237 1921 65293
rect 2007 65237 2063 65293
rect 2149 65237 2205 65293
rect 2291 65237 2347 65293
rect 2433 65237 2489 65293
rect 2575 65237 2631 65293
rect 2717 65237 2773 65293
rect 2859 65237 2915 65293
rect 3001 65237 3057 65293
rect 3143 65237 3199 65293
rect 3285 65237 3341 65293
rect 3427 65237 3483 65293
rect 3569 65237 3625 65293
rect 3711 65237 3767 65293
rect 3853 65237 3909 65293
rect 3995 65237 4051 65293
rect 4137 65237 4193 65293
rect 4279 65237 4335 65293
rect 4421 65237 4477 65293
rect 4563 65237 4619 65293
rect 4705 65237 4761 65293
rect 4847 65237 4903 65293
rect 4989 65237 5045 65293
rect 5131 65237 5187 65293
rect 5273 65237 5329 65293
rect 5415 65237 5471 65293
rect 5557 65237 5613 65293
rect 5699 65237 5755 65293
rect 5841 65237 5897 65293
rect 5983 65237 6039 65293
rect 6125 65237 6181 65293
rect 6267 65237 6323 65293
rect 6409 65237 6465 65293
rect 6551 65237 6607 65293
rect 6693 65237 6749 65293
rect 6835 65237 6891 65293
rect 6977 65237 7033 65293
rect 7119 65237 7175 65293
rect 7261 65237 7317 65293
rect 7403 65237 7459 65293
rect 7545 65237 7601 65293
rect 7687 65237 7743 65293
rect 7829 65237 7885 65293
rect 7971 65237 8027 65293
rect 8113 65237 8169 65293
rect 8255 65237 8311 65293
rect 8397 65237 8453 65293
rect 8539 65237 8595 65293
rect 8681 65237 8737 65293
rect 8823 65237 8879 65293
rect 8965 65237 9021 65293
rect 9107 65237 9163 65293
rect 9249 65237 9305 65293
rect 9391 65237 9447 65293
rect 9533 65237 9589 65293
rect 9675 65237 9731 65293
rect 9817 65237 9873 65293
rect 9959 65237 10015 65293
rect 10101 65237 10157 65293
rect 10243 65237 10299 65293
rect 10385 65237 10441 65293
rect 10527 65237 10583 65293
rect 10669 65237 10725 65293
rect 10811 65237 10867 65293
rect 10953 65237 11009 65293
rect 11095 65237 11151 65293
rect 11237 65237 11293 65293
rect 11379 65237 11435 65293
rect 11521 65237 11577 65293
rect 11663 65237 11719 65293
rect 11805 65237 11861 65293
rect 11947 65237 12003 65293
rect 12089 65237 12145 65293
rect 12231 65237 12287 65293
rect 12373 65237 12429 65293
rect 12515 65237 12571 65293
rect 12657 65237 12713 65293
rect 12799 65237 12855 65293
rect 12941 65237 12997 65293
rect 13083 65237 13139 65293
rect 13225 65237 13281 65293
rect 13367 65237 13423 65293
rect 13509 65237 13565 65293
rect 13651 65237 13707 65293
rect 13793 65237 13849 65293
rect 13935 65237 13991 65293
rect 14077 65237 14133 65293
rect 14219 65237 14275 65293
rect 14361 65237 14417 65293
rect 14503 65237 14559 65293
rect 14645 65237 14701 65293
rect 14787 65237 14843 65293
rect 161 64907 217 64963
rect 303 64907 359 64963
rect 445 64907 501 64963
rect 587 64907 643 64963
rect 729 64907 785 64963
rect 871 64907 927 64963
rect 1013 64907 1069 64963
rect 1155 64907 1211 64963
rect 1297 64907 1353 64963
rect 1439 64907 1495 64963
rect 1581 64907 1637 64963
rect 1723 64907 1779 64963
rect 1865 64907 1921 64963
rect 2007 64907 2063 64963
rect 2149 64907 2205 64963
rect 2291 64907 2347 64963
rect 2433 64907 2489 64963
rect 2575 64907 2631 64963
rect 2717 64907 2773 64963
rect 2859 64907 2915 64963
rect 3001 64907 3057 64963
rect 3143 64907 3199 64963
rect 3285 64907 3341 64963
rect 3427 64907 3483 64963
rect 3569 64907 3625 64963
rect 3711 64907 3767 64963
rect 3853 64907 3909 64963
rect 3995 64907 4051 64963
rect 4137 64907 4193 64963
rect 4279 64907 4335 64963
rect 4421 64907 4477 64963
rect 4563 64907 4619 64963
rect 4705 64907 4761 64963
rect 4847 64907 4903 64963
rect 4989 64907 5045 64963
rect 5131 64907 5187 64963
rect 5273 64907 5329 64963
rect 5415 64907 5471 64963
rect 5557 64907 5613 64963
rect 5699 64907 5755 64963
rect 5841 64907 5897 64963
rect 5983 64907 6039 64963
rect 6125 64907 6181 64963
rect 6267 64907 6323 64963
rect 6409 64907 6465 64963
rect 6551 64907 6607 64963
rect 6693 64907 6749 64963
rect 6835 64907 6891 64963
rect 6977 64907 7033 64963
rect 7119 64907 7175 64963
rect 7261 64907 7317 64963
rect 7403 64907 7459 64963
rect 7545 64907 7601 64963
rect 7687 64907 7743 64963
rect 7829 64907 7885 64963
rect 7971 64907 8027 64963
rect 8113 64907 8169 64963
rect 8255 64907 8311 64963
rect 8397 64907 8453 64963
rect 8539 64907 8595 64963
rect 8681 64907 8737 64963
rect 8823 64907 8879 64963
rect 8965 64907 9021 64963
rect 9107 64907 9163 64963
rect 9249 64907 9305 64963
rect 9391 64907 9447 64963
rect 9533 64907 9589 64963
rect 9675 64907 9731 64963
rect 9817 64907 9873 64963
rect 9959 64907 10015 64963
rect 10101 64907 10157 64963
rect 10243 64907 10299 64963
rect 10385 64907 10441 64963
rect 10527 64907 10583 64963
rect 10669 64907 10725 64963
rect 10811 64907 10867 64963
rect 10953 64907 11009 64963
rect 11095 64907 11151 64963
rect 11237 64907 11293 64963
rect 11379 64907 11435 64963
rect 11521 64907 11577 64963
rect 11663 64907 11719 64963
rect 11805 64907 11861 64963
rect 11947 64907 12003 64963
rect 12089 64907 12145 64963
rect 12231 64907 12287 64963
rect 12373 64907 12429 64963
rect 12515 64907 12571 64963
rect 12657 64907 12713 64963
rect 12799 64907 12855 64963
rect 12941 64907 12997 64963
rect 13083 64907 13139 64963
rect 13225 64907 13281 64963
rect 13367 64907 13423 64963
rect 13509 64907 13565 64963
rect 13651 64907 13707 64963
rect 13793 64907 13849 64963
rect 13935 64907 13991 64963
rect 14077 64907 14133 64963
rect 14219 64907 14275 64963
rect 14361 64907 14417 64963
rect 14503 64907 14559 64963
rect 14645 64907 14701 64963
rect 14787 64907 14843 64963
rect 161 64765 217 64821
rect 303 64765 359 64821
rect 445 64765 501 64821
rect 587 64765 643 64821
rect 729 64765 785 64821
rect 871 64765 927 64821
rect 1013 64765 1069 64821
rect 1155 64765 1211 64821
rect 1297 64765 1353 64821
rect 1439 64765 1495 64821
rect 1581 64765 1637 64821
rect 1723 64765 1779 64821
rect 1865 64765 1921 64821
rect 2007 64765 2063 64821
rect 2149 64765 2205 64821
rect 2291 64765 2347 64821
rect 2433 64765 2489 64821
rect 2575 64765 2631 64821
rect 2717 64765 2773 64821
rect 2859 64765 2915 64821
rect 3001 64765 3057 64821
rect 3143 64765 3199 64821
rect 3285 64765 3341 64821
rect 3427 64765 3483 64821
rect 3569 64765 3625 64821
rect 3711 64765 3767 64821
rect 3853 64765 3909 64821
rect 3995 64765 4051 64821
rect 4137 64765 4193 64821
rect 4279 64765 4335 64821
rect 4421 64765 4477 64821
rect 4563 64765 4619 64821
rect 4705 64765 4761 64821
rect 4847 64765 4903 64821
rect 4989 64765 5045 64821
rect 5131 64765 5187 64821
rect 5273 64765 5329 64821
rect 5415 64765 5471 64821
rect 5557 64765 5613 64821
rect 5699 64765 5755 64821
rect 5841 64765 5897 64821
rect 5983 64765 6039 64821
rect 6125 64765 6181 64821
rect 6267 64765 6323 64821
rect 6409 64765 6465 64821
rect 6551 64765 6607 64821
rect 6693 64765 6749 64821
rect 6835 64765 6891 64821
rect 6977 64765 7033 64821
rect 7119 64765 7175 64821
rect 7261 64765 7317 64821
rect 7403 64765 7459 64821
rect 7545 64765 7601 64821
rect 7687 64765 7743 64821
rect 7829 64765 7885 64821
rect 7971 64765 8027 64821
rect 8113 64765 8169 64821
rect 8255 64765 8311 64821
rect 8397 64765 8453 64821
rect 8539 64765 8595 64821
rect 8681 64765 8737 64821
rect 8823 64765 8879 64821
rect 8965 64765 9021 64821
rect 9107 64765 9163 64821
rect 9249 64765 9305 64821
rect 9391 64765 9447 64821
rect 9533 64765 9589 64821
rect 9675 64765 9731 64821
rect 9817 64765 9873 64821
rect 9959 64765 10015 64821
rect 10101 64765 10157 64821
rect 10243 64765 10299 64821
rect 10385 64765 10441 64821
rect 10527 64765 10583 64821
rect 10669 64765 10725 64821
rect 10811 64765 10867 64821
rect 10953 64765 11009 64821
rect 11095 64765 11151 64821
rect 11237 64765 11293 64821
rect 11379 64765 11435 64821
rect 11521 64765 11577 64821
rect 11663 64765 11719 64821
rect 11805 64765 11861 64821
rect 11947 64765 12003 64821
rect 12089 64765 12145 64821
rect 12231 64765 12287 64821
rect 12373 64765 12429 64821
rect 12515 64765 12571 64821
rect 12657 64765 12713 64821
rect 12799 64765 12855 64821
rect 12941 64765 12997 64821
rect 13083 64765 13139 64821
rect 13225 64765 13281 64821
rect 13367 64765 13423 64821
rect 13509 64765 13565 64821
rect 13651 64765 13707 64821
rect 13793 64765 13849 64821
rect 13935 64765 13991 64821
rect 14077 64765 14133 64821
rect 14219 64765 14275 64821
rect 14361 64765 14417 64821
rect 14503 64765 14559 64821
rect 14645 64765 14701 64821
rect 14787 64765 14843 64821
rect 161 64623 217 64679
rect 303 64623 359 64679
rect 445 64623 501 64679
rect 587 64623 643 64679
rect 729 64623 785 64679
rect 871 64623 927 64679
rect 1013 64623 1069 64679
rect 1155 64623 1211 64679
rect 1297 64623 1353 64679
rect 1439 64623 1495 64679
rect 1581 64623 1637 64679
rect 1723 64623 1779 64679
rect 1865 64623 1921 64679
rect 2007 64623 2063 64679
rect 2149 64623 2205 64679
rect 2291 64623 2347 64679
rect 2433 64623 2489 64679
rect 2575 64623 2631 64679
rect 2717 64623 2773 64679
rect 2859 64623 2915 64679
rect 3001 64623 3057 64679
rect 3143 64623 3199 64679
rect 3285 64623 3341 64679
rect 3427 64623 3483 64679
rect 3569 64623 3625 64679
rect 3711 64623 3767 64679
rect 3853 64623 3909 64679
rect 3995 64623 4051 64679
rect 4137 64623 4193 64679
rect 4279 64623 4335 64679
rect 4421 64623 4477 64679
rect 4563 64623 4619 64679
rect 4705 64623 4761 64679
rect 4847 64623 4903 64679
rect 4989 64623 5045 64679
rect 5131 64623 5187 64679
rect 5273 64623 5329 64679
rect 5415 64623 5471 64679
rect 5557 64623 5613 64679
rect 5699 64623 5755 64679
rect 5841 64623 5897 64679
rect 5983 64623 6039 64679
rect 6125 64623 6181 64679
rect 6267 64623 6323 64679
rect 6409 64623 6465 64679
rect 6551 64623 6607 64679
rect 6693 64623 6749 64679
rect 6835 64623 6891 64679
rect 6977 64623 7033 64679
rect 7119 64623 7175 64679
rect 7261 64623 7317 64679
rect 7403 64623 7459 64679
rect 7545 64623 7601 64679
rect 7687 64623 7743 64679
rect 7829 64623 7885 64679
rect 7971 64623 8027 64679
rect 8113 64623 8169 64679
rect 8255 64623 8311 64679
rect 8397 64623 8453 64679
rect 8539 64623 8595 64679
rect 8681 64623 8737 64679
rect 8823 64623 8879 64679
rect 8965 64623 9021 64679
rect 9107 64623 9163 64679
rect 9249 64623 9305 64679
rect 9391 64623 9447 64679
rect 9533 64623 9589 64679
rect 9675 64623 9731 64679
rect 9817 64623 9873 64679
rect 9959 64623 10015 64679
rect 10101 64623 10157 64679
rect 10243 64623 10299 64679
rect 10385 64623 10441 64679
rect 10527 64623 10583 64679
rect 10669 64623 10725 64679
rect 10811 64623 10867 64679
rect 10953 64623 11009 64679
rect 11095 64623 11151 64679
rect 11237 64623 11293 64679
rect 11379 64623 11435 64679
rect 11521 64623 11577 64679
rect 11663 64623 11719 64679
rect 11805 64623 11861 64679
rect 11947 64623 12003 64679
rect 12089 64623 12145 64679
rect 12231 64623 12287 64679
rect 12373 64623 12429 64679
rect 12515 64623 12571 64679
rect 12657 64623 12713 64679
rect 12799 64623 12855 64679
rect 12941 64623 12997 64679
rect 13083 64623 13139 64679
rect 13225 64623 13281 64679
rect 13367 64623 13423 64679
rect 13509 64623 13565 64679
rect 13651 64623 13707 64679
rect 13793 64623 13849 64679
rect 13935 64623 13991 64679
rect 14077 64623 14133 64679
rect 14219 64623 14275 64679
rect 14361 64623 14417 64679
rect 14503 64623 14559 64679
rect 14645 64623 14701 64679
rect 14787 64623 14843 64679
rect 161 64481 217 64537
rect 303 64481 359 64537
rect 445 64481 501 64537
rect 587 64481 643 64537
rect 729 64481 785 64537
rect 871 64481 927 64537
rect 1013 64481 1069 64537
rect 1155 64481 1211 64537
rect 1297 64481 1353 64537
rect 1439 64481 1495 64537
rect 1581 64481 1637 64537
rect 1723 64481 1779 64537
rect 1865 64481 1921 64537
rect 2007 64481 2063 64537
rect 2149 64481 2205 64537
rect 2291 64481 2347 64537
rect 2433 64481 2489 64537
rect 2575 64481 2631 64537
rect 2717 64481 2773 64537
rect 2859 64481 2915 64537
rect 3001 64481 3057 64537
rect 3143 64481 3199 64537
rect 3285 64481 3341 64537
rect 3427 64481 3483 64537
rect 3569 64481 3625 64537
rect 3711 64481 3767 64537
rect 3853 64481 3909 64537
rect 3995 64481 4051 64537
rect 4137 64481 4193 64537
rect 4279 64481 4335 64537
rect 4421 64481 4477 64537
rect 4563 64481 4619 64537
rect 4705 64481 4761 64537
rect 4847 64481 4903 64537
rect 4989 64481 5045 64537
rect 5131 64481 5187 64537
rect 5273 64481 5329 64537
rect 5415 64481 5471 64537
rect 5557 64481 5613 64537
rect 5699 64481 5755 64537
rect 5841 64481 5897 64537
rect 5983 64481 6039 64537
rect 6125 64481 6181 64537
rect 6267 64481 6323 64537
rect 6409 64481 6465 64537
rect 6551 64481 6607 64537
rect 6693 64481 6749 64537
rect 6835 64481 6891 64537
rect 6977 64481 7033 64537
rect 7119 64481 7175 64537
rect 7261 64481 7317 64537
rect 7403 64481 7459 64537
rect 7545 64481 7601 64537
rect 7687 64481 7743 64537
rect 7829 64481 7885 64537
rect 7971 64481 8027 64537
rect 8113 64481 8169 64537
rect 8255 64481 8311 64537
rect 8397 64481 8453 64537
rect 8539 64481 8595 64537
rect 8681 64481 8737 64537
rect 8823 64481 8879 64537
rect 8965 64481 9021 64537
rect 9107 64481 9163 64537
rect 9249 64481 9305 64537
rect 9391 64481 9447 64537
rect 9533 64481 9589 64537
rect 9675 64481 9731 64537
rect 9817 64481 9873 64537
rect 9959 64481 10015 64537
rect 10101 64481 10157 64537
rect 10243 64481 10299 64537
rect 10385 64481 10441 64537
rect 10527 64481 10583 64537
rect 10669 64481 10725 64537
rect 10811 64481 10867 64537
rect 10953 64481 11009 64537
rect 11095 64481 11151 64537
rect 11237 64481 11293 64537
rect 11379 64481 11435 64537
rect 11521 64481 11577 64537
rect 11663 64481 11719 64537
rect 11805 64481 11861 64537
rect 11947 64481 12003 64537
rect 12089 64481 12145 64537
rect 12231 64481 12287 64537
rect 12373 64481 12429 64537
rect 12515 64481 12571 64537
rect 12657 64481 12713 64537
rect 12799 64481 12855 64537
rect 12941 64481 12997 64537
rect 13083 64481 13139 64537
rect 13225 64481 13281 64537
rect 13367 64481 13423 64537
rect 13509 64481 13565 64537
rect 13651 64481 13707 64537
rect 13793 64481 13849 64537
rect 13935 64481 13991 64537
rect 14077 64481 14133 64537
rect 14219 64481 14275 64537
rect 14361 64481 14417 64537
rect 14503 64481 14559 64537
rect 14645 64481 14701 64537
rect 14787 64481 14843 64537
rect 161 64339 217 64395
rect 303 64339 359 64395
rect 445 64339 501 64395
rect 587 64339 643 64395
rect 729 64339 785 64395
rect 871 64339 927 64395
rect 1013 64339 1069 64395
rect 1155 64339 1211 64395
rect 1297 64339 1353 64395
rect 1439 64339 1495 64395
rect 1581 64339 1637 64395
rect 1723 64339 1779 64395
rect 1865 64339 1921 64395
rect 2007 64339 2063 64395
rect 2149 64339 2205 64395
rect 2291 64339 2347 64395
rect 2433 64339 2489 64395
rect 2575 64339 2631 64395
rect 2717 64339 2773 64395
rect 2859 64339 2915 64395
rect 3001 64339 3057 64395
rect 3143 64339 3199 64395
rect 3285 64339 3341 64395
rect 3427 64339 3483 64395
rect 3569 64339 3625 64395
rect 3711 64339 3767 64395
rect 3853 64339 3909 64395
rect 3995 64339 4051 64395
rect 4137 64339 4193 64395
rect 4279 64339 4335 64395
rect 4421 64339 4477 64395
rect 4563 64339 4619 64395
rect 4705 64339 4761 64395
rect 4847 64339 4903 64395
rect 4989 64339 5045 64395
rect 5131 64339 5187 64395
rect 5273 64339 5329 64395
rect 5415 64339 5471 64395
rect 5557 64339 5613 64395
rect 5699 64339 5755 64395
rect 5841 64339 5897 64395
rect 5983 64339 6039 64395
rect 6125 64339 6181 64395
rect 6267 64339 6323 64395
rect 6409 64339 6465 64395
rect 6551 64339 6607 64395
rect 6693 64339 6749 64395
rect 6835 64339 6891 64395
rect 6977 64339 7033 64395
rect 7119 64339 7175 64395
rect 7261 64339 7317 64395
rect 7403 64339 7459 64395
rect 7545 64339 7601 64395
rect 7687 64339 7743 64395
rect 7829 64339 7885 64395
rect 7971 64339 8027 64395
rect 8113 64339 8169 64395
rect 8255 64339 8311 64395
rect 8397 64339 8453 64395
rect 8539 64339 8595 64395
rect 8681 64339 8737 64395
rect 8823 64339 8879 64395
rect 8965 64339 9021 64395
rect 9107 64339 9163 64395
rect 9249 64339 9305 64395
rect 9391 64339 9447 64395
rect 9533 64339 9589 64395
rect 9675 64339 9731 64395
rect 9817 64339 9873 64395
rect 9959 64339 10015 64395
rect 10101 64339 10157 64395
rect 10243 64339 10299 64395
rect 10385 64339 10441 64395
rect 10527 64339 10583 64395
rect 10669 64339 10725 64395
rect 10811 64339 10867 64395
rect 10953 64339 11009 64395
rect 11095 64339 11151 64395
rect 11237 64339 11293 64395
rect 11379 64339 11435 64395
rect 11521 64339 11577 64395
rect 11663 64339 11719 64395
rect 11805 64339 11861 64395
rect 11947 64339 12003 64395
rect 12089 64339 12145 64395
rect 12231 64339 12287 64395
rect 12373 64339 12429 64395
rect 12515 64339 12571 64395
rect 12657 64339 12713 64395
rect 12799 64339 12855 64395
rect 12941 64339 12997 64395
rect 13083 64339 13139 64395
rect 13225 64339 13281 64395
rect 13367 64339 13423 64395
rect 13509 64339 13565 64395
rect 13651 64339 13707 64395
rect 13793 64339 13849 64395
rect 13935 64339 13991 64395
rect 14077 64339 14133 64395
rect 14219 64339 14275 64395
rect 14361 64339 14417 64395
rect 14503 64339 14559 64395
rect 14645 64339 14701 64395
rect 14787 64339 14843 64395
rect 161 64197 217 64253
rect 303 64197 359 64253
rect 445 64197 501 64253
rect 587 64197 643 64253
rect 729 64197 785 64253
rect 871 64197 927 64253
rect 1013 64197 1069 64253
rect 1155 64197 1211 64253
rect 1297 64197 1353 64253
rect 1439 64197 1495 64253
rect 1581 64197 1637 64253
rect 1723 64197 1779 64253
rect 1865 64197 1921 64253
rect 2007 64197 2063 64253
rect 2149 64197 2205 64253
rect 2291 64197 2347 64253
rect 2433 64197 2489 64253
rect 2575 64197 2631 64253
rect 2717 64197 2773 64253
rect 2859 64197 2915 64253
rect 3001 64197 3057 64253
rect 3143 64197 3199 64253
rect 3285 64197 3341 64253
rect 3427 64197 3483 64253
rect 3569 64197 3625 64253
rect 3711 64197 3767 64253
rect 3853 64197 3909 64253
rect 3995 64197 4051 64253
rect 4137 64197 4193 64253
rect 4279 64197 4335 64253
rect 4421 64197 4477 64253
rect 4563 64197 4619 64253
rect 4705 64197 4761 64253
rect 4847 64197 4903 64253
rect 4989 64197 5045 64253
rect 5131 64197 5187 64253
rect 5273 64197 5329 64253
rect 5415 64197 5471 64253
rect 5557 64197 5613 64253
rect 5699 64197 5755 64253
rect 5841 64197 5897 64253
rect 5983 64197 6039 64253
rect 6125 64197 6181 64253
rect 6267 64197 6323 64253
rect 6409 64197 6465 64253
rect 6551 64197 6607 64253
rect 6693 64197 6749 64253
rect 6835 64197 6891 64253
rect 6977 64197 7033 64253
rect 7119 64197 7175 64253
rect 7261 64197 7317 64253
rect 7403 64197 7459 64253
rect 7545 64197 7601 64253
rect 7687 64197 7743 64253
rect 7829 64197 7885 64253
rect 7971 64197 8027 64253
rect 8113 64197 8169 64253
rect 8255 64197 8311 64253
rect 8397 64197 8453 64253
rect 8539 64197 8595 64253
rect 8681 64197 8737 64253
rect 8823 64197 8879 64253
rect 8965 64197 9021 64253
rect 9107 64197 9163 64253
rect 9249 64197 9305 64253
rect 9391 64197 9447 64253
rect 9533 64197 9589 64253
rect 9675 64197 9731 64253
rect 9817 64197 9873 64253
rect 9959 64197 10015 64253
rect 10101 64197 10157 64253
rect 10243 64197 10299 64253
rect 10385 64197 10441 64253
rect 10527 64197 10583 64253
rect 10669 64197 10725 64253
rect 10811 64197 10867 64253
rect 10953 64197 11009 64253
rect 11095 64197 11151 64253
rect 11237 64197 11293 64253
rect 11379 64197 11435 64253
rect 11521 64197 11577 64253
rect 11663 64197 11719 64253
rect 11805 64197 11861 64253
rect 11947 64197 12003 64253
rect 12089 64197 12145 64253
rect 12231 64197 12287 64253
rect 12373 64197 12429 64253
rect 12515 64197 12571 64253
rect 12657 64197 12713 64253
rect 12799 64197 12855 64253
rect 12941 64197 12997 64253
rect 13083 64197 13139 64253
rect 13225 64197 13281 64253
rect 13367 64197 13423 64253
rect 13509 64197 13565 64253
rect 13651 64197 13707 64253
rect 13793 64197 13849 64253
rect 13935 64197 13991 64253
rect 14077 64197 14133 64253
rect 14219 64197 14275 64253
rect 14361 64197 14417 64253
rect 14503 64197 14559 64253
rect 14645 64197 14701 64253
rect 14787 64197 14843 64253
rect 161 64055 217 64111
rect 303 64055 359 64111
rect 445 64055 501 64111
rect 587 64055 643 64111
rect 729 64055 785 64111
rect 871 64055 927 64111
rect 1013 64055 1069 64111
rect 1155 64055 1211 64111
rect 1297 64055 1353 64111
rect 1439 64055 1495 64111
rect 1581 64055 1637 64111
rect 1723 64055 1779 64111
rect 1865 64055 1921 64111
rect 2007 64055 2063 64111
rect 2149 64055 2205 64111
rect 2291 64055 2347 64111
rect 2433 64055 2489 64111
rect 2575 64055 2631 64111
rect 2717 64055 2773 64111
rect 2859 64055 2915 64111
rect 3001 64055 3057 64111
rect 3143 64055 3199 64111
rect 3285 64055 3341 64111
rect 3427 64055 3483 64111
rect 3569 64055 3625 64111
rect 3711 64055 3767 64111
rect 3853 64055 3909 64111
rect 3995 64055 4051 64111
rect 4137 64055 4193 64111
rect 4279 64055 4335 64111
rect 4421 64055 4477 64111
rect 4563 64055 4619 64111
rect 4705 64055 4761 64111
rect 4847 64055 4903 64111
rect 4989 64055 5045 64111
rect 5131 64055 5187 64111
rect 5273 64055 5329 64111
rect 5415 64055 5471 64111
rect 5557 64055 5613 64111
rect 5699 64055 5755 64111
rect 5841 64055 5897 64111
rect 5983 64055 6039 64111
rect 6125 64055 6181 64111
rect 6267 64055 6323 64111
rect 6409 64055 6465 64111
rect 6551 64055 6607 64111
rect 6693 64055 6749 64111
rect 6835 64055 6891 64111
rect 6977 64055 7033 64111
rect 7119 64055 7175 64111
rect 7261 64055 7317 64111
rect 7403 64055 7459 64111
rect 7545 64055 7601 64111
rect 7687 64055 7743 64111
rect 7829 64055 7885 64111
rect 7971 64055 8027 64111
rect 8113 64055 8169 64111
rect 8255 64055 8311 64111
rect 8397 64055 8453 64111
rect 8539 64055 8595 64111
rect 8681 64055 8737 64111
rect 8823 64055 8879 64111
rect 8965 64055 9021 64111
rect 9107 64055 9163 64111
rect 9249 64055 9305 64111
rect 9391 64055 9447 64111
rect 9533 64055 9589 64111
rect 9675 64055 9731 64111
rect 9817 64055 9873 64111
rect 9959 64055 10015 64111
rect 10101 64055 10157 64111
rect 10243 64055 10299 64111
rect 10385 64055 10441 64111
rect 10527 64055 10583 64111
rect 10669 64055 10725 64111
rect 10811 64055 10867 64111
rect 10953 64055 11009 64111
rect 11095 64055 11151 64111
rect 11237 64055 11293 64111
rect 11379 64055 11435 64111
rect 11521 64055 11577 64111
rect 11663 64055 11719 64111
rect 11805 64055 11861 64111
rect 11947 64055 12003 64111
rect 12089 64055 12145 64111
rect 12231 64055 12287 64111
rect 12373 64055 12429 64111
rect 12515 64055 12571 64111
rect 12657 64055 12713 64111
rect 12799 64055 12855 64111
rect 12941 64055 12997 64111
rect 13083 64055 13139 64111
rect 13225 64055 13281 64111
rect 13367 64055 13423 64111
rect 13509 64055 13565 64111
rect 13651 64055 13707 64111
rect 13793 64055 13849 64111
rect 13935 64055 13991 64111
rect 14077 64055 14133 64111
rect 14219 64055 14275 64111
rect 14361 64055 14417 64111
rect 14503 64055 14559 64111
rect 14645 64055 14701 64111
rect 14787 64055 14843 64111
rect 161 63913 217 63969
rect 303 63913 359 63969
rect 445 63913 501 63969
rect 587 63913 643 63969
rect 729 63913 785 63969
rect 871 63913 927 63969
rect 1013 63913 1069 63969
rect 1155 63913 1211 63969
rect 1297 63913 1353 63969
rect 1439 63913 1495 63969
rect 1581 63913 1637 63969
rect 1723 63913 1779 63969
rect 1865 63913 1921 63969
rect 2007 63913 2063 63969
rect 2149 63913 2205 63969
rect 2291 63913 2347 63969
rect 2433 63913 2489 63969
rect 2575 63913 2631 63969
rect 2717 63913 2773 63969
rect 2859 63913 2915 63969
rect 3001 63913 3057 63969
rect 3143 63913 3199 63969
rect 3285 63913 3341 63969
rect 3427 63913 3483 63969
rect 3569 63913 3625 63969
rect 3711 63913 3767 63969
rect 3853 63913 3909 63969
rect 3995 63913 4051 63969
rect 4137 63913 4193 63969
rect 4279 63913 4335 63969
rect 4421 63913 4477 63969
rect 4563 63913 4619 63969
rect 4705 63913 4761 63969
rect 4847 63913 4903 63969
rect 4989 63913 5045 63969
rect 5131 63913 5187 63969
rect 5273 63913 5329 63969
rect 5415 63913 5471 63969
rect 5557 63913 5613 63969
rect 5699 63913 5755 63969
rect 5841 63913 5897 63969
rect 5983 63913 6039 63969
rect 6125 63913 6181 63969
rect 6267 63913 6323 63969
rect 6409 63913 6465 63969
rect 6551 63913 6607 63969
rect 6693 63913 6749 63969
rect 6835 63913 6891 63969
rect 6977 63913 7033 63969
rect 7119 63913 7175 63969
rect 7261 63913 7317 63969
rect 7403 63913 7459 63969
rect 7545 63913 7601 63969
rect 7687 63913 7743 63969
rect 7829 63913 7885 63969
rect 7971 63913 8027 63969
rect 8113 63913 8169 63969
rect 8255 63913 8311 63969
rect 8397 63913 8453 63969
rect 8539 63913 8595 63969
rect 8681 63913 8737 63969
rect 8823 63913 8879 63969
rect 8965 63913 9021 63969
rect 9107 63913 9163 63969
rect 9249 63913 9305 63969
rect 9391 63913 9447 63969
rect 9533 63913 9589 63969
rect 9675 63913 9731 63969
rect 9817 63913 9873 63969
rect 9959 63913 10015 63969
rect 10101 63913 10157 63969
rect 10243 63913 10299 63969
rect 10385 63913 10441 63969
rect 10527 63913 10583 63969
rect 10669 63913 10725 63969
rect 10811 63913 10867 63969
rect 10953 63913 11009 63969
rect 11095 63913 11151 63969
rect 11237 63913 11293 63969
rect 11379 63913 11435 63969
rect 11521 63913 11577 63969
rect 11663 63913 11719 63969
rect 11805 63913 11861 63969
rect 11947 63913 12003 63969
rect 12089 63913 12145 63969
rect 12231 63913 12287 63969
rect 12373 63913 12429 63969
rect 12515 63913 12571 63969
rect 12657 63913 12713 63969
rect 12799 63913 12855 63969
rect 12941 63913 12997 63969
rect 13083 63913 13139 63969
rect 13225 63913 13281 63969
rect 13367 63913 13423 63969
rect 13509 63913 13565 63969
rect 13651 63913 13707 63969
rect 13793 63913 13849 63969
rect 13935 63913 13991 63969
rect 14077 63913 14133 63969
rect 14219 63913 14275 63969
rect 14361 63913 14417 63969
rect 14503 63913 14559 63969
rect 14645 63913 14701 63969
rect 14787 63913 14843 63969
rect 161 63771 217 63827
rect 303 63771 359 63827
rect 445 63771 501 63827
rect 587 63771 643 63827
rect 729 63771 785 63827
rect 871 63771 927 63827
rect 1013 63771 1069 63827
rect 1155 63771 1211 63827
rect 1297 63771 1353 63827
rect 1439 63771 1495 63827
rect 1581 63771 1637 63827
rect 1723 63771 1779 63827
rect 1865 63771 1921 63827
rect 2007 63771 2063 63827
rect 2149 63771 2205 63827
rect 2291 63771 2347 63827
rect 2433 63771 2489 63827
rect 2575 63771 2631 63827
rect 2717 63771 2773 63827
rect 2859 63771 2915 63827
rect 3001 63771 3057 63827
rect 3143 63771 3199 63827
rect 3285 63771 3341 63827
rect 3427 63771 3483 63827
rect 3569 63771 3625 63827
rect 3711 63771 3767 63827
rect 3853 63771 3909 63827
rect 3995 63771 4051 63827
rect 4137 63771 4193 63827
rect 4279 63771 4335 63827
rect 4421 63771 4477 63827
rect 4563 63771 4619 63827
rect 4705 63771 4761 63827
rect 4847 63771 4903 63827
rect 4989 63771 5045 63827
rect 5131 63771 5187 63827
rect 5273 63771 5329 63827
rect 5415 63771 5471 63827
rect 5557 63771 5613 63827
rect 5699 63771 5755 63827
rect 5841 63771 5897 63827
rect 5983 63771 6039 63827
rect 6125 63771 6181 63827
rect 6267 63771 6323 63827
rect 6409 63771 6465 63827
rect 6551 63771 6607 63827
rect 6693 63771 6749 63827
rect 6835 63771 6891 63827
rect 6977 63771 7033 63827
rect 7119 63771 7175 63827
rect 7261 63771 7317 63827
rect 7403 63771 7459 63827
rect 7545 63771 7601 63827
rect 7687 63771 7743 63827
rect 7829 63771 7885 63827
rect 7971 63771 8027 63827
rect 8113 63771 8169 63827
rect 8255 63771 8311 63827
rect 8397 63771 8453 63827
rect 8539 63771 8595 63827
rect 8681 63771 8737 63827
rect 8823 63771 8879 63827
rect 8965 63771 9021 63827
rect 9107 63771 9163 63827
rect 9249 63771 9305 63827
rect 9391 63771 9447 63827
rect 9533 63771 9589 63827
rect 9675 63771 9731 63827
rect 9817 63771 9873 63827
rect 9959 63771 10015 63827
rect 10101 63771 10157 63827
rect 10243 63771 10299 63827
rect 10385 63771 10441 63827
rect 10527 63771 10583 63827
rect 10669 63771 10725 63827
rect 10811 63771 10867 63827
rect 10953 63771 11009 63827
rect 11095 63771 11151 63827
rect 11237 63771 11293 63827
rect 11379 63771 11435 63827
rect 11521 63771 11577 63827
rect 11663 63771 11719 63827
rect 11805 63771 11861 63827
rect 11947 63771 12003 63827
rect 12089 63771 12145 63827
rect 12231 63771 12287 63827
rect 12373 63771 12429 63827
rect 12515 63771 12571 63827
rect 12657 63771 12713 63827
rect 12799 63771 12855 63827
rect 12941 63771 12997 63827
rect 13083 63771 13139 63827
rect 13225 63771 13281 63827
rect 13367 63771 13423 63827
rect 13509 63771 13565 63827
rect 13651 63771 13707 63827
rect 13793 63771 13849 63827
rect 13935 63771 13991 63827
rect 14077 63771 14133 63827
rect 14219 63771 14275 63827
rect 14361 63771 14417 63827
rect 14503 63771 14559 63827
rect 14645 63771 14701 63827
rect 14787 63771 14843 63827
rect 161 63629 217 63685
rect 303 63629 359 63685
rect 445 63629 501 63685
rect 587 63629 643 63685
rect 729 63629 785 63685
rect 871 63629 927 63685
rect 1013 63629 1069 63685
rect 1155 63629 1211 63685
rect 1297 63629 1353 63685
rect 1439 63629 1495 63685
rect 1581 63629 1637 63685
rect 1723 63629 1779 63685
rect 1865 63629 1921 63685
rect 2007 63629 2063 63685
rect 2149 63629 2205 63685
rect 2291 63629 2347 63685
rect 2433 63629 2489 63685
rect 2575 63629 2631 63685
rect 2717 63629 2773 63685
rect 2859 63629 2915 63685
rect 3001 63629 3057 63685
rect 3143 63629 3199 63685
rect 3285 63629 3341 63685
rect 3427 63629 3483 63685
rect 3569 63629 3625 63685
rect 3711 63629 3767 63685
rect 3853 63629 3909 63685
rect 3995 63629 4051 63685
rect 4137 63629 4193 63685
rect 4279 63629 4335 63685
rect 4421 63629 4477 63685
rect 4563 63629 4619 63685
rect 4705 63629 4761 63685
rect 4847 63629 4903 63685
rect 4989 63629 5045 63685
rect 5131 63629 5187 63685
rect 5273 63629 5329 63685
rect 5415 63629 5471 63685
rect 5557 63629 5613 63685
rect 5699 63629 5755 63685
rect 5841 63629 5897 63685
rect 5983 63629 6039 63685
rect 6125 63629 6181 63685
rect 6267 63629 6323 63685
rect 6409 63629 6465 63685
rect 6551 63629 6607 63685
rect 6693 63629 6749 63685
rect 6835 63629 6891 63685
rect 6977 63629 7033 63685
rect 7119 63629 7175 63685
rect 7261 63629 7317 63685
rect 7403 63629 7459 63685
rect 7545 63629 7601 63685
rect 7687 63629 7743 63685
rect 7829 63629 7885 63685
rect 7971 63629 8027 63685
rect 8113 63629 8169 63685
rect 8255 63629 8311 63685
rect 8397 63629 8453 63685
rect 8539 63629 8595 63685
rect 8681 63629 8737 63685
rect 8823 63629 8879 63685
rect 8965 63629 9021 63685
rect 9107 63629 9163 63685
rect 9249 63629 9305 63685
rect 9391 63629 9447 63685
rect 9533 63629 9589 63685
rect 9675 63629 9731 63685
rect 9817 63629 9873 63685
rect 9959 63629 10015 63685
rect 10101 63629 10157 63685
rect 10243 63629 10299 63685
rect 10385 63629 10441 63685
rect 10527 63629 10583 63685
rect 10669 63629 10725 63685
rect 10811 63629 10867 63685
rect 10953 63629 11009 63685
rect 11095 63629 11151 63685
rect 11237 63629 11293 63685
rect 11379 63629 11435 63685
rect 11521 63629 11577 63685
rect 11663 63629 11719 63685
rect 11805 63629 11861 63685
rect 11947 63629 12003 63685
rect 12089 63629 12145 63685
rect 12231 63629 12287 63685
rect 12373 63629 12429 63685
rect 12515 63629 12571 63685
rect 12657 63629 12713 63685
rect 12799 63629 12855 63685
rect 12941 63629 12997 63685
rect 13083 63629 13139 63685
rect 13225 63629 13281 63685
rect 13367 63629 13423 63685
rect 13509 63629 13565 63685
rect 13651 63629 13707 63685
rect 13793 63629 13849 63685
rect 13935 63629 13991 63685
rect 14077 63629 14133 63685
rect 14219 63629 14275 63685
rect 14361 63629 14417 63685
rect 14503 63629 14559 63685
rect 14645 63629 14701 63685
rect 14787 63629 14843 63685
rect 161 63315 217 63371
rect 303 63315 359 63371
rect 445 63315 501 63371
rect 587 63315 643 63371
rect 729 63315 785 63371
rect 871 63315 927 63371
rect 1013 63315 1069 63371
rect 1155 63315 1211 63371
rect 1297 63315 1353 63371
rect 1439 63315 1495 63371
rect 1581 63315 1637 63371
rect 1723 63315 1779 63371
rect 1865 63315 1921 63371
rect 2007 63315 2063 63371
rect 2149 63315 2205 63371
rect 2291 63315 2347 63371
rect 2433 63315 2489 63371
rect 2575 63315 2631 63371
rect 2717 63315 2773 63371
rect 2859 63315 2915 63371
rect 3001 63315 3057 63371
rect 3143 63315 3199 63371
rect 3285 63315 3341 63371
rect 3427 63315 3483 63371
rect 3569 63315 3625 63371
rect 3711 63315 3767 63371
rect 3853 63315 3909 63371
rect 3995 63315 4051 63371
rect 4137 63315 4193 63371
rect 4279 63315 4335 63371
rect 4421 63315 4477 63371
rect 4563 63315 4619 63371
rect 4705 63315 4761 63371
rect 4847 63315 4903 63371
rect 4989 63315 5045 63371
rect 5131 63315 5187 63371
rect 5273 63315 5329 63371
rect 5415 63315 5471 63371
rect 5557 63315 5613 63371
rect 5699 63315 5755 63371
rect 5841 63315 5897 63371
rect 5983 63315 6039 63371
rect 6125 63315 6181 63371
rect 6267 63315 6323 63371
rect 6409 63315 6465 63371
rect 6551 63315 6607 63371
rect 6693 63315 6749 63371
rect 6835 63315 6891 63371
rect 6977 63315 7033 63371
rect 7119 63315 7175 63371
rect 7261 63315 7317 63371
rect 7403 63315 7459 63371
rect 7545 63315 7601 63371
rect 7687 63315 7743 63371
rect 7829 63315 7885 63371
rect 7971 63315 8027 63371
rect 8113 63315 8169 63371
rect 8255 63315 8311 63371
rect 8397 63315 8453 63371
rect 8539 63315 8595 63371
rect 8681 63315 8737 63371
rect 8823 63315 8879 63371
rect 8965 63315 9021 63371
rect 9107 63315 9163 63371
rect 9249 63315 9305 63371
rect 9391 63315 9447 63371
rect 9533 63315 9589 63371
rect 9675 63315 9731 63371
rect 9817 63315 9873 63371
rect 9959 63315 10015 63371
rect 10101 63315 10157 63371
rect 10243 63315 10299 63371
rect 10385 63315 10441 63371
rect 10527 63315 10583 63371
rect 10669 63315 10725 63371
rect 10811 63315 10867 63371
rect 10953 63315 11009 63371
rect 11095 63315 11151 63371
rect 11237 63315 11293 63371
rect 11379 63315 11435 63371
rect 11521 63315 11577 63371
rect 11663 63315 11719 63371
rect 11805 63315 11861 63371
rect 11947 63315 12003 63371
rect 12089 63315 12145 63371
rect 12231 63315 12287 63371
rect 12373 63315 12429 63371
rect 12515 63315 12571 63371
rect 12657 63315 12713 63371
rect 12799 63315 12855 63371
rect 12941 63315 12997 63371
rect 13083 63315 13139 63371
rect 13225 63315 13281 63371
rect 13367 63315 13423 63371
rect 13509 63315 13565 63371
rect 13651 63315 13707 63371
rect 13793 63315 13849 63371
rect 13935 63315 13991 63371
rect 14077 63315 14133 63371
rect 14219 63315 14275 63371
rect 14361 63315 14417 63371
rect 14503 63315 14559 63371
rect 14645 63315 14701 63371
rect 14787 63315 14843 63371
rect 161 63173 217 63229
rect 303 63173 359 63229
rect 445 63173 501 63229
rect 587 63173 643 63229
rect 729 63173 785 63229
rect 871 63173 927 63229
rect 1013 63173 1069 63229
rect 1155 63173 1211 63229
rect 1297 63173 1353 63229
rect 1439 63173 1495 63229
rect 1581 63173 1637 63229
rect 1723 63173 1779 63229
rect 1865 63173 1921 63229
rect 2007 63173 2063 63229
rect 2149 63173 2205 63229
rect 2291 63173 2347 63229
rect 2433 63173 2489 63229
rect 2575 63173 2631 63229
rect 2717 63173 2773 63229
rect 2859 63173 2915 63229
rect 3001 63173 3057 63229
rect 3143 63173 3199 63229
rect 3285 63173 3341 63229
rect 3427 63173 3483 63229
rect 3569 63173 3625 63229
rect 3711 63173 3767 63229
rect 3853 63173 3909 63229
rect 3995 63173 4051 63229
rect 4137 63173 4193 63229
rect 4279 63173 4335 63229
rect 4421 63173 4477 63229
rect 4563 63173 4619 63229
rect 4705 63173 4761 63229
rect 4847 63173 4903 63229
rect 4989 63173 5045 63229
rect 5131 63173 5187 63229
rect 5273 63173 5329 63229
rect 5415 63173 5471 63229
rect 5557 63173 5613 63229
rect 5699 63173 5755 63229
rect 5841 63173 5897 63229
rect 5983 63173 6039 63229
rect 6125 63173 6181 63229
rect 6267 63173 6323 63229
rect 6409 63173 6465 63229
rect 6551 63173 6607 63229
rect 6693 63173 6749 63229
rect 6835 63173 6891 63229
rect 6977 63173 7033 63229
rect 7119 63173 7175 63229
rect 7261 63173 7317 63229
rect 7403 63173 7459 63229
rect 7545 63173 7601 63229
rect 7687 63173 7743 63229
rect 7829 63173 7885 63229
rect 7971 63173 8027 63229
rect 8113 63173 8169 63229
rect 8255 63173 8311 63229
rect 8397 63173 8453 63229
rect 8539 63173 8595 63229
rect 8681 63173 8737 63229
rect 8823 63173 8879 63229
rect 8965 63173 9021 63229
rect 9107 63173 9163 63229
rect 9249 63173 9305 63229
rect 9391 63173 9447 63229
rect 9533 63173 9589 63229
rect 9675 63173 9731 63229
rect 9817 63173 9873 63229
rect 9959 63173 10015 63229
rect 10101 63173 10157 63229
rect 10243 63173 10299 63229
rect 10385 63173 10441 63229
rect 10527 63173 10583 63229
rect 10669 63173 10725 63229
rect 10811 63173 10867 63229
rect 10953 63173 11009 63229
rect 11095 63173 11151 63229
rect 11237 63173 11293 63229
rect 11379 63173 11435 63229
rect 11521 63173 11577 63229
rect 11663 63173 11719 63229
rect 11805 63173 11861 63229
rect 11947 63173 12003 63229
rect 12089 63173 12145 63229
rect 12231 63173 12287 63229
rect 12373 63173 12429 63229
rect 12515 63173 12571 63229
rect 12657 63173 12713 63229
rect 12799 63173 12855 63229
rect 12941 63173 12997 63229
rect 13083 63173 13139 63229
rect 13225 63173 13281 63229
rect 13367 63173 13423 63229
rect 13509 63173 13565 63229
rect 13651 63173 13707 63229
rect 13793 63173 13849 63229
rect 13935 63173 13991 63229
rect 14077 63173 14133 63229
rect 14219 63173 14275 63229
rect 14361 63173 14417 63229
rect 14503 63173 14559 63229
rect 14645 63173 14701 63229
rect 14787 63173 14843 63229
rect 161 63031 217 63087
rect 303 63031 359 63087
rect 445 63031 501 63087
rect 587 63031 643 63087
rect 729 63031 785 63087
rect 871 63031 927 63087
rect 1013 63031 1069 63087
rect 1155 63031 1211 63087
rect 1297 63031 1353 63087
rect 1439 63031 1495 63087
rect 1581 63031 1637 63087
rect 1723 63031 1779 63087
rect 1865 63031 1921 63087
rect 2007 63031 2063 63087
rect 2149 63031 2205 63087
rect 2291 63031 2347 63087
rect 2433 63031 2489 63087
rect 2575 63031 2631 63087
rect 2717 63031 2773 63087
rect 2859 63031 2915 63087
rect 3001 63031 3057 63087
rect 3143 63031 3199 63087
rect 3285 63031 3341 63087
rect 3427 63031 3483 63087
rect 3569 63031 3625 63087
rect 3711 63031 3767 63087
rect 3853 63031 3909 63087
rect 3995 63031 4051 63087
rect 4137 63031 4193 63087
rect 4279 63031 4335 63087
rect 4421 63031 4477 63087
rect 4563 63031 4619 63087
rect 4705 63031 4761 63087
rect 4847 63031 4903 63087
rect 4989 63031 5045 63087
rect 5131 63031 5187 63087
rect 5273 63031 5329 63087
rect 5415 63031 5471 63087
rect 5557 63031 5613 63087
rect 5699 63031 5755 63087
rect 5841 63031 5897 63087
rect 5983 63031 6039 63087
rect 6125 63031 6181 63087
rect 6267 63031 6323 63087
rect 6409 63031 6465 63087
rect 6551 63031 6607 63087
rect 6693 63031 6749 63087
rect 6835 63031 6891 63087
rect 6977 63031 7033 63087
rect 7119 63031 7175 63087
rect 7261 63031 7317 63087
rect 7403 63031 7459 63087
rect 7545 63031 7601 63087
rect 7687 63031 7743 63087
rect 7829 63031 7885 63087
rect 7971 63031 8027 63087
rect 8113 63031 8169 63087
rect 8255 63031 8311 63087
rect 8397 63031 8453 63087
rect 8539 63031 8595 63087
rect 8681 63031 8737 63087
rect 8823 63031 8879 63087
rect 8965 63031 9021 63087
rect 9107 63031 9163 63087
rect 9249 63031 9305 63087
rect 9391 63031 9447 63087
rect 9533 63031 9589 63087
rect 9675 63031 9731 63087
rect 9817 63031 9873 63087
rect 9959 63031 10015 63087
rect 10101 63031 10157 63087
rect 10243 63031 10299 63087
rect 10385 63031 10441 63087
rect 10527 63031 10583 63087
rect 10669 63031 10725 63087
rect 10811 63031 10867 63087
rect 10953 63031 11009 63087
rect 11095 63031 11151 63087
rect 11237 63031 11293 63087
rect 11379 63031 11435 63087
rect 11521 63031 11577 63087
rect 11663 63031 11719 63087
rect 11805 63031 11861 63087
rect 11947 63031 12003 63087
rect 12089 63031 12145 63087
rect 12231 63031 12287 63087
rect 12373 63031 12429 63087
rect 12515 63031 12571 63087
rect 12657 63031 12713 63087
rect 12799 63031 12855 63087
rect 12941 63031 12997 63087
rect 13083 63031 13139 63087
rect 13225 63031 13281 63087
rect 13367 63031 13423 63087
rect 13509 63031 13565 63087
rect 13651 63031 13707 63087
rect 13793 63031 13849 63087
rect 13935 63031 13991 63087
rect 14077 63031 14133 63087
rect 14219 63031 14275 63087
rect 14361 63031 14417 63087
rect 14503 63031 14559 63087
rect 14645 63031 14701 63087
rect 14787 63031 14843 63087
rect 161 62889 217 62945
rect 303 62889 359 62945
rect 445 62889 501 62945
rect 587 62889 643 62945
rect 729 62889 785 62945
rect 871 62889 927 62945
rect 1013 62889 1069 62945
rect 1155 62889 1211 62945
rect 1297 62889 1353 62945
rect 1439 62889 1495 62945
rect 1581 62889 1637 62945
rect 1723 62889 1779 62945
rect 1865 62889 1921 62945
rect 2007 62889 2063 62945
rect 2149 62889 2205 62945
rect 2291 62889 2347 62945
rect 2433 62889 2489 62945
rect 2575 62889 2631 62945
rect 2717 62889 2773 62945
rect 2859 62889 2915 62945
rect 3001 62889 3057 62945
rect 3143 62889 3199 62945
rect 3285 62889 3341 62945
rect 3427 62889 3483 62945
rect 3569 62889 3625 62945
rect 3711 62889 3767 62945
rect 3853 62889 3909 62945
rect 3995 62889 4051 62945
rect 4137 62889 4193 62945
rect 4279 62889 4335 62945
rect 4421 62889 4477 62945
rect 4563 62889 4619 62945
rect 4705 62889 4761 62945
rect 4847 62889 4903 62945
rect 4989 62889 5045 62945
rect 5131 62889 5187 62945
rect 5273 62889 5329 62945
rect 5415 62889 5471 62945
rect 5557 62889 5613 62945
rect 5699 62889 5755 62945
rect 5841 62889 5897 62945
rect 5983 62889 6039 62945
rect 6125 62889 6181 62945
rect 6267 62889 6323 62945
rect 6409 62889 6465 62945
rect 6551 62889 6607 62945
rect 6693 62889 6749 62945
rect 6835 62889 6891 62945
rect 6977 62889 7033 62945
rect 7119 62889 7175 62945
rect 7261 62889 7317 62945
rect 7403 62889 7459 62945
rect 7545 62889 7601 62945
rect 7687 62889 7743 62945
rect 7829 62889 7885 62945
rect 7971 62889 8027 62945
rect 8113 62889 8169 62945
rect 8255 62889 8311 62945
rect 8397 62889 8453 62945
rect 8539 62889 8595 62945
rect 8681 62889 8737 62945
rect 8823 62889 8879 62945
rect 8965 62889 9021 62945
rect 9107 62889 9163 62945
rect 9249 62889 9305 62945
rect 9391 62889 9447 62945
rect 9533 62889 9589 62945
rect 9675 62889 9731 62945
rect 9817 62889 9873 62945
rect 9959 62889 10015 62945
rect 10101 62889 10157 62945
rect 10243 62889 10299 62945
rect 10385 62889 10441 62945
rect 10527 62889 10583 62945
rect 10669 62889 10725 62945
rect 10811 62889 10867 62945
rect 10953 62889 11009 62945
rect 11095 62889 11151 62945
rect 11237 62889 11293 62945
rect 11379 62889 11435 62945
rect 11521 62889 11577 62945
rect 11663 62889 11719 62945
rect 11805 62889 11861 62945
rect 11947 62889 12003 62945
rect 12089 62889 12145 62945
rect 12231 62889 12287 62945
rect 12373 62889 12429 62945
rect 12515 62889 12571 62945
rect 12657 62889 12713 62945
rect 12799 62889 12855 62945
rect 12941 62889 12997 62945
rect 13083 62889 13139 62945
rect 13225 62889 13281 62945
rect 13367 62889 13423 62945
rect 13509 62889 13565 62945
rect 13651 62889 13707 62945
rect 13793 62889 13849 62945
rect 13935 62889 13991 62945
rect 14077 62889 14133 62945
rect 14219 62889 14275 62945
rect 14361 62889 14417 62945
rect 14503 62889 14559 62945
rect 14645 62889 14701 62945
rect 14787 62889 14843 62945
rect 161 62747 217 62803
rect 303 62747 359 62803
rect 445 62747 501 62803
rect 587 62747 643 62803
rect 729 62747 785 62803
rect 871 62747 927 62803
rect 1013 62747 1069 62803
rect 1155 62747 1211 62803
rect 1297 62747 1353 62803
rect 1439 62747 1495 62803
rect 1581 62747 1637 62803
rect 1723 62747 1779 62803
rect 1865 62747 1921 62803
rect 2007 62747 2063 62803
rect 2149 62747 2205 62803
rect 2291 62747 2347 62803
rect 2433 62747 2489 62803
rect 2575 62747 2631 62803
rect 2717 62747 2773 62803
rect 2859 62747 2915 62803
rect 3001 62747 3057 62803
rect 3143 62747 3199 62803
rect 3285 62747 3341 62803
rect 3427 62747 3483 62803
rect 3569 62747 3625 62803
rect 3711 62747 3767 62803
rect 3853 62747 3909 62803
rect 3995 62747 4051 62803
rect 4137 62747 4193 62803
rect 4279 62747 4335 62803
rect 4421 62747 4477 62803
rect 4563 62747 4619 62803
rect 4705 62747 4761 62803
rect 4847 62747 4903 62803
rect 4989 62747 5045 62803
rect 5131 62747 5187 62803
rect 5273 62747 5329 62803
rect 5415 62747 5471 62803
rect 5557 62747 5613 62803
rect 5699 62747 5755 62803
rect 5841 62747 5897 62803
rect 5983 62747 6039 62803
rect 6125 62747 6181 62803
rect 6267 62747 6323 62803
rect 6409 62747 6465 62803
rect 6551 62747 6607 62803
rect 6693 62747 6749 62803
rect 6835 62747 6891 62803
rect 6977 62747 7033 62803
rect 7119 62747 7175 62803
rect 7261 62747 7317 62803
rect 7403 62747 7459 62803
rect 7545 62747 7601 62803
rect 7687 62747 7743 62803
rect 7829 62747 7885 62803
rect 7971 62747 8027 62803
rect 8113 62747 8169 62803
rect 8255 62747 8311 62803
rect 8397 62747 8453 62803
rect 8539 62747 8595 62803
rect 8681 62747 8737 62803
rect 8823 62747 8879 62803
rect 8965 62747 9021 62803
rect 9107 62747 9163 62803
rect 9249 62747 9305 62803
rect 9391 62747 9447 62803
rect 9533 62747 9589 62803
rect 9675 62747 9731 62803
rect 9817 62747 9873 62803
rect 9959 62747 10015 62803
rect 10101 62747 10157 62803
rect 10243 62747 10299 62803
rect 10385 62747 10441 62803
rect 10527 62747 10583 62803
rect 10669 62747 10725 62803
rect 10811 62747 10867 62803
rect 10953 62747 11009 62803
rect 11095 62747 11151 62803
rect 11237 62747 11293 62803
rect 11379 62747 11435 62803
rect 11521 62747 11577 62803
rect 11663 62747 11719 62803
rect 11805 62747 11861 62803
rect 11947 62747 12003 62803
rect 12089 62747 12145 62803
rect 12231 62747 12287 62803
rect 12373 62747 12429 62803
rect 12515 62747 12571 62803
rect 12657 62747 12713 62803
rect 12799 62747 12855 62803
rect 12941 62747 12997 62803
rect 13083 62747 13139 62803
rect 13225 62747 13281 62803
rect 13367 62747 13423 62803
rect 13509 62747 13565 62803
rect 13651 62747 13707 62803
rect 13793 62747 13849 62803
rect 13935 62747 13991 62803
rect 14077 62747 14133 62803
rect 14219 62747 14275 62803
rect 14361 62747 14417 62803
rect 14503 62747 14559 62803
rect 14645 62747 14701 62803
rect 14787 62747 14843 62803
rect 161 62605 217 62661
rect 303 62605 359 62661
rect 445 62605 501 62661
rect 587 62605 643 62661
rect 729 62605 785 62661
rect 871 62605 927 62661
rect 1013 62605 1069 62661
rect 1155 62605 1211 62661
rect 1297 62605 1353 62661
rect 1439 62605 1495 62661
rect 1581 62605 1637 62661
rect 1723 62605 1779 62661
rect 1865 62605 1921 62661
rect 2007 62605 2063 62661
rect 2149 62605 2205 62661
rect 2291 62605 2347 62661
rect 2433 62605 2489 62661
rect 2575 62605 2631 62661
rect 2717 62605 2773 62661
rect 2859 62605 2915 62661
rect 3001 62605 3057 62661
rect 3143 62605 3199 62661
rect 3285 62605 3341 62661
rect 3427 62605 3483 62661
rect 3569 62605 3625 62661
rect 3711 62605 3767 62661
rect 3853 62605 3909 62661
rect 3995 62605 4051 62661
rect 4137 62605 4193 62661
rect 4279 62605 4335 62661
rect 4421 62605 4477 62661
rect 4563 62605 4619 62661
rect 4705 62605 4761 62661
rect 4847 62605 4903 62661
rect 4989 62605 5045 62661
rect 5131 62605 5187 62661
rect 5273 62605 5329 62661
rect 5415 62605 5471 62661
rect 5557 62605 5613 62661
rect 5699 62605 5755 62661
rect 5841 62605 5897 62661
rect 5983 62605 6039 62661
rect 6125 62605 6181 62661
rect 6267 62605 6323 62661
rect 6409 62605 6465 62661
rect 6551 62605 6607 62661
rect 6693 62605 6749 62661
rect 6835 62605 6891 62661
rect 6977 62605 7033 62661
rect 7119 62605 7175 62661
rect 7261 62605 7317 62661
rect 7403 62605 7459 62661
rect 7545 62605 7601 62661
rect 7687 62605 7743 62661
rect 7829 62605 7885 62661
rect 7971 62605 8027 62661
rect 8113 62605 8169 62661
rect 8255 62605 8311 62661
rect 8397 62605 8453 62661
rect 8539 62605 8595 62661
rect 8681 62605 8737 62661
rect 8823 62605 8879 62661
rect 8965 62605 9021 62661
rect 9107 62605 9163 62661
rect 9249 62605 9305 62661
rect 9391 62605 9447 62661
rect 9533 62605 9589 62661
rect 9675 62605 9731 62661
rect 9817 62605 9873 62661
rect 9959 62605 10015 62661
rect 10101 62605 10157 62661
rect 10243 62605 10299 62661
rect 10385 62605 10441 62661
rect 10527 62605 10583 62661
rect 10669 62605 10725 62661
rect 10811 62605 10867 62661
rect 10953 62605 11009 62661
rect 11095 62605 11151 62661
rect 11237 62605 11293 62661
rect 11379 62605 11435 62661
rect 11521 62605 11577 62661
rect 11663 62605 11719 62661
rect 11805 62605 11861 62661
rect 11947 62605 12003 62661
rect 12089 62605 12145 62661
rect 12231 62605 12287 62661
rect 12373 62605 12429 62661
rect 12515 62605 12571 62661
rect 12657 62605 12713 62661
rect 12799 62605 12855 62661
rect 12941 62605 12997 62661
rect 13083 62605 13139 62661
rect 13225 62605 13281 62661
rect 13367 62605 13423 62661
rect 13509 62605 13565 62661
rect 13651 62605 13707 62661
rect 13793 62605 13849 62661
rect 13935 62605 13991 62661
rect 14077 62605 14133 62661
rect 14219 62605 14275 62661
rect 14361 62605 14417 62661
rect 14503 62605 14559 62661
rect 14645 62605 14701 62661
rect 14787 62605 14843 62661
rect 161 62463 217 62519
rect 303 62463 359 62519
rect 445 62463 501 62519
rect 587 62463 643 62519
rect 729 62463 785 62519
rect 871 62463 927 62519
rect 1013 62463 1069 62519
rect 1155 62463 1211 62519
rect 1297 62463 1353 62519
rect 1439 62463 1495 62519
rect 1581 62463 1637 62519
rect 1723 62463 1779 62519
rect 1865 62463 1921 62519
rect 2007 62463 2063 62519
rect 2149 62463 2205 62519
rect 2291 62463 2347 62519
rect 2433 62463 2489 62519
rect 2575 62463 2631 62519
rect 2717 62463 2773 62519
rect 2859 62463 2915 62519
rect 3001 62463 3057 62519
rect 3143 62463 3199 62519
rect 3285 62463 3341 62519
rect 3427 62463 3483 62519
rect 3569 62463 3625 62519
rect 3711 62463 3767 62519
rect 3853 62463 3909 62519
rect 3995 62463 4051 62519
rect 4137 62463 4193 62519
rect 4279 62463 4335 62519
rect 4421 62463 4477 62519
rect 4563 62463 4619 62519
rect 4705 62463 4761 62519
rect 4847 62463 4903 62519
rect 4989 62463 5045 62519
rect 5131 62463 5187 62519
rect 5273 62463 5329 62519
rect 5415 62463 5471 62519
rect 5557 62463 5613 62519
rect 5699 62463 5755 62519
rect 5841 62463 5897 62519
rect 5983 62463 6039 62519
rect 6125 62463 6181 62519
rect 6267 62463 6323 62519
rect 6409 62463 6465 62519
rect 6551 62463 6607 62519
rect 6693 62463 6749 62519
rect 6835 62463 6891 62519
rect 6977 62463 7033 62519
rect 7119 62463 7175 62519
rect 7261 62463 7317 62519
rect 7403 62463 7459 62519
rect 7545 62463 7601 62519
rect 7687 62463 7743 62519
rect 7829 62463 7885 62519
rect 7971 62463 8027 62519
rect 8113 62463 8169 62519
rect 8255 62463 8311 62519
rect 8397 62463 8453 62519
rect 8539 62463 8595 62519
rect 8681 62463 8737 62519
rect 8823 62463 8879 62519
rect 8965 62463 9021 62519
rect 9107 62463 9163 62519
rect 9249 62463 9305 62519
rect 9391 62463 9447 62519
rect 9533 62463 9589 62519
rect 9675 62463 9731 62519
rect 9817 62463 9873 62519
rect 9959 62463 10015 62519
rect 10101 62463 10157 62519
rect 10243 62463 10299 62519
rect 10385 62463 10441 62519
rect 10527 62463 10583 62519
rect 10669 62463 10725 62519
rect 10811 62463 10867 62519
rect 10953 62463 11009 62519
rect 11095 62463 11151 62519
rect 11237 62463 11293 62519
rect 11379 62463 11435 62519
rect 11521 62463 11577 62519
rect 11663 62463 11719 62519
rect 11805 62463 11861 62519
rect 11947 62463 12003 62519
rect 12089 62463 12145 62519
rect 12231 62463 12287 62519
rect 12373 62463 12429 62519
rect 12515 62463 12571 62519
rect 12657 62463 12713 62519
rect 12799 62463 12855 62519
rect 12941 62463 12997 62519
rect 13083 62463 13139 62519
rect 13225 62463 13281 62519
rect 13367 62463 13423 62519
rect 13509 62463 13565 62519
rect 13651 62463 13707 62519
rect 13793 62463 13849 62519
rect 13935 62463 13991 62519
rect 14077 62463 14133 62519
rect 14219 62463 14275 62519
rect 14361 62463 14417 62519
rect 14503 62463 14559 62519
rect 14645 62463 14701 62519
rect 14787 62463 14843 62519
rect 161 62321 217 62377
rect 303 62321 359 62377
rect 445 62321 501 62377
rect 587 62321 643 62377
rect 729 62321 785 62377
rect 871 62321 927 62377
rect 1013 62321 1069 62377
rect 1155 62321 1211 62377
rect 1297 62321 1353 62377
rect 1439 62321 1495 62377
rect 1581 62321 1637 62377
rect 1723 62321 1779 62377
rect 1865 62321 1921 62377
rect 2007 62321 2063 62377
rect 2149 62321 2205 62377
rect 2291 62321 2347 62377
rect 2433 62321 2489 62377
rect 2575 62321 2631 62377
rect 2717 62321 2773 62377
rect 2859 62321 2915 62377
rect 3001 62321 3057 62377
rect 3143 62321 3199 62377
rect 3285 62321 3341 62377
rect 3427 62321 3483 62377
rect 3569 62321 3625 62377
rect 3711 62321 3767 62377
rect 3853 62321 3909 62377
rect 3995 62321 4051 62377
rect 4137 62321 4193 62377
rect 4279 62321 4335 62377
rect 4421 62321 4477 62377
rect 4563 62321 4619 62377
rect 4705 62321 4761 62377
rect 4847 62321 4903 62377
rect 4989 62321 5045 62377
rect 5131 62321 5187 62377
rect 5273 62321 5329 62377
rect 5415 62321 5471 62377
rect 5557 62321 5613 62377
rect 5699 62321 5755 62377
rect 5841 62321 5897 62377
rect 5983 62321 6039 62377
rect 6125 62321 6181 62377
rect 6267 62321 6323 62377
rect 6409 62321 6465 62377
rect 6551 62321 6607 62377
rect 6693 62321 6749 62377
rect 6835 62321 6891 62377
rect 6977 62321 7033 62377
rect 7119 62321 7175 62377
rect 7261 62321 7317 62377
rect 7403 62321 7459 62377
rect 7545 62321 7601 62377
rect 7687 62321 7743 62377
rect 7829 62321 7885 62377
rect 7971 62321 8027 62377
rect 8113 62321 8169 62377
rect 8255 62321 8311 62377
rect 8397 62321 8453 62377
rect 8539 62321 8595 62377
rect 8681 62321 8737 62377
rect 8823 62321 8879 62377
rect 8965 62321 9021 62377
rect 9107 62321 9163 62377
rect 9249 62321 9305 62377
rect 9391 62321 9447 62377
rect 9533 62321 9589 62377
rect 9675 62321 9731 62377
rect 9817 62321 9873 62377
rect 9959 62321 10015 62377
rect 10101 62321 10157 62377
rect 10243 62321 10299 62377
rect 10385 62321 10441 62377
rect 10527 62321 10583 62377
rect 10669 62321 10725 62377
rect 10811 62321 10867 62377
rect 10953 62321 11009 62377
rect 11095 62321 11151 62377
rect 11237 62321 11293 62377
rect 11379 62321 11435 62377
rect 11521 62321 11577 62377
rect 11663 62321 11719 62377
rect 11805 62321 11861 62377
rect 11947 62321 12003 62377
rect 12089 62321 12145 62377
rect 12231 62321 12287 62377
rect 12373 62321 12429 62377
rect 12515 62321 12571 62377
rect 12657 62321 12713 62377
rect 12799 62321 12855 62377
rect 12941 62321 12997 62377
rect 13083 62321 13139 62377
rect 13225 62321 13281 62377
rect 13367 62321 13423 62377
rect 13509 62321 13565 62377
rect 13651 62321 13707 62377
rect 13793 62321 13849 62377
rect 13935 62321 13991 62377
rect 14077 62321 14133 62377
rect 14219 62321 14275 62377
rect 14361 62321 14417 62377
rect 14503 62321 14559 62377
rect 14645 62321 14701 62377
rect 14787 62321 14843 62377
rect 161 62179 217 62235
rect 303 62179 359 62235
rect 445 62179 501 62235
rect 587 62179 643 62235
rect 729 62179 785 62235
rect 871 62179 927 62235
rect 1013 62179 1069 62235
rect 1155 62179 1211 62235
rect 1297 62179 1353 62235
rect 1439 62179 1495 62235
rect 1581 62179 1637 62235
rect 1723 62179 1779 62235
rect 1865 62179 1921 62235
rect 2007 62179 2063 62235
rect 2149 62179 2205 62235
rect 2291 62179 2347 62235
rect 2433 62179 2489 62235
rect 2575 62179 2631 62235
rect 2717 62179 2773 62235
rect 2859 62179 2915 62235
rect 3001 62179 3057 62235
rect 3143 62179 3199 62235
rect 3285 62179 3341 62235
rect 3427 62179 3483 62235
rect 3569 62179 3625 62235
rect 3711 62179 3767 62235
rect 3853 62179 3909 62235
rect 3995 62179 4051 62235
rect 4137 62179 4193 62235
rect 4279 62179 4335 62235
rect 4421 62179 4477 62235
rect 4563 62179 4619 62235
rect 4705 62179 4761 62235
rect 4847 62179 4903 62235
rect 4989 62179 5045 62235
rect 5131 62179 5187 62235
rect 5273 62179 5329 62235
rect 5415 62179 5471 62235
rect 5557 62179 5613 62235
rect 5699 62179 5755 62235
rect 5841 62179 5897 62235
rect 5983 62179 6039 62235
rect 6125 62179 6181 62235
rect 6267 62179 6323 62235
rect 6409 62179 6465 62235
rect 6551 62179 6607 62235
rect 6693 62179 6749 62235
rect 6835 62179 6891 62235
rect 6977 62179 7033 62235
rect 7119 62179 7175 62235
rect 7261 62179 7317 62235
rect 7403 62179 7459 62235
rect 7545 62179 7601 62235
rect 7687 62179 7743 62235
rect 7829 62179 7885 62235
rect 7971 62179 8027 62235
rect 8113 62179 8169 62235
rect 8255 62179 8311 62235
rect 8397 62179 8453 62235
rect 8539 62179 8595 62235
rect 8681 62179 8737 62235
rect 8823 62179 8879 62235
rect 8965 62179 9021 62235
rect 9107 62179 9163 62235
rect 9249 62179 9305 62235
rect 9391 62179 9447 62235
rect 9533 62179 9589 62235
rect 9675 62179 9731 62235
rect 9817 62179 9873 62235
rect 9959 62179 10015 62235
rect 10101 62179 10157 62235
rect 10243 62179 10299 62235
rect 10385 62179 10441 62235
rect 10527 62179 10583 62235
rect 10669 62179 10725 62235
rect 10811 62179 10867 62235
rect 10953 62179 11009 62235
rect 11095 62179 11151 62235
rect 11237 62179 11293 62235
rect 11379 62179 11435 62235
rect 11521 62179 11577 62235
rect 11663 62179 11719 62235
rect 11805 62179 11861 62235
rect 11947 62179 12003 62235
rect 12089 62179 12145 62235
rect 12231 62179 12287 62235
rect 12373 62179 12429 62235
rect 12515 62179 12571 62235
rect 12657 62179 12713 62235
rect 12799 62179 12855 62235
rect 12941 62179 12997 62235
rect 13083 62179 13139 62235
rect 13225 62179 13281 62235
rect 13367 62179 13423 62235
rect 13509 62179 13565 62235
rect 13651 62179 13707 62235
rect 13793 62179 13849 62235
rect 13935 62179 13991 62235
rect 14077 62179 14133 62235
rect 14219 62179 14275 62235
rect 14361 62179 14417 62235
rect 14503 62179 14559 62235
rect 14645 62179 14701 62235
rect 14787 62179 14843 62235
rect 161 62037 217 62093
rect 303 62037 359 62093
rect 445 62037 501 62093
rect 587 62037 643 62093
rect 729 62037 785 62093
rect 871 62037 927 62093
rect 1013 62037 1069 62093
rect 1155 62037 1211 62093
rect 1297 62037 1353 62093
rect 1439 62037 1495 62093
rect 1581 62037 1637 62093
rect 1723 62037 1779 62093
rect 1865 62037 1921 62093
rect 2007 62037 2063 62093
rect 2149 62037 2205 62093
rect 2291 62037 2347 62093
rect 2433 62037 2489 62093
rect 2575 62037 2631 62093
rect 2717 62037 2773 62093
rect 2859 62037 2915 62093
rect 3001 62037 3057 62093
rect 3143 62037 3199 62093
rect 3285 62037 3341 62093
rect 3427 62037 3483 62093
rect 3569 62037 3625 62093
rect 3711 62037 3767 62093
rect 3853 62037 3909 62093
rect 3995 62037 4051 62093
rect 4137 62037 4193 62093
rect 4279 62037 4335 62093
rect 4421 62037 4477 62093
rect 4563 62037 4619 62093
rect 4705 62037 4761 62093
rect 4847 62037 4903 62093
rect 4989 62037 5045 62093
rect 5131 62037 5187 62093
rect 5273 62037 5329 62093
rect 5415 62037 5471 62093
rect 5557 62037 5613 62093
rect 5699 62037 5755 62093
rect 5841 62037 5897 62093
rect 5983 62037 6039 62093
rect 6125 62037 6181 62093
rect 6267 62037 6323 62093
rect 6409 62037 6465 62093
rect 6551 62037 6607 62093
rect 6693 62037 6749 62093
rect 6835 62037 6891 62093
rect 6977 62037 7033 62093
rect 7119 62037 7175 62093
rect 7261 62037 7317 62093
rect 7403 62037 7459 62093
rect 7545 62037 7601 62093
rect 7687 62037 7743 62093
rect 7829 62037 7885 62093
rect 7971 62037 8027 62093
rect 8113 62037 8169 62093
rect 8255 62037 8311 62093
rect 8397 62037 8453 62093
rect 8539 62037 8595 62093
rect 8681 62037 8737 62093
rect 8823 62037 8879 62093
rect 8965 62037 9021 62093
rect 9107 62037 9163 62093
rect 9249 62037 9305 62093
rect 9391 62037 9447 62093
rect 9533 62037 9589 62093
rect 9675 62037 9731 62093
rect 9817 62037 9873 62093
rect 9959 62037 10015 62093
rect 10101 62037 10157 62093
rect 10243 62037 10299 62093
rect 10385 62037 10441 62093
rect 10527 62037 10583 62093
rect 10669 62037 10725 62093
rect 10811 62037 10867 62093
rect 10953 62037 11009 62093
rect 11095 62037 11151 62093
rect 11237 62037 11293 62093
rect 11379 62037 11435 62093
rect 11521 62037 11577 62093
rect 11663 62037 11719 62093
rect 11805 62037 11861 62093
rect 11947 62037 12003 62093
rect 12089 62037 12145 62093
rect 12231 62037 12287 62093
rect 12373 62037 12429 62093
rect 12515 62037 12571 62093
rect 12657 62037 12713 62093
rect 12799 62037 12855 62093
rect 12941 62037 12997 62093
rect 13083 62037 13139 62093
rect 13225 62037 13281 62093
rect 13367 62037 13423 62093
rect 13509 62037 13565 62093
rect 13651 62037 13707 62093
rect 13793 62037 13849 62093
rect 13935 62037 13991 62093
rect 14077 62037 14133 62093
rect 14219 62037 14275 62093
rect 14361 62037 14417 62093
rect 14503 62037 14559 62093
rect 14645 62037 14701 62093
rect 14787 62037 14843 62093
rect 161 61707 217 61763
rect 303 61707 359 61763
rect 445 61707 501 61763
rect 587 61707 643 61763
rect 729 61707 785 61763
rect 871 61707 927 61763
rect 1013 61707 1069 61763
rect 1155 61707 1211 61763
rect 1297 61707 1353 61763
rect 1439 61707 1495 61763
rect 1581 61707 1637 61763
rect 1723 61707 1779 61763
rect 1865 61707 1921 61763
rect 2007 61707 2063 61763
rect 2149 61707 2205 61763
rect 2291 61707 2347 61763
rect 2433 61707 2489 61763
rect 2575 61707 2631 61763
rect 2717 61707 2773 61763
rect 2859 61707 2915 61763
rect 3001 61707 3057 61763
rect 3143 61707 3199 61763
rect 3285 61707 3341 61763
rect 3427 61707 3483 61763
rect 3569 61707 3625 61763
rect 3711 61707 3767 61763
rect 3853 61707 3909 61763
rect 3995 61707 4051 61763
rect 4137 61707 4193 61763
rect 4279 61707 4335 61763
rect 4421 61707 4477 61763
rect 4563 61707 4619 61763
rect 4705 61707 4761 61763
rect 4847 61707 4903 61763
rect 4989 61707 5045 61763
rect 5131 61707 5187 61763
rect 5273 61707 5329 61763
rect 5415 61707 5471 61763
rect 5557 61707 5613 61763
rect 5699 61707 5755 61763
rect 5841 61707 5897 61763
rect 5983 61707 6039 61763
rect 6125 61707 6181 61763
rect 6267 61707 6323 61763
rect 6409 61707 6465 61763
rect 6551 61707 6607 61763
rect 6693 61707 6749 61763
rect 6835 61707 6891 61763
rect 6977 61707 7033 61763
rect 7119 61707 7175 61763
rect 7261 61707 7317 61763
rect 7403 61707 7459 61763
rect 7545 61707 7601 61763
rect 7687 61707 7743 61763
rect 7829 61707 7885 61763
rect 7971 61707 8027 61763
rect 8113 61707 8169 61763
rect 8255 61707 8311 61763
rect 8397 61707 8453 61763
rect 8539 61707 8595 61763
rect 8681 61707 8737 61763
rect 8823 61707 8879 61763
rect 8965 61707 9021 61763
rect 9107 61707 9163 61763
rect 9249 61707 9305 61763
rect 9391 61707 9447 61763
rect 9533 61707 9589 61763
rect 9675 61707 9731 61763
rect 9817 61707 9873 61763
rect 9959 61707 10015 61763
rect 10101 61707 10157 61763
rect 10243 61707 10299 61763
rect 10385 61707 10441 61763
rect 10527 61707 10583 61763
rect 10669 61707 10725 61763
rect 10811 61707 10867 61763
rect 10953 61707 11009 61763
rect 11095 61707 11151 61763
rect 11237 61707 11293 61763
rect 11379 61707 11435 61763
rect 11521 61707 11577 61763
rect 11663 61707 11719 61763
rect 11805 61707 11861 61763
rect 11947 61707 12003 61763
rect 12089 61707 12145 61763
rect 12231 61707 12287 61763
rect 12373 61707 12429 61763
rect 12515 61707 12571 61763
rect 12657 61707 12713 61763
rect 12799 61707 12855 61763
rect 12941 61707 12997 61763
rect 13083 61707 13139 61763
rect 13225 61707 13281 61763
rect 13367 61707 13423 61763
rect 13509 61707 13565 61763
rect 13651 61707 13707 61763
rect 13793 61707 13849 61763
rect 13935 61707 13991 61763
rect 14077 61707 14133 61763
rect 14219 61707 14275 61763
rect 14361 61707 14417 61763
rect 14503 61707 14559 61763
rect 14645 61707 14701 61763
rect 14787 61707 14843 61763
rect 161 61565 217 61621
rect 303 61565 359 61621
rect 445 61565 501 61621
rect 587 61565 643 61621
rect 729 61565 785 61621
rect 871 61565 927 61621
rect 1013 61565 1069 61621
rect 1155 61565 1211 61621
rect 1297 61565 1353 61621
rect 1439 61565 1495 61621
rect 1581 61565 1637 61621
rect 1723 61565 1779 61621
rect 1865 61565 1921 61621
rect 2007 61565 2063 61621
rect 2149 61565 2205 61621
rect 2291 61565 2347 61621
rect 2433 61565 2489 61621
rect 2575 61565 2631 61621
rect 2717 61565 2773 61621
rect 2859 61565 2915 61621
rect 3001 61565 3057 61621
rect 3143 61565 3199 61621
rect 3285 61565 3341 61621
rect 3427 61565 3483 61621
rect 3569 61565 3625 61621
rect 3711 61565 3767 61621
rect 3853 61565 3909 61621
rect 3995 61565 4051 61621
rect 4137 61565 4193 61621
rect 4279 61565 4335 61621
rect 4421 61565 4477 61621
rect 4563 61565 4619 61621
rect 4705 61565 4761 61621
rect 4847 61565 4903 61621
rect 4989 61565 5045 61621
rect 5131 61565 5187 61621
rect 5273 61565 5329 61621
rect 5415 61565 5471 61621
rect 5557 61565 5613 61621
rect 5699 61565 5755 61621
rect 5841 61565 5897 61621
rect 5983 61565 6039 61621
rect 6125 61565 6181 61621
rect 6267 61565 6323 61621
rect 6409 61565 6465 61621
rect 6551 61565 6607 61621
rect 6693 61565 6749 61621
rect 6835 61565 6891 61621
rect 6977 61565 7033 61621
rect 7119 61565 7175 61621
rect 7261 61565 7317 61621
rect 7403 61565 7459 61621
rect 7545 61565 7601 61621
rect 7687 61565 7743 61621
rect 7829 61565 7885 61621
rect 7971 61565 8027 61621
rect 8113 61565 8169 61621
rect 8255 61565 8311 61621
rect 8397 61565 8453 61621
rect 8539 61565 8595 61621
rect 8681 61565 8737 61621
rect 8823 61565 8879 61621
rect 8965 61565 9021 61621
rect 9107 61565 9163 61621
rect 9249 61565 9305 61621
rect 9391 61565 9447 61621
rect 9533 61565 9589 61621
rect 9675 61565 9731 61621
rect 9817 61565 9873 61621
rect 9959 61565 10015 61621
rect 10101 61565 10157 61621
rect 10243 61565 10299 61621
rect 10385 61565 10441 61621
rect 10527 61565 10583 61621
rect 10669 61565 10725 61621
rect 10811 61565 10867 61621
rect 10953 61565 11009 61621
rect 11095 61565 11151 61621
rect 11237 61565 11293 61621
rect 11379 61565 11435 61621
rect 11521 61565 11577 61621
rect 11663 61565 11719 61621
rect 11805 61565 11861 61621
rect 11947 61565 12003 61621
rect 12089 61565 12145 61621
rect 12231 61565 12287 61621
rect 12373 61565 12429 61621
rect 12515 61565 12571 61621
rect 12657 61565 12713 61621
rect 12799 61565 12855 61621
rect 12941 61565 12997 61621
rect 13083 61565 13139 61621
rect 13225 61565 13281 61621
rect 13367 61565 13423 61621
rect 13509 61565 13565 61621
rect 13651 61565 13707 61621
rect 13793 61565 13849 61621
rect 13935 61565 13991 61621
rect 14077 61565 14133 61621
rect 14219 61565 14275 61621
rect 14361 61565 14417 61621
rect 14503 61565 14559 61621
rect 14645 61565 14701 61621
rect 14787 61565 14843 61621
rect 161 61423 217 61479
rect 303 61423 359 61479
rect 445 61423 501 61479
rect 587 61423 643 61479
rect 729 61423 785 61479
rect 871 61423 927 61479
rect 1013 61423 1069 61479
rect 1155 61423 1211 61479
rect 1297 61423 1353 61479
rect 1439 61423 1495 61479
rect 1581 61423 1637 61479
rect 1723 61423 1779 61479
rect 1865 61423 1921 61479
rect 2007 61423 2063 61479
rect 2149 61423 2205 61479
rect 2291 61423 2347 61479
rect 2433 61423 2489 61479
rect 2575 61423 2631 61479
rect 2717 61423 2773 61479
rect 2859 61423 2915 61479
rect 3001 61423 3057 61479
rect 3143 61423 3199 61479
rect 3285 61423 3341 61479
rect 3427 61423 3483 61479
rect 3569 61423 3625 61479
rect 3711 61423 3767 61479
rect 3853 61423 3909 61479
rect 3995 61423 4051 61479
rect 4137 61423 4193 61479
rect 4279 61423 4335 61479
rect 4421 61423 4477 61479
rect 4563 61423 4619 61479
rect 4705 61423 4761 61479
rect 4847 61423 4903 61479
rect 4989 61423 5045 61479
rect 5131 61423 5187 61479
rect 5273 61423 5329 61479
rect 5415 61423 5471 61479
rect 5557 61423 5613 61479
rect 5699 61423 5755 61479
rect 5841 61423 5897 61479
rect 5983 61423 6039 61479
rect 6125 61423 6181 61479
rect 6267 61423 6323 61479
rect 6409 61423 6465 61479
rect 6551 61423 6607 61479
rect 6693 61423 6749 61479
rect 6835 61423 6891 61479
rect 6977 61423 7033 61479
rect 7119 61423 7175 61479
rect 7261 61423 7317 61479
rect 7403 61423 7459 61479
rect 7545 61423 7601 61479
rect 7687 61423 7743 61479
rect 7829 61423 7885 61479
rect 7971 61423 8027 61479
rect 8113 61423 8169 61479
rect 8255 61423 8311 61479
rect 8397 61423 8453 61479
rect 8539 61423 8595 61479
rect 8681 61423 8737 61479
rect 8823 61423 8879 61479
rect 8965 61423 9021 61479
rect 9107 61423 9163 61479
rect 9249 61423 9305 61479
rect 9391 61423 9447 61479
rect 9533 61423 9589 61479
rect 9675 61423 9731 61479
rect 9817 61423 9873 61479
rect 9959 61423 10015 61479
rect 10101 61423 10157 61479
rect 10243 61423 10299 61479
rect 10385 61423 10441 61479
rect 10527 61423 10583 61479
rect 10669 61423 10725 61479
rect 10811 61423 10867 61479
rect 10953 61423 11009 61479
rect 11095 61423 11151 61479
rect 11237 61423 11293 61479
rect 11379 61423 11435 61479
rect 11521 61423 11577 61479
rect 11663 61423 11719 61479
rect 11805 61423 11861 61479
rect 11947 61423 12003 61479
rect 12089 61423 12145 61479
rect 12231 61423 12287 61479
rect 12373 61423 12429 61479
rect 12515 61423 12571 61479
rect 12657 61423 12713 61479
rect 12799 61423 12855 61479
rect 12941 61423 12997 61479
rect 13083 61423 13139 61479
rect 13225 61423 13281 61479
rect 13367 61423 13423 61479
rect 13509 61423 13565 61479
rect 13651 61423 13707 61479
rect 13793 61423 13849 61479
rect 13935 61423 13991 61479
rect 14077 61423 14133 61479
rect 14219 61423 14275 61479
rect 14361 61423 14417 61479
rect 14503 61423 14559 61479
rect 14645 61423 14701 61479
rect 14787 61423 14843 61479
rect 161 61281 217 61337
rect 303 61281 359 61337
rect 445 61281 501 61337
rect 587 61281 643 61337
rect 729 61281 785 61337
rect 871 61281 927 61337
rect 1013 61281 1069 61337
rect 1155 61281 1211 61337
rect 1297 61281 1353 61337
rect 1439 61281 1495 61337
rect 1581 61281 1637 61337
rect 1723 61281 1779 61337
rect 1865 61281 1921 61337
rect 2007 61281 2063 61337
rect 2149 61281 2205 61337
rect 2291 61281 2347 61337
rect 2433 61281 2489 61337
rect 2575 61281 2631 61337
rect 2717 61281 2773 61337
rect 2859 61281 2915 61337
rect 3001 61281 3057 61337
rect 3143 61281 3199 61337
rect 3285 61281 3341 61337
rect 3427 61281 3483 61337
rect 3569 61281 3625 61337
rect 3711 61281 3767 61337
rect 3853 61281 3909 61337
rect 3995 61281 4051 61337
rect 4137 61281 4193 61337
rect 4279 61281 4335 61337
rect 4421 61281 4477 61337
rect 4563 61281 4619 61337
rect 4705 61281 4761 61337
rect 4847 61281 4903 61337
rect 4989 61281 5045 61337
rect 5131 61281 5187 61337
rect 5273 61281 5329 61337
rect 5415 61281 5471 61337
rect 5557 61281 5613 61337
rect 5699 61281 5755 61337
rect 5841 61281 5897 61337
rect 5983 61281 6039 61337
rect 6125 61281 6181 61337
rect 6267 61281 6323 61337
rect 6409 61281 6465 61337
rect 6551 61281 6607 61337
rect 6693 61281 6749 61337
rect 6835 61281 6891 61337
rect 6977 61281 7033 61337
rect 7119 61281 7175 61337
rect 7261 61281 7317 61337
rect 7403 61281 7459 61337
rect 7545 61281 7601 61337
rect 7687 61281 7743 61337
rect 7829 61281 7885 61337
rect 7971 61281 8027 61337
rect 8113 61281 8169 61337
rect 8255 61281 8311 61337
rect 8397 61281 8453 61337
rect 8539 61281 8595 61337
rect 8681 61281 8737 61337
rect 8823 61281 8879 61337
rect 8965 61281 9021 61337
rect 9107 61281 9163 61337
rect 9249 61281 9305 61337
rect 9391 61281 9447 61337
rect 9533 61281 9589 61337
rect 9675 61281 9731 61337
rect 9817 61281 9873 61337
rect 9959 61281 10015 61337
rect 10101 61281 10157 61337
rect 10243 61281 10299 61337
rect 10385 61281 10441 61337
rect 10527 61281 10583 61337
rect 10669 61281 10725 61337
rect 10811 61281 10867 61337
rect 10953 61281 11009 61337
rect 11095 61281 11151 61337
rect 11237 61281 11293 61337
rect 11379 61281 11435 61337
rect 11521 61281 11577 61337
rect 11663 61281 11719 61337
rect 11805 61281 11861 61337
rect 11947 61281 12003 61337
rect 12089 61281 12145 61337
rect 12231 61281 12287 61337
rect 12373 61281 12429 61337
rect 12515 61281 12571 61337
rect 12657 61281 12713 61337
rect 12799 61281 12855 61337
rect 12941 61281 12997 61337
rect 13083 61281 13139 61337
rect 13225 61281 13281 61337
rect 13367 61281 13423 61337
rect 13509 61281 13565 61337
rect 13651 61281 13707 61337
rect 13793 61281 13849 61337
rect 13935 61281 13991 61337
rect 14077 61281 14133 61337
rect 14219 61281 14275 61337
rect 14361 61281 14417 61337
rect 14503 61281 14559 61337
rect 14645 61281 14701 61337
rect 14787 61281 14843 61337
rect 161 61139 217 61195
rect 303 61139 359 61195
rect 445 61139 501 61195
rect 587 61139 643 61195
rect 729 61139 785 61195
rect 871 61139 927 61195
rect 1013 61139 1069 61195
rect 1155 61139 1211 61195
rect 1297 61139 1353 61195
rect 1439 61139 1495 61195
rect 1581 61139 1637 61195
rect 1723 61139 1779 61195
rect 1865 61139 1921 61195
rect 2007 61139 2063 61195
rect 2149 61139 2205 61195
rect 2291 61139 2347 61195
rect 2433 61139 2489 61195
rect 2575 61139 2631 61195
rect 2717 61139 2773 61195
rect 2859 61139 2915 61195
rect 3001 61139 3057 61195
rect 3143 61139 3199 61195
rect 3285 61139 3341 61195
rect 3427 61139 3483 61195
rect 3569 61139 3625 61195
rect 3711 61139 3767 61195
rect 3853 61139 3909 61195
rect 3995 61139 4051 61195
rect 4137 61139 4193 61195
rect 4279 61139 4335 61195
rect 4421 61139 4477 61195
rect 4563 61139 4619 61195
rect 4705 61139 4761 61195
rect 4847 61139 4903 61195
rect 4989 61139 5045 61195
rect 5131 61139 5187 61195
rect 5273 61139 5329 61195
rect 5415 61139 5471 61195
rect 5557 61139 5613 61195
rect 5699 61139 5755 61195
rect 5841 61139 5897 61195
rect 5983 61139 6039 61195
rect 6125 61139 6181 61195
rect 6267 61139 6323 61195
rect 6409 61139 6465 61195
rect 6551 61139 6607 61195
rect 6693 61139 6749 61195
rect 6835 61139 6891 61195
rect 6977 61139 7033 61195
rect 7119 61139 7175 61195
rect 7261 61139 7317 61195
rect 7403 61139 7459 61195
rect 7545 61139 7601 61195
rect 7687 61139 7743 61195
rect 7829 61139 7885 61195
rect 7971 61139 8027 61195
rect 8113 61139 8169 61195
rect 8255 61139 8311 61195
rect 8397 61139 8453 61195
rect 8539 61139 8595 61195
rect 8681 61139 8737 61195
rect 8823 61139 8879 61195
rect 8965 61139 9021 61195
rect 9107 61139 9163 61195
rect 9249 61139 9305 61195
rect 9391 61139 9447 61195
rect 9533 61139 9589 61195
rect 9675 61139 9731 61195
rect 9817 61139 9873 61195
rect 9959 61139 10015 61195
rect 10101 61139 10157 61195
rect 10243 61139 10299 61195
rect 10385 61139 10441 61195
rect 10527 61139 10583 61195
rect 10669 61139 10725 61195
rect 10811 61139 10867 61195
rect 10953 61139 11009 61195
rect 11095 61139 11151 61195
rect 11237 61139 11293 61195
rect 11379 61139 11435 61195
rect 11521 61139 11577 61195
rect 11663 61139 11719 61195
rect 11805 61139 11861 61195
rect 11947 61139 12003 61195
rect 12089 61139 12145 61195
rect 12231 61139 12287 61195
rect 12373 61139 12429 61195
rect 12515 61139 12571 61195
rect 12657 61139 12713 61195
rect 12799 61139 12855 61195
rect 12941 61139 12997 61195
rect 13083 61139 13139 61195
rect 13225 61139 13281 61195
rect 13367 61139 13423 61195
rect 13509 61139 13565 61195
rect 13651 61139 13707 61195
rect 13793 61139 13849 61195
rect 13935 61139 13991 61195
rect 14077 61139 14133 61195
rect 14219 61139 14275 61195
rect 14361 61139 14417 61195
rect 14503 61139 14559 61195
rect 14645 61139 14701 61195
rect 14787 61139 14843 61195
rect 161 60997 217 61053
rect 303 60997 359 61053
rect 445 60997 501 61053
rect 587 60997 643 61053
rect 729 60997 785 61053
rect 871 60997 927 61053
rect 1013 60997 1069 61053
rect 1155 60997 1211 61053
rect 1297 60997 1353 61053
rect 1439 60997 1495 61053
rect 1581 60997 1637 61053
rect 1723 60997 1779 61053
rect 1865 60997 1921 61053
rect 2007 60997 2063 61053
rect 2149 60997 2205 61053
rect 2291 60997 2347 61053
rect 2433 60997 2489 61053
rect 2575 60997 2631 61053
rect 2717 60997 2773 61053
rect 2859 60997 2915 61053
rect 3001 60997 3057 61053
rect 3143 60997 3199 61053
rect 3285 60997 3341 61053
rect 3427 60997 3483 61053
rect 3569 60997 3625 61053
rect 3711 60997 3767 61053
rect 3853 60997 3909 61053
rect 3995 60997 4051 61053
rect 4137 60997 4193 61053
rect 4279 60997 4335 61053
rect 4421 60997 4477 61053
rect 4563 60997 4619 61053
rect 4705 60997 4761 61053
rect 4847 60997 4903 61053
rect 4989 60997 5045 61053
rect 5131 60997 5187 61053
rect 5273 60997 5329 61053
rect 5415 60997 5471 61053
rect 5557 60997 5613 61053
rect 5699 60997 5755 61053
rect 5841 60997 5897 61053
rect 5983 60997 6039 61053
rect 6125 60997 6181 61053
rect 6267 60997 6323 61053
rect 6409 60997 6465 61053
rect 6551 60997 6607 61053
rect 6693 60997 6749 61053
rect 6835 60997 6891 61053
rect 6977 60997 7033 61053
rect 7119 60997 7175 61053
rect 7261 60997 7317 61053
rect 7403 60997 7459 61053
rect 7545 60997 7601 61053
rect 7687 60997 7743 61053
rect 7829 60997 7885 61053
rect 7971 60997 8027 61053
rect 8113 60997 8169 61053
rect 8255 60997 8311 61053
rect 8397 60997 8453 61053
rect 8539 60997 8595 61053
rect 8681 60997 8737 61053
rect 8823 60997 8879 61053
rect 8965 60997 9021 61053
rect 9107 60997 9163 61053
rect 9249 60997 9305 61053
rect 9391 60997 9447 61053
rect 9533 60997 9589 61053
rect 9675 60997 9731 61053
rect 9817 60997 9873 61053
rect 9959 60997 10015 61053
rect 10101 60997 10157 61053
rect 10243 60997 10299 61053
rect 10385 60997 10441 61053
rect 10527 60997 10583 61053
rect 10669 60997 10725 61053
rect 10811 60997 10867 61053
rect 10953 60997 11009 61053
rect 11095 60997 11151 61053
rect 11237 60997 11293 61053
rect 11379 60997 11435 61053
rect 11521 60997 11577 61053
rect 11663 60997 11719 61053
rect 11805 60997 11861 61053
rect 11947 60997 12003 61053
rect 12089 60997 12145 61053
rect 12231 60997 12287 61053
rect 12373 60997 12429 61053
rect 12515 60997 12571 61053
rect 12657 60997 12713 61053
rect 12799 60997 12855 61053
rect 12941 60997 12997 61053
rect 13083 60997 13139 61053
rect 13225 60997 13281 61053
rect 13367 60997 13423 61053
rect 13509 60997 13565 61053
rect 13651 60997 13707 61053
rect 13793 60997 13849 61053
rect 13935 60997 13991 61053
rect 14077 60997 14133 61053
rect 14219 60997 14275 61053
rect 14361 60997 14417 61053
rect 14503 60997 14559 61053
rect 14645 60997 14701 61053
rect 14787 60997 14843 61053
rect 161 60855 217 60911
rect 303 60855 359 60911
rect 445 60855 501 60911
rect 587 60855 643 60911
rect 729 60855 785 60911
rect 871 60855 927 60911
rect 1013 60855 1069 60911
rect 1155 60855 1211 60911
rect 1297 60855 1353 60911
rect 1439 60855 1495 60911
rect 1581 60855 1637 60911
rect 1723 60855 1779 60911
rect 1865 60855 1921 60911
rect 2007 60855 2063 60911
rect 2149 60855 2205 60911
rect 2291 60855 2347 60911
rect 2433 60855 2489 60911
rect 2575 60855 2631 60911
rect 2717 60855 2773 60911
rect 2859 60855 2915 60911
rect 3001 60855 3057 60911
rect 3143 60855 3199 60911
rect 3285 60855 3341 60911
rect 3427 60855 3483 60911
rect 3569 60855 3625 60911
rect 3711 60855 3767 60911
rect 3853 60855 3909 60911
rect 3995 60855 4051 60911
rect 4137 60855 4193 60911
rect 4279 60855 4335 60911
rect 4421 60855 4477 60911
rect 4563 60855 4619 60911
rect 4705 60855 4761 60911
rect 4847 60855 4903 60911
rect 4989 60855 5045 60911
rect 5131 60855 5187 60911
rect 5273 60855 5329 60911
rect 5415 60855 5471 60911
rect 5557 60855 5613 60911
rect 5699 60855 5755 60911
rect 5841 60855 5897 60911
rect 5983 60855 6039 60911
rect 6125 60855 6181 60911
rect 6267 60855 6323 60911
rect 6409 60855 6465 60911
rect 6551 60855 6607 60911
rect 6693 60855 6749 60911
rect 6835 60855 6891 60911
rect 6977 60855 7033 60911
rect 7119 60855 7175 60911
rect 7261 60855 7317 60911
rect 7403 60855 7459 60911
rect 7545 60855 7601 60911
rect 7687 60855 7743 60911
rect 7829 60855 7885 60911
rect 7971 60855 8027 60911
rect 8113 60855 8169 60911
rect 8255 60855 8311 60911
rect 8397 60855 8453 60911
rect 8539 60855 8595 60911
rect 8681 60855 8737 60911
rect 8823 60855 8879 60911
rect 8965 60855 9021 60911
rect 9107 60855 9163 60911
rect 9249 60855 9305 60911
rect 9391 60855 9447 60911
rect 9533 60855 9589 60911
rect 9675 60855 9731 60911
rect 9817 60855 9873 60911
rect 9959 60855 10015 60911
rect 10101 60855 10157 60911
rect 10243 60855 10299 60911
rect 10385 60855 10441 60911
rect 10527 60855 10583 60911
rect 10669 60855 10725 60911
rect 10811 60855 10867 60911
rect 10953 60855 11009 60911
rect 11095 60855 11151 60911
rect 11237 60855 11293 60911
rect 11379 60855 11435 60911
rect 11521 60855 11577 60911
rect 11663 60855 11719 60911
rect 11805 60855 11861 60911
rect 11947 60855 12003 60911
rect 12089 60855 12145 60911
rect 12231 60855 12287 60911
rect 12373 60855 12429 60911
rect 12515 60855 12571 60911
rect 12657 60855 12713 60911
rect 12799 60855 12855 60911
rect 12941 60855 12997 60911
rect 13083 60855 13139 60911
rect 13225 60855 13281 60911
rect 13367 60855 13423 60911
rect 13509 60855 13565 60911
rect 13651 60855 13707 60911
rect 13793 60855 13849 60911
rect 13935 60855 13991 60911
rect 14077 60855 14133 60911
rect 14219 60855 14275 60911
rect 14361 60855 14417 60911
rect 14503 60855 14559 60911
rect 14645 60855 14701 60911
rect 14787 60855 14843 60911
rect 161 60713 217 60769
rect 303 60713 359 60769
rect 445 60713 501 60769
rect 587 60713 643 60769
rect 729 60713 785 60769
rect 871 60713 927 60769
rect 1013 60713 1069 60769
rect 1155 60713 1211 60769
rect 1297 60713 1353 60769
rect 1439 60713 1495 60769
rect 1581 60713 1637 60769
rect 1723 60713 1779 60769
rect 1865 60713 1921 60769
rect 2007 60713 2063 60769
rect 2149 60713 2205 60769
rect 2291 60713 2347 60769
rect 2433 60713 2489 60769
rect 2575 60713 2631 60769
rect 2717 60713 2773 60769
rect 2859 60713 2915 60769
rect 3001 60713 3057 60769
rect 3143 60713 3199 60769
rect 3285 60713 3341 60769
rect 3427 60713 3483 60769
rect 3569 60713 3625 60769
rect 3711 60713 3767 60769
rect 3853 60713 3909 60769
rect 3995 60713 4051 60769
rect 4137 60713 4193 60769
rect 4279 60713 4335 60769
rect 4421 60713 4477 60769
rect 4563 60713 4619 60769
rect 4705 60713 4761 60769
rect 4847 60713 4903 60769
rect 4989 60713 5045 60769
rect 5131 60713 5187 60769
rect 5273 60713 5329 60769
rect 5415 60713 5471 60769
rect 5557 60713 5613 60769
rect 5699 60713 5755 60769
rect 5841 60713 5897 60769
rect 5983 60713 6039 60769
rect 6125 60713 6181 60769
rect 6267 60713 6323 60769
rect 6409 60713 6465 60769
rect 6551 60713 6607 60769
rect 6693 60713 6749 60769
rect 6835 60713 6891 60769
rect 6977 60713 7033 60769
rect 7119 60713 7175 60769
rect 7261 60713 7317 60769
rect 7403 60713 7459 60769
rect 7545 60713 7601 60769
rect 7687 60713 7743 60769
rect 7829 60713 7885 60769
rect 7971 60713 8027 60769
rect 8113 60713 8169 60769
rect 8255 60713 8311 60769
rect 8397 60713 8453 60769
rect 8539 60713 8595 60769
rect 8681 60713 8737 60769
rect 8823 60713 8879 60769
rect 8965 60713 9021 60769
rect 9107 60713 9163 60769
rect 9249 60713 9305 60769
rect 9391 60713 9447 60769
rect 9533 60713 9589 60769
rect 9675 60713 9731 60769
rect 9817 60713 9873 60769
rect 9959 60713 10015 60769
rect 10101 60713 10157 60769
rect 10243 60713 10299 60769
rect 10385 60713 10441 60769
rect 10527 60713 10583 60769
rect 10669 60713 10725 60769
rect 10811 60713 10867 60769
rect 10953 60713 11009 60769
rect 11095 60713 11151 60769
rect 11237 60713 11293 60769
rect 11379 60713 11435 60769
rect 11521 60713 11577 60769
rect 11663 60713 11719 60769
rect 11805 60713 11861 60769
rect 11947 60713 12003 60769
rect 12089 60713 12145 60769
rect 12231 60713 12287 60769
rect 12373 60713 12429 60769
rect 12515 60713 12571 60769
rect 12657 60713 12713 60769
rect 12799 60713 12855 60769
rect 12941 60713 12997 60769
rect 13083 60713 13139 60769
rect 13225 60713 13281 60769
rect 13367 60713 13423 60769
rect 13509 60713 13565 60769
rect 13651 60713 13707 60769
rect 13793 60713 13849 60769
rect 13935 60713 13991 60769
rect 14077 60713 14133 60769
rect 14219 60713 14275 60769
rect 14361 60713 14417 60769
rect 14503 60713 14559 60769
rect 14645 60713 14701 60769
rect 14787 60713 14843 60769
rect 161 60571 217 60627
rect 303 60571 359 60627
rect 445 60571 501 60627
rect 587 60571 643 60627
rect 729 60571 785 60627
rect 871 60571 927 60627
rect 1013 60571 1069 60627
rect 1155 60571 1211 60627
rect 1297 60571 1353 60627
rect 1439 60571 1495 60627
rect 1581 60571 1637 60627
rect 1723 60571 1779 60627
rect 1865 60571 1921 60627
rect 2007 60571 2063 60627
rect 2149 60571 2205 60627
rect 2291 60571 2347 60627
rect 2433 60571 2489 60627
rect 2575 60571 2631 60627
rect 2717 60571 2773 60627
rect 2859 60571 2915 60627
rect 3001 60571 3057 60627
rect 3143 60571 3199 60627
rect 3285 60571 3341 60627
rect 3427 60571 3483 60627
rect 3569 60571 3625 60627
rect 3711 60571 3767 60627
rect 3853 60571 3909 60627
rect 3995 60571 4051 60627
rect 4137 60571 4193 60627
rect 4279 60571 4335 60627
rect 4421 60571 4477 60627
rect 4563 60571 4619 60627
rect 4705 60571 4761 60627
rect 4847 60571 4903 60627
rect 4989 60571 5045 60627
rect 5131 60571 5187 60627
rect 5273 60571 5329 60627
rect 5415 60571 5471 60627
rect 5557 60571 5613 60627
rect 5699 60571 5755 60627
rect 5841 60571 5897 60627
rect 5983 60571 6039 60627
rect 6125 60571 6181 60627
rect 6267 60571 6323 60627
rect 6409 60571 6465 60627
rect 6551 60571 6607 60627
rect 6693 60571 6749 60627
rect 6835 60571 6891 60627
rect 6977 60571 7033 60627
rect 7119 60571 7175 60627
rect 7261 60571 7317 60627
rect 7403 60571 7459 60627
rect 7545 60571 7601 60627
rect 7687 60571 7743 60627
rect 7829 60571 7885 60627
rect 7971 60571 8027 60627
rect 8113 60571 8169 60627
rect 8255 60571 8311 60627
rect 8397 60571 8453 60627
rect 8539 60571 8595 60627
rect 8681 60571 8737 60627
rect 8823 60571 8879 60627
rect 8965 60571 9021 60627
rect 9107 60571 9163 60627
rect 9249 60571 9305 60627
rect 9391 60571 9447 60627
rect 9533 60571 9589 60627
rect 9675 60571 9731 60627
rect 9817 60571 9873 60627
rect 9959 60571 10015 60627
rect 10101 60571 10157 60627
rect 10243 60571 10299 60627
rect 10385 60571 10441 60627
rect 10527 60571 10583 60627
rect 10669 60571 10725 60627
rect 10811 60571 10867 60627
rect 10953 60571 11009 60627
rect 11095 60571 11151 60627
rect 11237 60571 11293 60627
rect 11379 60571 11435 60627
rect 11521 60571 11577 60627
rect 11663 60571 11719 60627
rect 11805 60571 11861 60627
rect 11947 60571 12003 60627
rect 12089 60571 12145 60627
rect 12231 60571 12287 60627
rect 12373 60571 12429 60627
rect 12515 60571 12571 60627
rect 12657 60571 12713 60627
rect 12799 60571 12855 60627
rect 12941 60571 12997 60627
rect 13083 60571 13139 60627
rect 13225 60571 13281 60627
rect 13367 60571 13423 60627
rect 13509 60571 13565 60627
rect 13651 60571 13707 60627
rect 13793 60571 13849 60627
rect 13935 60571 13991 60627
rect 14077 60571 14133 60627
rect 14219 60571 14275 60627
rect 14361 60571 14417 60627
rect 14503 60571 14559 60627
rect 14645 60571 14701 60627
rect 14787 60571 14843 60627
rect 161 60429 217 60485
rect 303 60429 359 60485
rect 445 60429 501 60485
rect 587 60429 643 60485
rect 729 60429 785 60485
rect 871 60429 927 60485
rect 1013 60429 1069 60485
rect 1155 60429 1211 60485
rect 1297 60429 1353 60485
rect 1439 60429 1495 60485
rect 1581 60429 1637 60485
rect 1723 60429 1779 60485
rect 1865 60429 1921 60485
rect 2007 60429 2063 60485
rect 2149 60429 2205 60485
rect 2291 60429 2347 60485
rect 2433 60429 2489 60485
rect 2575 60429 2631 60485
rect 2717 60429 2773 60485
rect 2859 60429 2915 60485
rect 3001 60429 3057 60485
rect 3143 60429 3199 60485
rect 3285 60429 3341 60485
rect 3427 60429 3483 60485
rect 3569 60429 3625 60485
rect 3711 60429 3767 60485
rect 3853 60429 3909 60485
rect 3995 60429 4051 60485
rect 4137 60429 4193 60485
rect 4279 60429 4335 60485
rect 4421 60429 4477 60485
rect 4563 60429 4619 60485
rect 4705 60429 4761 60485
rect 4847 60429 4903 60485
rect 4989 60429 5045 60485
rect 5131 60429 5187 60485
rect 5273 60429 5329 60485
rect 5415 60429 5471 60485
rect 5557 60429 5613 60485
rect 5699 60429 5755 60485
rect 5841 60429 5897 60485
rect 5983 60429 6039 60485
rect 6125 60429 6181 60485
rect 6267 60429 6323 60485
rect 6409 60429 6465 60485
rect 6551 60429 6607 60485
rect 6693 60429 6749 60485
rect 6835 60429 6891 60485
rect 6977 60429 7033 60485
rect 7119 60429 7175 60485
rect 7261 60429 7317 60485
rect 7403 60429 7459 60485
rect 7545 60429 7601 60485
rect 7687 60429 7743 60485
rect 7829 60429 7885 60485
rect 7971 60429 8027 60485
rect 8113 60429 8169 60485
rect 8255 60429 8311 60485
rect 8397 60429 8453 60485
rect 8539 60429 8595 60485
rect 8681 60429 8737 60485
rect 8823 60429 8879 60485
rect 8965 60429 9021 60485
rect 9107 60429 9163 60485
rect 9249 60429 9305 60485
rect 9391 60429 9447 60485
rect 9533 60429 9589 60485
rect 9675 60429 9731 60485
rect 9817 60429 9873 60485
rect 9959 60429 10015 60485
rect 10101 60429 10157 60485
rect 10243 60429 10299 60485
rect 10385 60429 10441 60485
rect 10527 60429 10583 60485
rect 10669 60429 10725 60485
rect 10811 60429 10867 60485
rect 10953 60429 11009 60485
rect 11095 60429 11151 60485
rect 11237 60429 11293 60485
rect 11379 60429 11435 60485
rect 11521 60429 11577 60485
rect 11663 60429 11719 60485
rect 11805 60429 11861 60485
rect 11947 60429 12003 60485
rect 12089 60429 12145 60485
rect 12231 60429 12287 60485
rect 12373 60429 12429 60485
rect 12515 60429 12571 60485
rect 12657 60429 12713 60485
rect 12799 60429 12855 60485
rect 12941 60429 12997 60485
rect 13083 60429 13139 60485
rect 13225 60429 13281 60485
rect 13367 60429 13423 60485
rect 13509 60429 13565 60485
rect 13651 60429 13707 60485
rect 13793 60429 13849 60485
rect 13935 60429 13991 60485
rect 14077 60429 14133 60485
rect 14219 60429 14275 60485
rect 14361 60429 14417 60485
rect 14503 60429 14559 60485
rect 14645 60429 14701 60485
rect 14787 60429 14843 60485
rect 161 60115 217 60171
rect 303 60115 359 60171
rect 445 60115 501 60171
rect 587 60115 643 60171
rect 729 60115 785 60171
rect 871 60115 927 60171
rect 1013 60115 1069 60171
rect 1155 60115 1211 60171
rect 1297 60115 1353 60171
rect 1439 60115 1495 60171
rect 1581 60115 1637 60171
rect 1723 60115 1779 60171
rect 1865 60115 1921 60171
rect 2007 60115 2063 60171
rect 2149 60115 2205 60171
rect 2291 60115 2347 60171
rect 2433 60115 2489 60171
rect 2575 60115 2631 60171
rect 2717 60115 2773 60171
rect 2859 60115 2915 60171
rect 3001 60115 3057 60171
rect 3143 60115 3199 60171
rect 3285 60115 3341 60171
rect 3427 60115 3483 60171
rect 3569 60115 3625 60171
rect 3711 60115 3767 60171
rect 3853 60115 3909 60171
rect 3995 60115 4051 60171
rect 4137 60115 4193 60171
rect 4279 60115 4335 60171
rect 4421 60115 4477 60171
rect 4563 60115 4619 60171
rect 4705 60115 4761 60171
rect 4847 60115 4903 60171
rect 4989 60115 5045 60171
rect 5131 60115 5187 60171
rect 5273 60115 5329 60171
rect 5415 60115 5471 60171
rect 5557 60115 5613 60171
rect 5699 60115 5755 60171
rect 5841 60115 5897 60171
rect 5983 60115 6039 60171
rect 6125 60115 6181 60171
rect 6267 60115 6323 60171
rect 6409 60115 6465 60171
rect 6551 60115 6607 60171
rect 6693 60115 6749 60171
rect 6835 60115 6891 60171
rect 6977 60115 7033 60171
rect 7119 60115 7175 60171
rect 7261 60115 7317 60171
rect 7403 60115 7459 60171
rect 7545 60115 7601 60171
rect 7687 60115 7743 60171
rect 7829 60115 7885 60171
rect 7971 60115 8027 60171
rect 8113 60115 8169 60171
rect 8255 60115 8311 60171
rect 8397 60115 8453 60171
rect 8539 60115 8595 60171
rect 8681 60115 8737 60171
rect 8823 60115 8879 60171
rect 8965 60115 9021 60171
rect 9107 60115 9163 60171
rect 9249 60115 9305 60171
rect 9391 60115 9447 60171
rect 9533 60115 9589 60171
rect 9675 60115 9731 60171
rect 9817 60115 9873 60171
rect 9959 60115 10015 60171
rect 10101 60115 10157 60171
rect 10243 60115 10299 60171
rect 10385 60115 10441 60171
rect 10527 60115 10583 60171
rect 10669 60115 10725 60171
rect 10811 60115 10867 60171
rect 10953 60115 11009 60171
rect 11095 60115 11151 60171
rect 11237 60115 11293 60171
rect 11379 60115 11435 60171
rect 11521 60115 11577 60171
rect 11663 60115 11719 60171
rect 11805 60115 11861 60171
rect 11947 60115 12003 60171
rect 12089 60115 12145 60171
rect 12231 60115 12287 60171
rect 12373 60115 12429 60171
rect 12515 60115 12571 60171
rect 12657 60115 12713 60171
rect 12799 60115 12855 60171
rect 12941 60115 12997 60171
rect 13083 60115 13139 60171
rect 13225 60115 13281 60171
rect 13367 60115 13423 60171
rect 13509 60115 13565 60171
rect 13651 60115 13707 60171
rect 13793 60115 13849 60171
rect 13935 60115 13991 60171
rect 14077 60115 14133 60171
rect 14219 60115 14275 60171
rect 14361 60115 14417 60171
rect 14503 60115 14559 60171
rect 14645 60115 14701 60171
rect 14787 60115 14843 60171
rect 161 59973 217 60029
rect 303 59973 359 60029
rect 445 59973 501 60029
rect 587 59973 643 60029
rect 729 59973 785 60029
rect 871 59973 927 60029
rect 1013 59973 1069 60029
rect 1155 59973 1211 60029
rect 1297 59973 1353 60029
rect 1439 59973 1495 60029
rect 1581 59973 1637 60029
rect 1723 59973 1779 60029
rect 1865 59973 1921 60029
rect 2007 59973 2063 60029
rect 2149 59973 2205 60029
rect 2291 59973 2347 60029
rect 2433 59973 2489 60029
rect 2575 59973 2631 60029
rect 2717 59973 2773 60029
rect 2859 59973 2915 60029
rect 3001 59973 3057 60029
rect 3143 59973 3199 60029
rect 3285 59973 3341 60029
rect 3427 59973 3483 60029
rect 3569 59973 3625 60029
rect 3711 59973 3767 60029
rect 3853 59973 3909 60029
rect 3995 59973 4051 60029
rect 4137 59973 4193 60029
rect 4279 59973 4335 60029
rect 4421 59973 4477 60029
rect 4563 59973 4619 60029
rect 4705 59973 4761 60029
rect 4847 59973 4903 60029
rect 4989 59973 5045 60029
rect 5131 59973 5187 60029
rect 5273 59973 5329 60029
rect 5415 59973 5471 60029
rect 5557 59973 5613 60029
rect 5699 59973 5755 60029
rect 5841 59973 5897 60029
rect 5983 59973 6039 60029
rect 6125 59973 6181 60029
rect 6267 59973 6323 60029
rect 6409 59973 6465 60029
rect 6551 59973 6607 60029
rect 6693 59973 6749 60029
rect 6835 59973 6891 60029
rect 6977 59973 7033 60029
rect 7119 59973 7175 60029
rect 7261 59973 7317 60029
rect 7403 59973 7459 60029
rect 7545 59973 7601 60029
rect 7687 59973 7743 60029
rect 7829 59973 7885 60029
rect 7971 59973 8027 60029
rect 8113 59973 8169 60029
rect 8255 59973 8311 60029
rect 8397 59973 8453 60029
rect 8539 59973 8595 60029
rect 8681 59973 8737 60029
rect 8823 59973 8879 60029
rect 8965 59973 9021 60029
rect 9107 59973 9163 60029
rect 9249 59973 9305 60029
rect 9391 59973 9447 60029
rect 9533 59973 9589 60029
rect 9675 59973 9731 60029
rect 9817 59973 9873 60029
rect 9959 59973 10015 60029
rect 10101 59973 10157 60029
rect 10243 59973 10299 60029
rect 10385 59973 10441 60029
rect 10527 59973 10583 60029
rect 10669 59973 10725 60029
rect 10811 59973 10867 60029
rect 10953 59973 11009 60029
rect 11095 59973 11151 60029
rect 11237 59973 11293 60029
rect 11379 59973 11435 60029
rect 11521 59973 11577 60029
rect 11663 59973 11719 60029
rect 11805 59973 11861 60029
rect 11947 59973 12003 60029
rect 12089 59973 12145 60029
rect 12231 59973 12287 60029
rect 12373 59973 12429 60029
rect 12515 59973 12571 60029
rect 12657 59973 12713 60029
rect 12799 59973 12855 60029
rect 12941 59973 12997 60029
rect 13083 59973 13139 60029
rect 13225 59973 13281 60029
rect 13367 59973 13423 60029
rect 13509 59973 13565 60029
rect 13651 59973 13707 60029
rect 13793 59973 13849 60029
rect 13935 59973 13991 60029
rect 14077 59973 14133 60029
rect 14219 59973 14275 60029
rect 14361 59973 14417 60029
rect 14503 59973 14559 60029
rect 14645 59973 14701 60029
rect 14787 59973 14843 60029
rect 161 59831 217 59887
rect 303 59831 359 59887
rect 445 59831 501 59887
rect 587 59831 643 59887
rect 729 59831 785 59887
rect 871 59831 927 59887
rect 1013 59831 1069 59887
rect 1155 59831 1211 59887
rect 1297 59831 1353 59887
rect 1439 59831 1495 59887
rect 1581 59831 1637 59887
rect 1723 59831 1779 59887
rect 1865 59831 1921 59887
rect 2007 59831 2063 59887
rect 2149 59831 2205 59887
rect 2291 59831 2347 59887
rect 2433 59831 2489 59887
rect 2575 59831 2631 59887
rect 2717 59831 2773 59887
rect 2859 59831 2915 59887
rect 3001 59831 3057 59887
rect 3143 59831 3199 59887
rect 3285 59831 3341 59887
rect 3427 59831 3483 59887
rect 3569 59831 3625 59887
rect 3711 59831 3767 59887
rect 3853 59831 3909 59887
rect 3995 59831 4051 59887
rect 4137 59831 4193 59887
rect 4279 59831 4335 59887
rect 4421 59831 4477 59887
rect 4563 59831 4619 59887
rect 4705 59831 4761 59887
rect 4847 59831 4903 59887
rect 4989 59831 5045 59887
rect 5131 59831 5187 59887
rect 5273 59831 5329 59887
rect 5415 59831 5471 59887
rect 5557 59831 5613 59887
rect 5699 59831 5755 59887
rect 5841 59831 5897 59887
rect 5983 59831 6039 59887
rect 6125 59831 6181 59887
rect 6267 59831 6323 59887
rect 6409 59831 6465 59887
rect 6551 59831 6607 59887
rect 6693 59831 6749 59887
rect 6835 59831 6891 59887
rect 6977 59831 7033 59887
rect 7119 59831 7175 59887
rect 7261 59831 7317 59887
rect 7403 59831 7459 59887
rect 7545 59831 7601 59887
rect 7687 59831 7743 59887
rect 7829 59831 7885 59887
rect 7971 59831 8027 59887
rect 8113 59831 8169 59887
rect 8255 59831 8311 59887
rect 8397 59831 8453 59887
rect 8539 59831 8595 59887
rect 8681 59831 8737 59887
rect 8823 59831 8879 59887
rect 8965 59831 9021 59887
rect 9107 59831 9163 59887
rect 9249 59831 9305 59887
rect 9391 59831 9447 59887
rect 9533 59831 9589 59887
rect 9675 59831 9731 59887
rect 9817 59831 9873 59887
rect 9959 59831 10015 59887
rect 10101 59831 10157 59887
rect 10243 59831 10299 59887
rect 10385 59831 10441 59887
rect 10527 59831 10583 59887
rect 10669 59831 10725 59887
rect 10811 59831 10867 59887
rect 10953 59831 11009 59887
rect 11095 59831 11151 59887
rect 11237 59831 11293 59887
rect 11379 59831 11435 59887
rect 11521 59831 11577 59887
rect 11663 59831 11719 59887
rect 11805 59831 11861 59887
rect 11947 59831 12003 59887
rect 12089 59831 12145 59887
rect 12231 59831 12287 59887
rect 12373 59831 12429 59887
rect 12515 59831 12571 59887
rect 12657 59831 12713 59887
rect 12799 59831 12855 59887
rect 12941 59831 12997 59887
rect 13083 59831 13139 59887
rect 13225 59831 13281 59887
rect 13367 59831 13423 59887
rect 13509 59831 13565 59887
rect 13651 59831 13707 59887
rect 13793 59831 13849 59887
rect 13935 59831 13991 59887
rect 14077 59831 14133 59887
rect 14219 59831 14275 59887
rect 14361 59831 14417 59887
rect 14503 59831 14559 59887
rect 14645 59831 14701 59887
rect 14787 59831 14843 59887
rect 161 59689 217 59745
rect 303 59689 359 59745
rect 445 59689 501 59745
rect 587 59689 643 59745
rect 729 59689 785 59745
rect 871 59689 927 59745
rect 1013 59689 1069 59745
rect 1155 59689 1211 59745
rect 1297 59689 1353 59745
rect 1439 59689 1495 59745
rect 1581 59689 1637 59745
rect 1723 59689 1779 59745
rect 1865 59689 1921 59745
rect 2007 59689 2063 59745
rect 2149 59689 2205 59745
rect 2291 59689 2347 59745
rect 2433 59689 2489 59745
rect 2575 59689 2631 59745
rect 2717 59689 2773 59745
rect 2859 59689 2915 59745
rect 3001 59689 3057 59745
rect 3143 59689 3199 59745
rect 3285 59689 3341 59745
rect 3427 59689 3483 59745
rect 3569 59689 3625 59745
rect 3711 59689 3767 59745
rect 3853 59689 3909 59745
rect 3995 59689 4051 59745
rect 4137 59689 4193 59745
rect 4279 59689 4335 59745
rect 4421 59689 4477 59745
rect 4563 59689 4619 59745
rect 4705 59689 4761 59745
rect 4847 59689 4903 59745
rect 4989 59689 5045 59745
rect 5131 59689 5187 59745
rect 5273 59689 5329 59745
rect 5415 59689 5471 59745
rect 5557 59689 5613 59745
rect 5699 59689 5755 59745
rect 5841 59689 5897 59745
rect 5983 59689 6039 59745
rect 6125 59689 6181 59745
rect 6267 59689 6323 59745
rect 6409 59689 6465 59745
rect 6551 59689 6607 59745
rect 6693 59689 6749 59745
rect 6835 59689 6891 59745
rect 6977 59689 7033 59745
rect 7119 59689 7175 59745
rect 7261 59689 7317 59745
rect 7403 59689 7459 59745
rect 7545 59689 7601 59745
rect 7687 59689 7743 59745
rect 7829 59689 7885 59745
rect 7971 59689 8027 59745
rect 8113 59689 8169 59745
rect 8255 59689 8311 59745
rect 8397 59689 8453 59745
rect 8539 59689 8595 59745
rect 8681 59689 8737 59745
rect 8823 59689 8879 59745
rect 8965 59689 9021 59745
rect 9107 59689 9163 59745
rect 9249 59689 9305 59745
rect 9391 59689 9447 59745
rect 9533 59689 9589 59745
rect 9675 59689 9731 59745
rect 9817 59689 9873 59745
rect 9959 59689 10015 59745
rect 10101 59689 10157 59745
rect 10243 59689 10299 59745
rect 10385 59689 10441 59745
rect 10527 59689 10583 59745
rect 10669 59689 10725 59745
rect 10811 59689 10867 59745
rect 10953 59689 11009 59745
rect 11095 59689 11151 59745
rect 11237 59689 11293 59745
rect 11379 59689 11435 59745
rect 11521 59689 11577 59745
rect 11663 59689 11719 59745
rect 11805 59689 11861 59745
rect 11947 59689 12003 59745
rect 12089 59689 12145 59745
rect 12231 59689 12287 59745
rect 12373 59689 12429 59745
rect 12515 59689 12571 59745
rect 12657 59689 12713 59745
rect 12799 59689 12855 59745
rect 12941 59689 12997 59745
rect 13083 59689 13139 59745
rect 13225 59689 13281 59745
rect 13367 59689 13423 59745
rect 13509 59689 13565 59745
rect 13651 59689 13707 59745
rect 13793 59689 13849 59745
rect 13935 59689 13991 59745
rect 14077 59689 14133 59745
rect 14219 59689 14275 59745
rect 14361 59689 14417 59745
rect 14503 59689 14559 59745
rect 14645 59689 14701 59745
rect 14787 59689 14843 59745
rect 161 59547 217 59603
rect 303 59547 359 59603
rect 445 59547 501 59603
rect 587 59547 643 59603
rect 729 59547 785 59603
rect 871 59547 927 59603
rect 1013 59547 1069 59603
rect 1155 59547 1211 59603
rect 1297 59547 1353 59603
rect 1439 59547 1495 59603
rect 1581 59547 1637 59603
rect 1723 59547 1779 59603
rect 1865 59547 1921 59603
rect 2007 59547 2063 59603
rect 2149 59547 2205 59603
rect 2291 59547 2347 59603
rect 2433 59547 2489 59603
rect 2575 59547 2631 59603
rect 2717 59547 2773 59603
rect 2859 59547 2915 59603
rect 3001 59547 3057 59603
rect 3143 59547 3199 59603
rect 3285 59547 3341 59603
rect 3427 59547 3483 59603
rect 3569 59547 3625 59603
rect 3711 59547 3767 59603
rect 3853 59547 3909 59603
rect 3995 59547 4051 59603
rect 4137 59547 4193 59603
rect 4279 59547 4335 59603
rect 4421 59547 4477 59603
rect 4563 59547 4619 59603
rect 4705 59547 4761 59603
rect 4847 59547 4903 59603
rect 4989 59547 5045 59603
rect 5131 59547 5187 59603
rect 5273 59547 5329 59603
rect 5415 59547 5471 59603
rect 5557 59547 5613 59603
rect 5699 59547 5755 59603
rect 5841 59547 5897 59603
rect 5983 59547 6039 59603
rect 6125 59547 6181 59603
rect 6267 59547 6323 59603
rect 6409 59547 6465 59603
rect 6551 59547 6607 59603
rect 6693 59547 6749 59603
rect 6835 59547 6891 59603
rect 6977 59547 7033 59603
rect 7119 59547 7175 59603
rect 7261 59547 7317 59603
rect 7403 59547 7459 59603
rect 7545 59547 7601 59603
rect 7687 59547 7743 59603
rect 7829 59547 7885 59603
rect 7971 59547 8027 59603
rect 8113 59547 8169 59603
rect 8255 59547 8311 59603
rect 8397 59547 8453 59603
rect 8539 59547 8595 59603
rect 8681 59547 8737 59603
rect 8823 59547 8879 59603
rect 8965 59547 9021 59603
rect 9107 59547 9163 59603
rect 9249 59547 9305 59603
rect 9391 59547 9447 59603
rect 9533 59547 9589 59603
rect 9675 59547 9731 59603
rect 9817 59547 9873 59603
rect 9959 59547 10015 59603
rect 10101 59547 10157 59603
rect 10243 59547 10299 59603
rect 10385 59547 10441 59603
rect 10527 59547 10583 59603
rect 10669 59547 10725 59603
rect 10811 59547 10867 59603
rect 10953 59547 11009 59603
rect 11095 59547 11151 59603
rect 11237 59547 11293 59603
rect 11379 59547 11435 59603
rect 11521 59547 11577 59603
rect 11663 59547 11719 59603
rect 11805 59547 11861 59603
rect 11947 59547 12003 59603
rect 12089 59547 12145 59603
rect 12231 59547 12287 59603
rect 12373 59547 12429 59603
rect 12515 59547 12571 59603
rect 12657 59547 12713 59603
rect 12799 59547 12855 59603
rect 12941 59547 12997 59603
rect 13083 59547 13139 59603
rect 13225 59547 13281 59603
rect 13367 59547 13423 59603
rect 13509 59547 13565 59603
rect 13651 59547 13707 59603
rect 13793 59547 13849 59603
rect 13935 59547 13991 59603
rect 14077 59547 14133 59603
rect 14219 59547 14275 59603
rect 14361 59547 14417 59603
rect 14503 59547 14559 59603
rect 14645 59547 14701 59603
rect 14787 59547 14843 59603
rect 161 59405 217 59461
rect 303 59405 359 59461
rect 445 59405 501 59461
rect 587 59405 643 59461
rect 729 59405 785 59461
rect 871 59405 927 59461
rect 1013 59405 1069 59461
rect 1155 59405 1211 59461
rect 1297 59405 1353 59461
rect 1439 59405 1495 59461
rect 1581 59405 1637 59461
rect 1723 59405 1779 59461
rect 1865 59405 1921 59461
rect 2007 59405 2063 59461
rect 2149 59405 2205 59461
rect 2291 59405 2347 59461
rect 2433 59405 2489 59461
rect 2575 59405 2631 59461
rect 2717 59405 2773 59461
rect 2859 59405 2915 59461
rect 3001 59405 3057 59461
rect 3143 59405 3199 59461
rect 3285 59405 3341 59461
rect 3427 59405 3483 59461
rect 3569 59405 3625 59461
rect 3711 59405 3767 59461
rect 3853 59405 3909 59461
rect 3995 59405 4051 59461
rect 4137 59405 4193 59461
rect 4279 59405 4335 59461
rect 4421 59405 4477 59461
rect 4563 59405 4619 59461
rect 4705 59405 4761 59461
rect 4847 59405 4903 59461
rect 4989 59405 5045 59461
rect 5131 59405 5187 59461
rect 5273 59405 5329 59461
rect 5415 59405 5471 59461
rect 5557 59405 5613 59461
rect 5699 59405 5755 59461
rect 5841 59405 5897 59461
rect 5983 59405 6039 59461
rect 6125 59405 6181 59461
rect 6267 59405 6323 59461
rect 6409 59405 6465 59461
rect 6551 59405 6607 59461
rect 6693 59405 6749 59461
rect 6835 59405 6891 59461
rect 6977 59405 7033 59461
rect 7119 59405 7175 59461
rect 7261 59405 7317 59461
rect 7403 59405 7459 59461
rect 7545 59405 7601 59461
rect 7687 59405 7743 59461
rect 7829 59405 7885 59461
rect 7971 59405 8027 59461
rect 8113 59405 8169 59461
rect 8255 59405 8311 59461
rect 8397 59405 8453 59461
rect 8539 59405 8595 59461
rect 8681 59405 8737 59461
rect 8823 59405 8879 59461
rect 8965 59405 9021 59461
rect 9107 59405 9163 59461
rect 9249 59405 9305 59461
rect 9391 59405 9447 59461
rect 9533 59405 9589 59461
rect 9675 59405 9731 59461
rect 9817 59405 9873 59461
rect 9959 59405 10015 59461
rect 10101 59405 10157 59461
rect 10243 59405 10299 59461
rect 10385 59405 10441 59461
rect 10527 59405 10583 59461
rect 10669 59405 10725 59461
rect 10811 59405 10867 59461
rect 10953 59405 11009 59461
rect 11095 59405 11151 59461
rect 11237 59405 11293 59461
rect 11379 59405 11435 59461
rect 11521 59405 11577 59461
rect 11663 59405 11719 59461
rect 11805 59405 11861 59461
rect 11947 59405 12003 59461
rect 12089 59405 12145 59461
rect 12231 59405 12287 59461
rect 12373 59405 12429 59461
rect 12515 59405 12571 59461
rect 12657 59405 12713 59461
rect 12799 59405 12855 59461
rect 12941 59405 12997 59461
rect 13083 59405 13139 59461
rect 13225 59405 13281 59461
rect 13367 59405 13423 59461
rect 13509 59405 13565 59461
rect 13651 59405 13707 59461
rect 13793 59405 13849 59461
rect 13935 59405 13991 59461
rect 14077 59405 14133 59461
rect 14219 59405 14275 59461
rect 14361 59405 14417 59461
rect 14503 59405 14559 59461
rect 14645 59405 14701 59461
rect 14787 59405 14843 59461
rect 161 59263 217 59319
rect 303 59263 359 59319
rect 445 59263 501 59319
rect 587 59263 643 59319
rect 729 59263 785 59319
rect 871 59263 927 59319
rect 1013 59263 1069 59319
rect 1155 59263 1211 59319
rect 1297 59263 1353 59319
rect 1439 59263 1495 59319
rect 1581 59263 1637 59319
rect 1723 59263 1779 59319
rect 1865 59263 1921 59319
rect 2007 59263 2063 59319
rect 2149 59263 2205 59319
rect 2291 59263 2347 59319
rect 2433 59263 2489 59319
rect 2575 59263 2631 59319
rect 2717 59263 2773 59319
rect 2859 59263 2915 59319
rect 3001 59263 3057 59319
rect 3143 59263 3199 59319
rect 3285 59263 3341 59319
rect 3427 59263 3483 59319
rect 3569 59263 3625 59319
rect 3711 59263 3767 59319
rect 3853 59263 3909 59319
rect 3995 59263 4051 59319
rect 4137 59263 4193 59319
rect 4279 59263 4335 59319
rect 4421 59263 4477 59319
rect 4563 59263 4619 59319
rect 4705 59263 4761 59319
rect 4847 59263 4903 59319
rect 4989 59263 5045 59319
rect 5131 59263 5187 59319
rect 5273 59263 5329 59319
rect 5415 59263 5471 59319
rect 5557 59263 5613 59319
rect 5699 59263 5755 59319
rect 5841 59263 5897 59319
rect 5983 59263 6039 59319
rect 6125 59263 6181 59319
rect 6267 59263 6323 59319
rect 6409 59263 6465 59319
rect 6551 59263 6607 59319
rect 6693 59263 6749 59319
rect 6835 59263 6891 59319
rect 6977 59263 7033 59319
rect 7119 59263 7175 59319
rect 7261 59263 7317 59319
rect 7403 59263 7459 59319
rect 7545 59263 7601 59319
rect 7687 59263 7743 59319
rect 7829 59263 7885 59319
rect 7971 59263 8027 59319
rect 8113 59263 8169 59319
rect 8255 59263 8311 59319
rect 8397 59263 8453 59319
rect 8539 59263 8595 59319
rect 8681 59263 8737 59319
rect 8823 59263 8879 59319
rect 8965 59263 9021 59319
rect 9107 59263 9163 59319
rect 9249 59263 9305 59319
rect 9391 59263 9447 59319
rect 9533 59263 9589 59319
rect 9675 59263 9731 59319
rect 9817 59263 9873 59319
rect 9959 59263 10015 59319
rect 10101 59263 10157 59319
rect 10243 59263 10299 59319
rect 10385 59263 10441 59319
rect 10527 59263 10583 59319
rect 10669 59263 10725 59319
rect 10811 59263 10867 59319
rect 10953 59263 11009 59319
rect 11095 59263 11151 59319
rect 11237 59263 11293 59319
rect 11379 59263 11435 59319
rect 11521 59263 11577 59319
rect 11663 59263 11719 59319
rect 11805 59263 11861 59319
rect 11947 59263 12003 59319
rect 12089 59263 12145 59319
rect 12231 59263 12287 59319
rect 12373 59263 12429 59319
rect 12515 59263 12571 59319
rect 12657 59263 12713 59319
rect 12799 59263 12855 59319
rect 12941 59263 12997 59319
rect 13083 59263 13139 59319
rect 13225 59263 13281 59319
rect 13367 59263 13423 59319
rect 13509 59263 13565 59319
rect 13651 59263 13707 59319
rect 13793 59263 13849 59319
rect 13935 59263 13991 59319
rect 14077 59263 14133 59319
rect 14219 59263 14275 59319
rect 14361 59263 14417 59319
rect 14503 59263 14559 59319
rect 14645 59263 14701 59319
rect 14787 59263 14843 59319
rect 161 59121 217 59177
rect 303 59121 359 59177
rect 445 59121 501 59177
rect 587 59121 643 59177
rect 729 59121 785 59177
rect 871 59121 927 59177
rect 1013 59121 1069 59177
rect 1155 59121 1211 59177
rect 1297 59121 1353 59177
rect 1439 59121 1495 59177
rect 1581 59121 1637 59177
rect 1723 59121 1779 59177
rect 1865 59121 1921 59177
rect 2007 59121 2063 59177
rect 2149 59121 2205 59177
rect 2291 59121 2347 59177
rect 2433 59121 2489 59177
rect 2575 59121 2631 59177
rect 2717 59121 2773 59177
rect 2859 59121 2915 59177
rect 3001 59121 3057 59177
rect 3143 59121 3199 59177
rect 3285 59121 3341 59177
rect 3427 59121 3483 59177
rect 3569 59121 3625 59177
rect 3711 59121 3767 59177
rect 3853 59121 3909 59177
rect 3995 59121 4051 59177
rect 4137 59121 4193 59177
rect 4279 59121 4335 59177
rect 4421 59121 4477 59177
rect 4563 59121 4619 59177
rect 4705 59121 4761 59177
rect 4847 59121 4903 59177
rect 4989 59121 5045 59177
rect 5131 59121 5187 59177
rect 5273 59121 5329 59177
rect 5415 59121 5471 59177
rect 5557 59121 5613 59177
rect 5699 59121 5755 59177
rect 5841 59121 5897 59177
rect 5983 59121 6039 59177
rect 6125 59121 6181 59177
rect 6267 59121 6323 59177
rect 6409 59121 6465 59177
rect 6551 59121 6607 59177
rect 6693 59121 6749 59177
rect 6835 59121 6891 59177
rect 6977 59121 7033 59177
rect 7119 59121 7175 59177
rect 7261 59121 7317 59177
rect 7403 59121 7459 59177
rect 7545 59121 7601 59177
rect 7687 59121 7743 59177
rect 7829 59121 7885 59177
rect 7971 59121 8027 59177
rect 8113 59121 8169 59177
rect 8255 59121 8311 59177
rect 8397 59121 8453 59177
rect 8539 59121 8595 59177
rect 8681 59121 8737 59177
rect 8823 59121 8879 59177
rect 8965 59121 9021 59177
rect 9107 59121 9163 59177
rect 9249 59121 9305 59177
rect 9391 59121 9447 59177
rect 9533 59121 9589 59177
rect 9675 59121 9731 59177
rect 9817 59121 9873 59177
rect 9959 59121 10015 59177
rect 10101 59121 10157 59177
rect 10243 59121 10299 59177
rect 10385 59121 10441 59177
rect 10527 59121 10583 59177
rect 10669 59121 10725 59177
rect 10811 59121 10867 59177
rect 10953 59121 11009 59177
rect 11095 59121 11151 59177
rect 11237 59121 11293 59177
rect 11379 59121 11435 59177
rect 11521 59121 11577 59177
rect 11663 59121 11719 59177
rect 11805 59121 11861 59177
rect 11947 59121 12003 59177
rect 12089 59121 12145 59177
rect 12231 59121 12287 59177
rect 12373 59121 12429 59177
rect 12515 59121 12571 59177
rect 12657 59121 12713 59177
rect 12799 59121 12855 59177
rect 12941 59121 12997 59177
rect 13083 59121 13139 59177
rect 13225 59121 13281 59177
rect 13367 59121 13423 59177
rect 13509 59121 13565 59177
rect 13651 59121 13707 59177
rect 13793 59121 13849 59177
rect 13935 59121 13991 59177
rect 14077 59121 14133 59177
rect 14219 59121 14275 59177
rect 14361 59121 14417 59177
rect 14503 59121 14559 59177
rect 14645 59121 14701 59177
rect 14787 59121 14843 59177
rect 161 58979 217 59035
rect 303 58979 359 59035
rect 445 58979 501 59035
rect 587 58979 643 59035
rect 729 58979 785 59035
rect 871 58979 927 59035
rect 1013 58979 1069 59035
rect 1155 58979 1211 59035
rect 1297 58979 1353 59035
rect 1439 58979 1495 59035
rect 1581 58979 1637 59035
rect 1723 58979 1779 59035
rect 1865 58979 1921 59035
rect 2007 58979 2063 59035
rect 2149 58979 2205 59035
rect 2291 58979 2347 59035
rect 2433 58979 2489 59035
rect 2575 58979 2631 59035
rect 2717 58979 2773 59035
rect 2859 58979 2915 59035
rect 3001 58979 3057 59035
rect 3143 58979 3199 59035
rect 3285 58979 3341 59035
rect 3427 58979 3483 59035
rect 3569 58979 3625 59035
rect 3711 58979 3767 59035
rect 3853 58979 3909 59035
rect 3995 58979 4051 59035
rect 4137 58979 4193 59035
rect 4279 58979 4335 59035
rect 4421 58979 4477 59035
rect 4563 58979 4619 59035
rect 4705 58979 4761 59035
rect 4847 58979 4903 59035
rect 4989 58979 5045 59035
rect 5131 58979 5187 59035
rect 5273 58979 5329 59035
rect 5415 58979 5471 59035
rect 5557 58979 5613 59035
rect 5699 58979 5755 59035
rect 5841 58979 5897 59035
rect 5983 58979 6039 59035
rect 6125 58979 6181 59035
rect 6267 58979 6323 59035
rect 6409 58979 6465 59035
rect 6551 58979 6607 59035
rect 6693 58979 6749 59035
rect 6835 58979 6891 59035
rect 6977 58979 7033 59035
rect 7119 58979 7175 59035
rect 7261 58979 7317 59035
rect 7403 58979 7459 59035
rect 7545 58979 7601 59035
rect 7687 58979 7743 59035
rect 7829 58979 7885 59035
rect 7971 58979 8027 59035
rect 8113 58979 8169 59035
rect 8255 58979 8311 59035
rect 8397 58979 8453 59035
rect 8539 58979 8595 59035
rect 8681 58979 8737 59035
rect 8823 58979 8879 59035
rect 8965 58979 9021 59035
rect 9107 58979 9163 59035
rect 9249 58979 9305 59035
rect 9391 58979 9447 59035
rect 9533 58979 9589 59035
rect 9675 58979 9731 59035
rect 9817 58979 9873 59035
rect 9959 58979 10015 59035
rect 10101 58979 10157 59035
rect 10243 58979 10299 59035
rect 10385 58979 10441 59035
rect 10527 58979 10583 59035
rect 10669 58979 10725 59035
rect 10811 58979 10867 59035
rect 10953 58979 11009 59035
rect 11095 58979 11151 59035
rect 11237 58979 11293 59035
rect 11379 58979 11435 59035
rect 11521 58979 11577 59035
rect 11663 58979 11719 59035
rect 11805 58979 11861 59035
rect 11947 58979 12003 59035
rect 12089 58979 12145 59035
rect 12231 58979 12287 59035
rect 12373 58979 12429 59035
rect 12515 58979 12571 59035
rect 12657 58979 12713 59035
rect 12799 58979 12855 59035
rect 12941 58979 12997 59035
rect 13083 58979 13139 59035
rect 13225 58979 13281 59035
rect 13367 58979 13423 59035
rect 13509 58979 13565 59035
rect 13651 58979 13707 59035
rect 13793 58979 13849 59035
rect 13935 58979 13991 59035
rect 14077 58979 14133 59035
rect 14219 58979 14275 59035
rect 14361 58979 14417 59035
rect 14503 58979 14559 59035
rect 14645 58979 14701 59035
rect 14787 58979 14843 59035
rect 161 58837 217 58893
rect 303 58837 359 58893
rect 445 58837 501 58893
rect 587 58837 643 58893
rect 729 58837 785 58893
rect 871 58837 927 58893
rect 1013 58837 1069 58893
rect 1155 58837 1211 58893
rect 1297 58837 1353 58893
rect 1439 58837 1495 58893
rect 1581 58837 1637 58893
rect 1723 58837 1779 58893
rect 1865 58837 1921 58893
rect 2007 58837 2063 58893
rect 2149 58837 2205 58893
rect 2291 58837 2347 58893
rect 2433 58837 2489 58893
rect 2575 58837 2631 58893
rect 2717 58837 2773 58893
rect 2859 58837 2915 58893
rect 3001 58837 3057 58893
rect 3143 58837 3199 58893
rect 3285 58837 3341 58893
rect 3427 58837 3483 58893
rect 3569 58837 3625 58893
rect 3711 58837 3767 58893
rect 3853 58837 3909 58893
rect 3995 58837 4051 58893
rect 4137 58837 4193 58893
rect 4279 58837 4335 58893
rect 4421 58837 4477 58893
rect 4563 58837 4619 58893
rect 4705 58837 4761 58893
rect 4847 58837 4903 58893
rect 4989 58837 5045 58893
rect 5131 58837 5187 58893
rect 5273 58837 5329 58893
rect 5415 58837 5471 58893
rect 5557 58837 5613 58893
rect 5699 58837 5755 58893
rect 5841 58837 5897 58893
rect 5983 58837 6039 58893
rect 6125 58837 6181 58893
rect 6267 58837 6323 58893
rect 6409 58837 6465 58893
rect 6551 58837 6607 58893
rect 6693 58837 6749 58893
rect 6835 58837 6891 58893
rect 6977 58837 7033 58893
rect 7119 58837 7175 58893
rect 7261 58837 7317 58893
rect 7403 58837 7459 58893
rect 7545 58837 7601 58893
rect 7687 58837 7743 58893
rect 7829 58837 7885 58893
rect 7971 58837 8027 58893
rect 8113 58837 8169 58893
rect 8255 58837 8311 58893
rect 8397 58837 8453 58893
rect 8539 58837 8595 58893
rect 8681 58837 8737 58893
rect 8823 58837 8879 58893
rect 8965 58837 9021 58893
rect 9107 58837 9163 58893
rect 9249 58837 9305 58893
rect 9391 58837 9447 58893
rect 9533 58837 9589 58893
rect 9675 58837 9731 58893
rect 9817 58837 9873 58893
rect 9959 58837 10015 58893
rect 10101 58837 10157 58893
rect 10243 58837 10299 58893
rect 10385 58837 10441 58893
rect 10527 58837 10583 58893
rect 10669 58837 10725 58893
rect 10811 58837 10867 58893
rect 10953 58837 11009 58893
rect 11095 58837 11151 58893
rect 11237 58837 11293 58893
rect 11379 58837 11435 58893
rect 11521 58837 11577 58893
rect 11663 58837 11719 58893
rect 11805 58837 11861 58893
rect 11947 58837 12003 58893
rect 12089 58837 12145 58893
rect 12231 58837 12287 58893
rect 12373 58837 12429 58893
rect 12515 58837 12571 58893
rect 12657 58837 12713 58893
rect 12799 58837 12855 58893
rect 12941 58837 12997 58893
rect 13083 58837 13139 58893
rect 13225 58837 13281 58893
rect 13367 58837 13423 58893
rect 13509 58837 13565 58893
rect 13651 58837 13707 58893
rect 13793 58837 13849 58893
rect 13935 58837 13991 58893
rect 14077 58837 14133 58893
rect 14219 58837 14275 58893
rect 14361 58837 14417 58893
rect 14503 58837 14559 58893
rect 14645 58837 14701 58893
rect 14787 58837 14843 58893
rect 161 58507 217 58563
rect 303 58507 359 58563
rect 445 58507 501 58563
rect 587 58507 643 58563
rect 729 58507 785 58563
rect 871 58507 927 58563
rect 1013 58507 1069 58563
rect 1155 58507 1211 58563
rect 1297 58507 1353 58563
rect 1439 58507 1495 58563
rect 1581 58507 1637 58563
rect 1723 58507 1779 58563
rect 1865 58507 1921 58563
rect 2007 58507 2063 58563
rect 2149 58507 2205 58563
rect 2291 58507 2347 58563
rect 2433 58507 2489 58563
rect 2575 58507 2631 58563
rect 2717 58507 2773 58563
rect 2859 58507 2915 58563
rect 3001 58507 3057 58563
rect 3143 58507 3199 58563
rect 3285 58507 3341 58563
rect 3427 58507 3483 58563
rect 3569 58507 3625 58563
rect 3711 58507 3767 58563
rect 3853 58507 3909 58563
rect 3995 58507 4051 58563
rect 4137 58507 4193 58563
rect 4279 58507 4335 58563
rect 4421 58507 4477 58563
rect 4563 58507 4619 58563
rect 4705 58507 4761 58563
rect 4847 58507 4903 58563
rect 4989 58507 5045 58563
rect 5131 58507 5187 58563
rect 5273 58507 5329 58563
rect 5415 58507 5471 58563
rect 5557 58507 5613 58563
rect 5699 58507 5755 58563
rect 5841 58507 5897 58563
rect 5983 58507 6039 58563
rect 6125 58507 6181 58563
rect 6267 58507 6323 58563
rect 6409 58507 6465 58563
rect 6551 58507 6607 58563
rect 6693 58507 6749 58563
rect 6835 58507 6891 58563
rect 6977 58507 7033 58563
rect 7119 58507 7175 58563
rect 7261 58507 7317 58563
rect 7403 58507 7459 58563
rect 7545 58507 7601 58563
rect 7687 58507 7743 58563
rect 7829 58507 7885 58563
rect 7971 58507 8027 58563
rect 8113 58507 8169 58563
rect 8255 58507 8311 58563
rect 8397 58507 8453 58563
rect 8539 58507 8595 58563
rect 8681 58507 8737 58563
rect 8823 58507 8879 58563
rect 8965 58507 9021 58563
rect 9107 58507 9163 58563
rect 9249 58507 9305 58563
rect 9391 58507 9447 58563
rect 9533 58507 9589 58563
rect 9675 58507 9731 58563
rect 9817 58507 9873 58563
rect 9959 58507 10015 58563
rect 10101 58507 10157 58563
rect 10243 58507 10299 58563
rect 10385 58507 10441 58563
rect 10527 58507 10583 58563
rect 10669 58507 10725 58563
rect 10811 58507 10867 58563
rect 10953 58507 11009 58563
rect 11095 58507 11151 58563
rect 11237 58507 11293 58563
rect 11379 58507 11435 58563
rect 11521 58507 11577 58563
rect 11663 58507 11719 58563
rect 11805 58507 11861 58563
rect 11947 58507 12003 58563
rect 12089 58507 12145 58563
rect 12231 58507 12287 58563
rect 12373 58507 12429 58563
rect 12515 58507 12571 58563
rect 12657 58507 12713 58563
rect 12799 58507 12855 58563
rect 12941 58507 12997 58563
rect 13083 58507 13139 58563
rect 13225 58507 13281 58563
rect 13367 58507 13423 58563
rect 13509 58507 13565 58563
rect 13651 58507 13707 58563
rect 13793 58507 13849 58563
rect 13935 58507 13991 58563
rect 14077 58507 14133 58563
rect 14219 58507 14275 58563
rect 14361 58507 14417 58563
rect 14503 58507 14559 58563
rect 14645 58507 14701 58563
rect 14787 58507 14843 58563
rect 161 58365 217 58421
rect 303 58365 359 58421
rect 445 58365 501 58421
rect 587 58365 643 58421
rect 729 58365 785 58421
rect 871 58365 927 58421
rect 1013 58365 1069 58421
rect 1155 58365 1211 58421
rect 1297 58365 1353 58421
rect 1439 58365 1495 58421
rect 1581 58365 1637 58421
rect 1723 58365 1779 58421
rect 1865 58365 1921 58421
rect 2007 58365 2063 58421
rect 2149 58365 2205 58421
rect 2291 58365 2347 58421
rect 2433 58365 2489 58421
rect 2575 58365 2631 58421
rect 2717 58365 2773 58421
rect 2859 58365 2915 58421
rect 3001 58365 3057 58421
rect 3143 58365 3199 58421
rect 3285 58365 3341 58421
rect 3427 58365 3483 58421
rect 3569 58365 3625 58421
rect 3711 58365 3767 58421
rect 3853 58365 3909 58421
rect 3995 58365 4051 58421
rect 4137 58365 4193 58421
rect 4279 58365 4335 58421
rect 4421 58365 4477 58421
rect 4563 58365 4619 58421
rect 4705 58365 4761 58421
rect 4847 58365 4903 58421
rect 4989 58365 5045 58421
rect 5131 58365 5187 58421
rect 5273 58365 5329 58421
rect 5415 58365 5471 58421
rect 5557 58365 5613 58421
rect 5699 58365 5755 58421
rect 5841 58365 5897 58421
rect 5983 58365 6039 58421
rect 6125 58365 6181 58421
rect 6267 58365 6323 58421
rect 6409 58365 6465 58421
rect 6551 58365 6607 58421
rect 6693 58365 6749 58421
rect 6835 58365 6891 58421
rect 6977 58365 7033 58421
rect 7119 58365 7175 58421
rect 7261 58365 7317 58421
rect 7403 58365 7459 58421
rect 7545 58365 7601 58421
rect 7687 58365 7743 58421
rect 7829 58365 7885 58421
rect 7971 58365 8027 58421
rect 8113 58365 8169 58421
rect 8255 58365 8311 58421
rect 8397 58365 8453 58421
rect 8539 58365 8595 58421
rect 8681 58365 8737 58421
rect 8823 58365 8879 58421
rect 8965 58365 9021 58421
rect 9107 58365 9163 58421
rect 9249 58365 9305 58421
rect 9391 58365 9447 58421
rect 9533 58365 9589 58421
rect 9675 58365 9731 58421
rect 9817 58365 9873 58421
rect 9959 58365 10015 58421
rect 10101 58365 10157 58421
rect 10243 58365 10299 58421
rect 10385 58365 10441 58421
rect 10527 58365 10583 58421
rect 10669 58365 10725 58421
rect 10811 58365 10867 58421
rect 10953 58365 11009 58421
rect 11095 58365 11151 58421
rect 11237 58365 11293 58421
rect 11379 58365 11435 58421
rect 11521 58365 11577 58421
rect 11663 58365 11719 58421
rect 11805 58365 11861 58421
rect 11947 58365 12003 58421
rect 12089 58365 12145 58421
rect 12231 58365 12287 58421
rect 12373 58365 12429 58421
rect 12515 58365 12571 58421
rect 12657 58365 12713 58421
rect 12799 58365 12855 58421
rect 12941 58365 12997 58421
rect 13083 58365 13139 58421
rect 13225 58365 13281 58421
rect 13367 58365 13423 58421
rect 13509 58365 13565 58421
rect 13651 58365 13707 58421
rect 13793 58365 13849 58421
rect 13935 58365 13991 58421
rect 14077 58365 14133 58421
rect 14219 58365 14275 58421
rect 14361 58365 14417 58421
rect 14503 58365 14559 58421
rect 14645 58365 14701 58421
rect 14787 58365 14843 58421
rect 161 58223 217 58279
rect 303 58223 359 58279
rect 445 58223 501 58279
rect 587 58223 643 58279
rect 729 58223 785 58279
rect 871 58223 927 58279
rect 1013 58223 1069 58279
rect 1155 58223 1211 58279
rect 1297 58223 1353 58279
rect 1439 58223 1495 58279
rect 1581 58223 1637 58279
rect 1723 58223 1779 58279
rect 1865 58223 1921 58279
rect 2007 58223 2063 58279
rect 2149 58223 2205 58279
rect 2291 58223 2347 58279
rect 2433 58223 2489 58279
rect 2575 58223 2631 58279
rect 2717 58223 2773 58279
rect 2859 58223 2915 58279
rect 3001 58223 3057 58279
rect 3143 58223 3199 58279
rect 3285 58223 3341 58279
rect 3427 58223 3483 58279
rect 3569 58223 3625 58279
rect 3711 58223 3767 58279
rect 3853 58223 3909 58279
rect 3995 58223 4051 58279
rect 4137 58223 4193 58279
rect 4279 58223 4335 58279
rect 4421 58223 4477 58279
rect 4563 58223 4619 58279
rect 4705 58223 4761 58279
rect 4847 58223 4903 58279
rect 4989 58223 5045 58279
rect 5131 58223 5187 58279
rect 5273 58223 5329 58279
rect 5415 58223 5471 58279
rect 5557 58223 5613 58279
rect 5699 58223 5755 58279
rect 5841 58223 5897 58279
rect 5983 58223 6039 58279
rect 6125 58223 6181 58279
rect 6267 58223 6323 58279
rect 6409 58223 6465 58279
rect 6551 58223 6607 58279
rect 6693 58223 6749 58279
rect 6835 58223 6891 58279
rect 6977 58223 7033 58279
rect 7119 58223 7175 58279
rect 7261 58223 7317 58279
rect 7403 58223 7459 58279
rect 7545 58223 7601 58279
rect 7687 58223 7743 58279
rect 7829 58223 7885 58279
rect 7971 58223 8027 58279
rect 8113 58223 8169 58279
rect 8255 58223 8311 58279
rect 8397 58223 8453 58279
rect 8539 58223 8595 58279
rect 8681 58223 8737 58279
rect 8823 58223 8879 58279
rect 8965 58223 9021 58279
rect 9107 58223 9163 58279
rect 9249 58223 9305 58279
rect 9391 58223 9447 58279
rect 9533 58223 9589 58279
rect 9675 58223 9731 58279
rect 9817 58223 9873 58279
rect 9959 58223 10015 58279
rect 10101 58223 10157 58279
rect 10243 58223 10299 58279
rect 10385 58223 10441 58279
rect 10527 58223 10583 58279
rect 10669 58223 10725 58279
rect 10811 58223 10867 58279
rect 10953 58223 11009 58279
rect 11095 58223 11151 58279
rect 11237 58223 11293 58279
rect 11379 58223 11435 58279
rect 11521 58223 11577 58279
rect 11663 58223 11719 58279
rect 11805 58223 11861 58279
rect 11947 58223 12003 58279
rect 12089 58223 12145 58279
rect 12231 58223 12287 58279
rect 12373 58223 12429 58279
rect 12515 58223 12571 58279
rect 12657 58223 12713 58279
rect 12799 58223 12855 58279
rect 12941 58223 12997 58279
rect 13083 58223 13139 58279
rect 13225 58223 13281 58279
rect 13367 58223 13423 58279
rect 13509 58223 13565 58279
rect 13651 58223 13707 58279
rect 13793 58223 13849 58279
rect 13935 58223 13991 58279
rect 14077 58223 14133 58279
rect 14219 58223 14275 58279
rect 14361 58223 14417 58279
rect 14503 58223 14559 58279
rect 14645 58223 14701 58279
rect 14787 58223 14843 58279
rect 161 58081 217 58137
rect 303 58081 359 58137
rect 445 58081 501 58137
rect 587 58081 643 58137
rect 729 58081 785 58137
rect 871 58081 927 58137
rect 1013 58081 1069 58137
rect 1155 58081 1211 58137
rect 1297 58081 1353 58137
rect 1439 58081 1495 58137
rect 1581 58081 1637 58137
rect 1723 58081 1779 58137
rect 1865 58081 1921 58137
rect 2007 58081 2063 58137
rect 2149 58081 2205 58137
rect 2291 58081 2347 58137
rect 2433 58081 2489 58137
rect 2575 58081 2631 58137
rect 2717 58081 2773 58137
rect 2859 58081 2915 58137
rect 3001 58081 3057 58137
rect 3143 58081 3199 58137
rect 3285 58081 3341 58137
rect 3427 58081 3483 58137
rect 3569 58081 3625 58137
rect 3711 58081 3767 58137
rect 3853 58081 3909 58137
rect 3995 58081 4051 58137
rect 4137 58081 4193 58137
rect 4279 58081 4335 58137
rect 4421 58081 4477 58137
rect 4563 58081 4619 58137
rect 4705 58081 4761 58137
rect 4847 58081 4903 58137
rect 4989 58081 5045 58137
rect 5131 58081 5187 58137
rect 5273 58081 5329 58137
rect 5415 58081 5471 58137
rect 5557 58081 5613 58137
rect 5699 58081 5755 58137
rect 5841 58081 5897 58137
rect 5983 58081 6039 58137
rect 6125 58081 6181 58137
rect 6267 58081 6323 58137
rect 6409 58081 6465 58137
rect 6551 58081 6607 58137
rect 6693 58081 6749 58137
rect 6835 58081 6891 58137
rect 6977 58081 7033 58137
rect 7119 58081 7175 58137
rect 7261 58081 7317 58137
rect 7403 58081 7459 58137
rect 7545 58081 7601 58137
rect 7687 58081 7743 58137
rect 7829 58081 7885 58137
rect 7971 58081 8027 58137
rect 8113 58081 8169 58137
rect 8255 58081 8311 58137
rect 8397 58081 8453 58137
rect 8539 58081 8595 58137
rect 8681 58081 8737 58137
rect 8823 58081 8879 58137
rect 8965 58081 9021 58137
rect 9107 58081 9163 58137
rect 9249 58081 9305 58137
rect 9391 58081 9447 58137
rect 9533 58081 9589 58137
rect 9675 58081 9731 58137
rect 9817 58081 9873 58137
rect 9959 58081 10015 58137
rect 10101 58081 10157 58137
rect 10243 58081 10299 58137
rect 10385 58081 10441 58137
rect 10527 58081 10583 58137
rect 10669 58081 10725 58137
rect 10811 58081 10867 58137
rect 10953 58081 11009 58137
rect 11095 58081 11151 58137
rect 11237 58081 11293 58137
rect 11379 58081 11435 58137
rect 11521 58081 11577 58137
rect 11663 58081 11719 58137
rect 11805 58081 11861 58137
rect 11947 58081 12003 58137
rect 12089 58081 12145 58137
rect 12231 58081 12287 58137
rect 12373 58081 12429 58137
rect 12515 58081 12571 58137
rect 12657 58081 12713 58137
rect 12799 58081 12855 58137
rect 12941 58081 12997 58137
rect 13083 58081 13139 58137
rect 13225 58081 13281 58137
rect 13367 58081 13423 58137
rect 13509 58081 13565 58137
rect 13651 58081 13707 58137
rect 13793 58081 13849 58137
rect 13935 58081 13991 58137
rect 14077 58081 14133 58137
rect 14219 58081 14275 58137
rect 14361 58081 14417 58137
rect 14503 58081 14559 58137
rect 14645 58081 14701 58137
rect 14787 58081 14843 58137
rect 161 57939 217 57995
rect 303 57939 359 57995
rect 445 57939 501 57995
rect 587 57939 643 57995
rect 729 57939 785 57995
rect 871 57939 927 57995
rect 1013 57939 1069 57995
rect 1155 57939 1211 57995
rect 1297 57939 1353 57995
rect 1439 57939 1495 57995
rect 1581 57939 1637 57995
rect 1723 57939 1779 57995
rect 1865 57939 1921 57995
rect 2007 57939 2063 57995
rect 2149 57939 2205 57995
rect 2291 57939 2347 57995
rect 2433 57939 2489 57995
rect 2575 57939 2631 57995
rect 2717 57939 2773 57995
rect 2859 57939 2915 57995
rect 3001 57939 3057 57995
rect 3143 57939 3199 57995
rect 3285 57939 3341 57995
rect 3427 57939 3483 57995
rect 3569 57939 3625 57995
rect 3711 57939 3767 57995
rect 3853 57939 3909 57995
rect 3995 57939 4051 57995
rect 4137 57939 4193 57995
rect 4279 57939 4335 57995
rect 4421 57939 4477 57995
rect 4563 57939 4619 57995
rect 4705 57939 4761 57995
rect 4847 57939 4903 57995
rect 4989 57939 5045 57995
rect 5131 57939 5187 57995
rect 5273 57939 5329 57995
rect 5415 57939 5471 57995
rect 5557 57939 5613 57995
rect 5699 57939 5755 57995
rect 5841 57939 5897 57995
rect 5983 57939 6039 57995
rect 6125 57939 6181 57995
rect 6267 57939 6323 57995
rect 6409 57939 6465 57995
rect 6551 57939 6607 57995
rect 6693 57939 6749 57995
rect 6835 57939 6891 57995
rect 6977 57939 7033 57995
rect 7119 57939 7175 57995
rect 7261 57939 7317 57995
rect 7403 57939 7459 57995
rect 7545 57939 7601 57995
rect 7687 57939 7743 57995
rect 7829 57939 7885 57995
rect 7971 57939 8027 57995
rect 8113 57939 8169 57995
rect 8255 57939 8311 57995
rect 8397 57939 8453 57995
rect 8539 57939 8595 57995
rect 8681 57939 8737 57995
rect 8823 57939 8879 57995
rect 8965 57939 9021 57995
rect 9107 57939 9163 57995
rect 9249 57939 9305 57995
rect 9391 57939 9447 57995
rect 9533 57939 9589 57995
rect 9675 57939 9731 57995
rect 9817 57939 9873 57995
rect 9959 57939 10015 57995
rect 10101 57939 10157 57995
rect 10243 57939 10299 57995
rect 10385 57939 10441 57995
rect 10527 57939 10583 57995
rect 10669 57939 10725 57995
rect 10811 57939 10867 57995
rect 10953 57939 11009 57995
rect 11095 57939 11151 57995
rect 11237 57939 11293 57995
rect 11379 57939 11435 57995
rect 11521 57939 11577 57995
rect 11663 57939 11719 57995
rect 11805 57939 11861 57995
rect 11947 57939 12003 57995
rect 12089 57939 12145 57995
rect 12231 57939 12287 57995
rect 12373 57939 12429 57995
rect 12515 57939 12571 57995
rect 12657 57939 12713 57995
rect 12799 57939 12855 57995
rect 12941 57939 12997 57995
rect 13083 57939 13139 57995
rect 13225 57939 13281 57995
rect 13367 57939 13423 57995
rect 13509 57939 13565 57995
rect 13651 57939 13707 57995
rect 13793 57939 13849 57995
rect 13935 57939 13991 57995
rect 14077 57939 14133 57995
rect 14219 57939 14275 57995
rect 14361 57939 14417 57995
rect 14503 57939 14559 57995
rect 14645 57939 14701 57995
rect 14787 57939 14843 57995
rect 161 57797 217 57853
rect 303 57797 359 57853
rect 445 57797 501 57853
rect 587 57797 643 57853
rect 729 57797 785 57853
rect 871 57797 927 57853
rect 1013 57797 1069 57853
rect 1155 57797 1211 57853
rect 1297 57797 1353 57853
rect 1439 57797 1495 57853
rect 1581 57797 1637 57853
rect 1723 57797 1779 57853
rect 1865 57797 1921 57853
rect 2007 57797 2063 57853
rect 2149 57797 2205 57853
rect 2291 57797 2347 57853
rect 2433 57797 2489 57853
rect 2575 57797 2631 57853
rect 2717 57797 2773 57853
rect 2859 57797 2915 57853
rect 3001 57797 3057 57853
rect 3143 57797 3199 57853
rect 3285 57797 3341 57853
rect 3427 57797 3483 57853
rect 3569 57797 3625 57853
rect 3711 57797 3767 57853
rect 3853 57797 3909 57853
rect 3995 57797 4051 57853
rect 4137 57797 4193 57853
rect 4279 57797 4335 57853
rect 4421 57797 4477 57853
rect 4563 57797 4619 57853
rect 4705 57797 4761 57853
rect 4847 57797 4903 57853
rect 4989 57797 5045 57853
rect 5131 57797 5187 57853
rect 5273 57797 5329 57853
rect 5415 57797 5471 57853
rect 5557 57797 5613 57853
rect 5699 57797 5755 57853
rect 5841 57797 5897 57853
rect 5983 57797 6039 57853
rect 6125 57797 6181 57853
rect 6267 57797 6323 57853
rect 6409 57797 6465 57853
rect 6551 57797 6607 57853
rect 6693 57797 6749 57853
rect 6835 57797 6891 57853
rect 6977 57797 7033 57853
rect 7119 57797 7175 57853
rect 7261 57797 7317 57853
rect 7403 57797 7459 57853
rect 7545 57797 7601 57853
rect 7687 57797 7743 57853
rect 7829 57797 7885 57853
rect 7971 57797 8027 57853
rect 8113 57797 8169 57853
rect 8255 57797 8311 57853
rect 8397 57797 8453 57853
rect 8539 57797 8595 57853
rect 8681 57797 8737 57853
rect 8823 57797 8879 57853
rect 8965 57797 9021 57853
rect 9107 57797 9163 57853
rect 9249 57797 9305 57853
rect 9391 57797 9447 57853
rect 9533 57797 9589 57853
rect 9675 57797 9731 57853
rect 9817 57797 9873 57853
rect 9959 57797 10015 57853
rect 10101 57797 10157 57853
rect 10243 57797 10299 57853
rect 10385 57797 10441 57853
rect 10527 57797 10583 57853
rect 10669 57797 10725 57853
rect 10811 57797 10867 57853
rect 10953 57797 11009 57853
rect 11095 57797 11151 57853
rect 11237 57797 11293 57853
rect 11379 57797 11435 57853
rect 11521 57797 11577 57853
rect 11663 57797 11719 57853
rect 11805 57797 11861 57853
rect 11947 57797 12003 57853
rect 12089 57797 12145 57853
rect 12231 57797 12287 57853
rect 12373 57797 12429 57853
rect 12515 57797 12571 57853
rect 12657 57797 12713 57853
rect 12799 57797 12855 57853
rect 12941 57797 12997 57853
rect 13083 57797 13139 57853
rect 13225 57797 13281 57853
rect 13367 57797 13423 57853
rect 13509 57797 13565 57853
rect 13651 57797 13707 57853
rect 13793 57797 13849 57853
rect 13935 57797 13991 57853
rect 14077 57797 14133 57853
rect 14219 57797 14275 57853
rect 14361 57797 14417 57853
rect 14503 57797 14559 57853
rect 14645 57797 14701 57853
rect 14787 57797 14843 57853
rect 161 57655 217 57711
rect 303 57655 359 57711
rect 445 57655 501 57711
rect 587 57655 643 57711
rect 729 57655 785 57711
rect 871 57655 927 57711
rect 1013 57655 1069 57711
rect 1155 57655 1211 57711
rect 1297 57655 1353 57711
rect 1439 57655 1495 57711
rect 1581 57655 1637 57711
rect 1723 57655 1779 57711
rect 1865 57655 1921 57711
rect 2007 57655 2063 57711
rect 2149 57655 2205 57711
rect 2291 57655 2347 57711
rect 2433 57655 2489 57711
rect 2575 57655 2631 57711
rect 2717 57655 2773 57711
rect 2859 57655 2915 57711
rect 3001 57655 3057 57711
rect 3143 57655 3199 57711
rect 3285 57655 3341 57711
rect 3427 57655 3483 57711
rect 3569 57655 3625 57711
rect 3711 57655 3767 57711
rect 3853 57655 3909 57711
rect 3995 57655 4051 57711
rect 4137 57655 4193 57711
rect 4279 57655 4335 57711
rect 4421 57655 4477 57711
rect 4563 57655 4619 57711
rect 4705 57655 4761 57711
rect 4847 57655 4903 57711
rect 4989 57655 5045 57711
rect 5131 57655 5187 57711
rect 5273 57655 5329 57711
rect 5415 57655 5471 57711
rect 5557 57655 5613 57711
rect 5699 57655 5755 57711
rect 5841 57655 5897 57711
rect 5983 57655 6039 57711
rect 6125 57655 6181 57711
rect 6267 57655 6323 57711
rect 6409 57655 6465 57711
rect 6551 57655 6607 57711
rect 6693 57655 6749 57711
rect 6835 57655 6891 57711
rect 6977 57655 7033 57711
rect 7119 57655 7175 57711
rect 7261 57655 7317 57711
rect 7403 57655 7459 57711
rect 7545 57655 7601 57711
rect 7687 57655 7743 57711
rect 7829 57655 7885 57711
rect 7971 57655 8027 57711
rect 8113 57655 8169 57711
rect 8255 57655 8311 57711
rect 8397 57655 8453 57711
rect 8539 57655 8595 57711
rect 8681 57655 8737 57711
rect 8823 57655 8879 57711
rect 8965 57655 9021 57711
rect 9107 57655 9163 57711
rect 9249 57655 9305 57711
rect 9391 57655 9447 57711
rect 9533 57655 9589 57711
rect 9675 57655 9731 57711
rect 9817 57655 9873 57711
rect 9959 57655 10015 57711
rect 10101 57655 10157 57711
rect 10243 57655 10299 57711
rect 10385 57655 10441 57711
rect 10527 57655 10583 57711
rect 10669 57655 10725 57711
rect 10811 57655 10867 57711
rect 10953 57655 11009 57711
rect 11095 57655 11151 57711
rect 11237 57655 11293 57711
rect 11379 57655 11435 57711
rect 11521 57655 11577 57711
rect 11663 57655 11719 57711
rect 11805 57655 11861 57711
rect 11947 57655 12003 57711
rect 12089 57655 12145 57711
rect 12231 57655 12287 57711
rect 12373 57655 12429 57711
rect 12515 57655 12571 57711
rect 12657 57655 12713 57711
rect 12799 57655 12855 57711
rect 12941 57655 12997 57711
rect 13083 57655 13139 57711
rect 13225 57655 13281 57711
rect 13367 57655 13423 57711
rect 13509 57655 13565 57711
rect 13651 57655 13707 57711
rect 13793 57655 13849 57711
rect 13935 57655 13991 57711
rect 14077 57655 14133 57711
rect 14219 57655 14275 57711
rect 14361 57655 14417 57711
rect 14503 57655 14559 57711
rect 14645 57655 14701 57711
rect 14787 57655 14843 57711
rect 161 57513 217 57569
rect 303 57513 359 57569
rect 445 57513 501 57569
rect 587 57513 643 57569
rect 729 57513 785 57569
rect 871 57513 927 57569
rect 1013 57513 1069 57569
rect 1155 57513 1211 57569
rect 1297 57513 1353 57569
rect 1439 57513 1495 57569
rect 1581 57513 1637 57569
rect 1723 57513 1779 57569
rect 1865 57513 1921 57569
rect 2007 57513 2063 57569
rect 2149 57513 2205 57569
rect 2291 57513 2347 57569
rect 2433 57513 2489 57569
rect 2575 57513 2631 57569
rect 2717 57513 2773 57569
rect 2859 57513 2915 57569
rect 3001 57513 3057 57569
rect 3143 57513 3199 57569
rect 3285 57513 3341 57569
rect 3427 57513 3483 57569
rect 3569 57513 3625 57569
rect 3711 57513 3767 57569
rect 3853 57513 3909 57569
rect 3995 57513 4051 57569
rect 4137 57513 4193 57569
rect 4279 57513 4335 57569
rect 4421 57513 4477 57569
rect 4563 57513 4619 57569
rect 4705 57513 4761 57569
rect 4847 57513 4903 57569
rect 4989 57513 5045 57569
rect 5131 57513 5187 57569
rect 5273 57513 5329 57569
rect 5415 57513 5471 57569
rect 5557 57513 5613 57569
rect 5699 57513 5755 57569
rect 5841 57513 5897 57569
rect 5983 57513 6039 57569
rect 6125 57513 6181 57569
rect 6267 57513 6323 57569
rect 6409 57513 6465 57569
rect 6551 57513 6607 57569
rect 6693 57513 6749 57569
rect 6835 57513 6891 57569
rect 6977 57513 7033 57569
rect 7119 57513 7175 57569
rect 7261 57513 7317 57569
rect 7403 57513 7459 57569
rect 7545 57513 7601 57569
rect 7687 57513 7743 57569
rect 7829 57513 7885 57569
rect 7971 57513 8027 57569
rect 8113 57513 8169 57569
rect 8255 57513 8311 57569
rect 8397 57513 8453 57569
rect 8539 57513 8595 57569
rect 8681 57513 8737 57569
rect 8823 57513 8879 57569
rect 8965 57513 9021 57569
rect 9107 57513 9163 57569
rect 9249 57513 9305 57569
rect 9391 57513 9447 57569
rect 9533 57513 9589 57569
rect 9675 57513 9731 57569
rect 9817 57513 9873 57569
rect 9959 57513 10015 57569
rect 10101 57513 10157 57569
rect 10243 57513 10299 57569
rect 10385 57513 10441 57569
rect 10527 57513 10583 57569
rect 10669 57513 10725 57569
rect 10811 57513 10867 57569
rect 10953 57513 11009 57569
rect 11095 57513 11151 57569
rect 11237 57513 11293 57569
rect 11379 57513 11435 57569
rect 11521 57513 11577 57569
rect 11663 57513 11719 57569
rect 11805 57513 11861 57569
rect 11947 57513 12003 57569
rect 12089 57513 12145 57569
rect 12231 57513 12287 57569
rect 12373 57513 12429 57569
rect 12515 57513 12571 57569
rect 12657 57513 12713 57569
rect 12799 57513 12855 57569
rect 12941 57513 12997 57569
rect 13083 57513 13139 57569
rect 13225 57513 13281 57569
rect 13367 57513 13423 57569
rect 13509 57513 13565 57569
rect 13651 57513 13707 57569
rect 13793 57513 13849 57569
rect 13935 57513 13991 57569
rect 14077 57513 14133 57569
rect 14219 57513 14275 57569
rect 14361 57513 14417 57569
rect 14503 57513 14559 57569
rect 14645 57513 14701 57569
rect 14787 57513 14843 57569
rect 161 57371 217 57427
rect 303 57371 359 57427
rect 445 57371 501 57427
rect 587 57371 643 57427
rect 729 57371 785 57427
rect 871 57371 927 57427
rect 1013 57371 1069 57427
rect 1155 57371 1211 57427
rect 1297 57371 1353 57427
rect 1439 57371 1495 57427
rect 1581 57371 1637 57427
rect 1723 57371 1779 57427
rect 1865 57371 1921 57427
rect 2007 57371 2063 57427
rect 2149 57371 2205 57427
rect 2291 57371 2347 57427
rect 2433 57371 2489 57427
rect 2575 57371 2631 57427
rect 2717 57371 2773 57427
rect 2859 57371 2915 57427
rect 3001 57371 3057 57427
rect 3143 57371 3199 57427
rect 3285 57371 3341 57427
rect 3427 57371 3483 57427
rect 3569 57371 3625 57427
rect 3711 57371 3767 57427
rect 3853 57371 3909 57427
rect 3995 57371 4051 57427
rect 4137 57371 4193 57427
rect 4279 57371 4335 57427
rect 4421 57371 4477 57427
rect 4563 57371 4619 57427
rect 4705 57371 4761 57427
rect 4847 57371 4903 57427
rect 4989 57371 5045 57427
rect 5131 57371 5187 57427
rect 5273 57371 5329 57427
rect 5415 57371 5471 57427
rect 5557 57371 5613 57427
rect 5699 57371 5755 57427
rect 5841 57371 5897 57427
rect 5983 57371 6039 57427
rect 6125 57371 6181 57427
rect 6267 57371 6323 57427
rect 6409 57371 6465 57427
rect 6551 57371 6607 57427
rect 6693 57371 6749 57427
rect 6835 57371 6891 57427
rect 6977 57371 7033 57427
rect 7119 57371 7175 57427
rect 7261 57371 7317 57427
rect 7403 57371 7459 57427
rect 7545 57371 7601 57427
rect 7687 57371 7743 57427
rect 7829 57371 7885 57427
rect 7971 57371 8027 57427
rect 8113 57371 8169 57427
rect 8255 57371 8311 57427
rect 8397 57371 8453 57427
rect 8539 57371 8595 57427
rect 8681 57371 8737 57427
rect 8823 57371 8879 57427
rect 8965 57371 9021 57427
rect 9107 57371 9163 57427
rect 9249 57371 9305 57427
rect 9391 57371 9447 57427
rect 9533 57371 9589 57427
rect 9675 57371 9731 57427
rect 9817 57371 9873 57427
rect 9959 57371 10015 57427
rect 10101 57371 10157 57427
rect 10243 57371 10299 57427
rect 10385 57371 10441 57427
rect 10527 57371 10583 57427
rect 10669 57371 10725 57427
rect 10811 57371 10867 57427
rect 10953 57371 11009 57427
rect 11095 57371 11151 57427
rect 11237 57371 11293 57427
rect 11379 57371 11435 57427
rect 11521 57371 11577 57427
rect 11663 57371 11719 57427
rect 11805 57371 11861 57427
rect 11947 57371 12003 57427
rect 12089 57371 12145 57427
rect 12231 57371 12287 57427
rect 12373 57371 12429 57427
rect 12515 57371 12571 57427
rect 12657 57371 12713 57427
rect 12799 57371 12855 57427
rect 12941 57371 12997 57427
rect 13083 57371 13139 57427
rect 13225 57371 13281 57427
rect 13367 57371 13423 57427
rect 13509 57371 13565 57427
rect 13651 57371 13707 57427
rect 13793 57371 13849 57427
rect 13935 57371 13991 57427
rect 14077 57371 14133 57427
rect 14219 57371 14275 57427
rect 14361 57371 14417 57427
rect 14503 57371 14559 57427
rect 14645 57371 14701 57427
rect 14787 57371 14843 57427
rect 161 57229 217 57285
rect 303 57229 359 57285
rect 445 57229 501 57285
rect 587 57229 643 57285
rect 729 57229 785 57285
rect 871 57229 927 57285
rect 1013 57229 1069 57285
rect 1155 57229 1211 57285
rect 1297 57229 1353 57285
rect 1439 57229 1495 57285
rect 1581 57229 1637 57285
rect 1723 57229 1779 57285
rect 1865 57229 1921 57285
rect 2007 57229 2063 57285
rect 2149 57229 2205 57285
rect 2291 57229 2347 57285
rect 2433 57229 2489 57285
rect 2575 57229 2631 57285
rect 2717 57229 2773 57285
rect 2859 57229 2915 57285
rect 3001 57229 3057 57285
rect 3143 57229 3199 57285
rect 3285 57229 3341 57285
rect 3427 57229 3483 57285
rect 3569 57229 3625 57285
rect 3711 57229 3767 57285
rect 3853 57229 3909 57285
rect 3995 57229 4051 57285
rect 4137 57229 4193 57285
rect 4279 57229 4335 57285
rect 4421 57229 4477 57285
rect 4563 57229 4619 57285
rect 4705 57229 4761 57285
rect 4847 57229 4903 57285
rect 4989 57229 5045 57285
rect 5131 57229 5187 57285
rect 5273 57229 5329 57285
rect 5415 57229 5471 57285
rect 5557 57229 5613 57285
rect 5699 57229 5755 57285
rect 5841 57229 5897 57285
rect 5983 57229 6039 57285
rect 6125 57229 6181 57285
rect 6267 57229 6323 57285
rect 6409 57229 6465 57285
rect 6551 57229 6607 57285
rect 6693 57229 6749 57285
rect 6835 57229 6891 57285
rect 6977 57229 7033 57285
rect 7119 57229 7175 57285
rect 7261 57229 7317 57285
rect 7403 57229 7459 57285
rect 7545 57229 7601 57285
rect 7687 57229 7743 57285
rect 7829 57229 7885 57285
rect 7971 57229 8027 57285
rect 8113 57229 8169 57285
rect 8255 57229 8311 57285
rect 8397 57229 8453 57285
rect 8539 57229 8595 57285
rect 8681 57229 8737 57285
rect 8823 57229 8879 57285
rect 8965 57229 9021 57285
rect 9107 57229 9163 57285
rect 9249 57229 9305 57285
rect 9391 57229 9447 57285
rect 9533 57229 9589 57285
rect 9675 57229 9731 57285
rect 9817 57229 9873 57285
rect 9959 57229 10015 57285
rect 10101 57229 10157 57285
rect 10243 57229 10299 57285
rect 10385 57229 10441 57285
rect 10527 57229 10583 57285
rect 10669 57229 10725 57285
rect 10811 57229 10867 57285
rect 10953 57229 11009 57285
rect 11095 57229 11151 57285
rect 11237 57229 11293 57285
rect 11379 57229 11435 57285
rect 11521 57229 11577 57285
rect 11663 57229 11719 57285
rect 11805 57229 11861 57285
rect 11947 57229 12003 57285
rect 12089 57229 12145 57285
rect 12231 57229 12287 57285
rect 12373 57229 12429 57285
rect 12515 57229 12571 57285
rect 12657 57229 12713 57285
rect 12799 57229 12855 57285
rect 12941 57229 12997 57285
rect 13083 57229 13139 57285
rect 13225 57229 13281 57285
rect 13367 57229 13423 57285
rect 13509 57229 13565 57285
rect 13651 57229 13707 57285
rect 13793 57229 13849 57285
rect 13935 57229 13991 57285
rect 14077 57229 14133 57285
rect 14219 57229 14275 57285
rect 14361 57229 14417 57285
rect 14503 57229 14559 57285
rect 14645 57229 14701 57285
rect 14787 57229 14843 57285
rect 161 56915 217 56971
rect 303 56915 359 56971
rect 445 56915 501 56971
rect 587 56915 643 56971
rect 729 56915 785 56971
rect 871 56915 927 56971
rect 1013 56915 1069 56971
rect 1155 56915 1211 56971
rect 1297 56915 1353 56971
rect 1439 56915 1495 56971
rect 1581 56915 1637 56971
rect 1723 56915 1779 56971
rect 1865 56915 1921 56971
rect 2007 56915 2063 56971
rect 2149 56915 2205 56971
rect 2291 56915 2347 56971
rect 2433 56915 2489 56971
rect 2575 56915 2631 56971
rect 2717 56915 2773 56971
rect 2859 56915 2915 56971
rect 3001 56915 3057 56971
rect 3143 56915 3199 56971
rect 3285 56915 3341 56971
rect 3427 56915 3483 56971
rect 3569 56915 3625 56971
rect 3711 56915 3767 56971
rect 3853 56915 3909 56971
rect 3995 56915 4051 56971
rect 4137 56915 4193 56971
rect 4279 56915 4335 56971
rect 4421 56915 4477 56971
rect 4563 56915 4619 56971
rect 4705 56915 4761 56971
rect 4847 56915 4903 56971
rect 4989 56915 5045 56971
rect 5131 56915 5187 56971
rect 5273 56915 5329 56971
rect 5415 56915 5471 56971
rect 5557 56915 5613 56971
rect 5699 56915 5755 56971
rect 5841 56915 5897 56971
rect 5983 56915 6039 56971
rect 6125 56915 6181 56971
rect 6267 56915 6323 56971
rect 6409 56915 6465 56971
rect 6551 56915 6607 56971
rect 6693 56915 6749 56971
rect 6835 56915 6891 56971
rect 6977 56915 7033 56971
rect 7119 56915 7175 56971
rect 7261 56915 7317 56971
rect 7403 56915 7459 56971
rect 7545 56915 7601 56971
rect 7687 56915 7743 56971
rect 7829 56915 7885 56971
rect 7971 56915 8027 56971
rect 8113 56915 8169 56971
rect 8255 56915 8311 56971
rect 8397 56915 8453 56971
rect 8539 56915 8595 56971
rect 8681 56915 8737 56971
rect 8823 56915 8879 56971
rect 8965 56915 9021 56971
rect 9107 56915 9163 56971
rect 9249 56915 9305 56971
rect 9391 56915 9447 56971
rect 9533 56915 9589 56971
rect 9675 56915 9731 56971
rect 9817 56915 9873 56971
rect 9959 56915 10015 56971
rect 10101 56915 10157 56971
rect 10243 56915 10299 56971
rect 10385 56915 10441 56971
rect 10527 56915 10583 56971
rect 10669 56915 10725 56971
rect 10811 56915 10867 56971
rect 10953 56915 11009 56971
rect 11095 56915 11151 56971
rect 11237 56915 11293 56971
rect 11379 56915 11435 56971
rect 11521 56915 11577 56971
rect 11663 56915 11719 56971
rect 11805 56915 11861 56971
rect 11947 56915 12003 56971
rect 12089 56915 12145 56971
rect 12231 56915 12287 56971
rect 12373 56915 12429 56971
rect 12515 56915 12571 56971
rect 12657 56915 12713 56971
rect 12799 56915 12855 56971
rect 12941 56915 12997 56971
rect 13083 56915 13139 56971
rect 13225 56915 13281 56971
rect 13367 56915 13423 56971
rect 13509 56915 13565 56971
rect 13651 56915 13707 56971
rect 13793 56915 13849 56971
rect 13935 56915 13991 56971
rect 14077 56915 14133 56971
rect 14219 56915 14275 56971
rect 14361 56915 14417 56971
rect 14503 56915 14559 56971
rect 14645 56915 14701 56971
rect 14787 56915 14843 56971
rect 161 56773 217 56829
rect 303 56773 359 56829
rect 445 56773 501 56829
rect 587 56773 643 56829
rect 729 56773 785 56829
rect 871 56773 927 56829
rect 1013 56773 1069 56829
rect 1155 56773 1211 56829
rect 1297 56773 1353 56829
rect 1439 56773 1495 56829
rect 1581 56773 1637 56829
rect 1723 56773 1779 56829
rect 1865 56773 1921 56829
rect 2007 56773 2063 56829
rect 2149 56773 2205 56829
rect 2291 56773 2347 56829
rect 2433 56773 2489 56829
rect 2575 56773 2631 56829
rect 2717 56773 2773 56829
rect 2859 56773 2915 56829
rect 3001 56773 3057 56829
rect 3143 56773 3199 56829
rect 3285 56773 3341 56829
rect 3427 56773 3483 56829
rect 3569 56773 3625 56829
rect 3711 56773 3767 56829
rect 3853 56773 3909 56829
rect 3995 56773 4051 56829
rect 4137 56773 4193 56829
rect 4279 56773 4335 56829
rect 4421 56773 4477 56829
rect 4563 56773 4619 56829
rect 4705 56773 4761 56829
rect 4847 56773 4903 56829
rect 4989 56773 5045 56829
rect 5131 56773 5187 56829
rect 5273 56773 5329 56829
rect 5415 56773 5471 56829
rect 5557 56773 5613 56829
rect 5699 56773 5755 56829
rect 5841 56773 5897 56829
rect 5983 56773 6039 56829
rect 6125 56773 6181 56829
rect 6267 56773 6323 56829
rect 6409 56773 6465 56829
rect 6551 56773 6607 56829
rect 6693 56773 6749 56829
rect 6835 56773 6891 56829
rect 6977 56773 7033 56829
rect 7119 56773 7175 56829
rect 7261 56773 7317 56829
rect 7403 56773 7459 56829
rect 7545 56773 7601 56829
rect 7687 56773 7743 56829
rect 7829 56773 7885 56829
rect 7971 56773 8027 56829
rect 8113 56773 8169 56829
rect 8255 56773 8311 56829
rect 8397 56773 8453 56829
rect 8539 56773 8595 56829
rect 8681 56773 8737 56829
rect 8823 56773 8879 56829
rect 8965 56773 9021 56829
rect 9107 56773 9163 56829
rect 9249 56773 9305 56829
rect 9391 56773 9447 56829
rect 9533 56773 9589 56829
rect 9675 56773 9731 56829
rect 9817 56773 9873 56829
rect 9959 56773 10015 56829
rect 10101 56773 10157 56829
rect 10243 56773 10299 56829
rect 10385 56773 10441 56829
rect 10527 56773 10583 56829
rect 10669 56773 10725 56829
rect 10811 56773 10867 56829
rect 10953 56773 11009 56829
rect 11095 56773 11151 56829
rect 11237 56773 11293 56829
rect 11379 56773 11435 56829
rect 11521 56773 11577 56829
rect 11663 56773 11719 56829
rect 11805 56773 11861 56829
rect 11947 56773 12003 56829
rect 12089 56773 12145 56829
rect 12231 56773 12287 56829
rect 12373 56773 12429 56829
rect 12515 56773 12571 56829
rect 12657 56773 12713 56829
rect 12799 56773 12855 56829
rect 12941 56773 12997 56829
rect 13083 56773 13139 56829
rect 13225 56773 13281 56829
rect 13367 56773 13423 56829
rect 13509 56773 13565 56829
rect 13651 56773 13707 56829
rect 13793 56773 13849 56829
rect 13935 56773 13991 56829
rect 14077 56773 14133 56829
rect 14219 56773 14275 56829
rect 14361 56773 14417 56829
rect 14503 56773 14559 56829
rect 14645 56773 14701 56829
rect 14787 56773 14843 56829
rect 161 56631 217 56687
rect 303 56631 359 56687
rect 445 56631 501 56687
rect 587 56631 643 56687
rect 729 56631 785 56687
rect 871 56631 927 56687
rect 1013 56631 1069 56687
rect 1155 56631 1211 56687
rect 1297 56631 1353 56687
rect 1439 56631 1495 56687
rect 1581 56631 1637 56687
rect 1723 56631 1779 56687
rect 1865 56631 1921 56687
rect 2007 56631 2063 56687
rect 2149 56631 2205 56687
rect 2291 56631 2347 56687
rect 2433 56631 2489 56687
rect 2575 56631 2631 56687
rect 2717 56631 2773 56687
rect 2859 56631 2915 56687
rect 3001 56631 3057 56687
rect 3143 56631 3199 56687
rect 3285 56631 3341 56687
rect 3427 56631 3483 56687
rect 3569 56631 3625 56687
rect 3711 56631 3767 56687
rect 3853 56631 3909 56687
rect 3995 56631 4051 56687
rect 4137 56631 4193 56687
rect 4279 56631 4335 56687
rect 4421 56631 4477 56687
rect 4563 56631 4619 56687
rect 4705 56631 4761 56687
rect 4847 56631 4903 56687
rect 4989 56631 5045 56687
rect 5131 56631 5187 56687
rect 5273 56631 5329 56687
rect 5415 56631 5471 56687
rect 5557 56631 5613 56687
rect 5699 56631 5755 56687
rect 5841 56631 5897 56687
rect 5983 56631 6039 56687
rect 6125 56631 6181 56687
rect 6267 56631 6323 56687
rect 6409 56631 6465 56687
rect 6551 56631 6607 56687
rect 6693 56631 6749 56687
rect 6835 56631 6891 56687
rect 6977 56631 7033 56687
rect 7119 56631 7175 56687
rect 7261 56631 7317 56687
rect 7403 56631 7459 56687
rect 7545 56631 7601 56687
rect 7687 56631 7743 56687
rect 7829 56631 7885 56687
rect 7971 56631 8027 56687
rect 8113 56631 8169 56687
rect 8255 56631 8311 56687
rect 8397 56631 8453 56687
rect 8539 56631 8595 56687
rect 8681 56631 8737 56687
rect 8823 56631 8879 56687
rect 8965 56631 9021 56687
rect 9107 56631 9163 56687
rect 9249 56631 9305 56687
rect 9391 56631 9447 56687
rect 9533 56631 9589 56687
rect 9675 56631 9731 56687
rect 9817 56631 9873 56687
rect 9959 56631 10015 56687
rect 10101 56631 10157 56687
rect 10243 56631 10299 56687
rect 10385 56631 10441 56687
rect 10527 56631 10583 56687
rect 10669 56631 10725 56687
rect 10811 56631 10867 56687
rect 10953 56631 11009 56687
rect 11095 56631 11151 56687
rect 11237 56631 11293 56687
rect 11379 56631 11435 56687
rect 11521 56631 11577 56687
rect 11663 56631 11719 56687
rect 11805 56631 11861 56687
rect 11947 56631 12003 56687
rect 12089 56631 12145 56687
rect 12231 56631 12287 56687
rect 12373 56631 12429 56687
rect 12515 56631 12571 56687
rect 12657 56631 12713 56687
rect 12799 56631 12855 56687
rect 12941 56631 12997 56687
rect 13083 56631 13139 56687
rect 13225 56631 13281 56687
rect 13367 56631 13423 56687
rect 13509 56631 13565 56687
rect 13651 56631 13707 56687
rect 13793 56631 13849 56687
rect 13935 56631 13991 56687
rect 14077 56631 14133 56687
rect 14219 56631 14275 56687
rect 14361 56631 14417 56687
rect 14503 56631 14559 56687
rect 14645 56631 14701 56687
rect 14787 56631 14843 56687
rect 161 56489 217 56545
rect 303 56489 359 56545
rect 445 56489 501 56545
rect 587 56489 643 56545
rect 729 56489 785 56545
rect 871 56489 927 56545
rect 1013 56489 1069 56545
rect 1155 56489 1211 56545
rect 1297 56489 1353 56545
rect 1439 56489 1495 56545
rect 1581 56489 1637 56545
rect 1723 56489 1779 56545
rect 1865 56489 1921 56545
rect 2007 56489 2063 56545
rect 2149 56489 2205 56545
rect 2291 56489 2347 56545
rect 2433 56489 2489 56545
rect 2575 56489 2631 56545
rect 2717 56489 2773 56545
rect 2859 56489 2915 56545
rect 3001 56489 3057 56545
rect 3143 56489 3199 56545
rect 3285 56489 3341 56545
rect 3427 56489 3483 56545
rect 3569 56489 3625 56545
rect 3711 56489 3767 56545
rect 3853 56489 3909 56545
rect 3995 56489 4051 56545
rect 4137 56489 4193 56545
rect 4279 56489 4335 56545
rect 4421 56489 4477 56545
rect 4563 56489 4619 56545
rect 4705 56489 4761 56545
rect 4847 56489 4903 56545
rect 4989 56489 5045 56545
rect 5131 56489 5187 56545
rect 5273 56489 5329 56545
rect 5415 56489 5471 56545
rect 5557 56489 5613 56545
rect 5699 56489 5755 56545
rect 5841 56489 5897 56545
rect 5983 56489 6039 56545
rect 6125 56489 6181 56545
rect 6267 56489 6323 56545
rect 6409 56489 6465 56545
rect 6551 56489 6607 56545
rect 6693 56489 6749 56545
rect 6835 56489 6891 56545
rect 6977 56489 7033 56545
rect 7119 56489 7175 56545
rect 7261 56489 7317 56545
rect 7403 56489 7459 56545
rect 7545 56489 7601 56545
rect 7687 56489 7743 56545
rect 7829 56489 7885 56545
rect 7971 56489 8027 56545
rect 8113 56489 8169 56545
rect 8255 56489 8311 56545
rect 8397 56489 8453 56545
rect 8539 56489 8595 56545
rect 8681 56489 8737 56545
rect 8823 56489 8879 56545
rect 8965 56489 9021 56545
rect 9107 56489 9163 56545
rect 9249 56489 9305 56545
rect 9391 56489 9447 56545
rect 9533 56489 9589 56545
rect 9675 56489 9731 56545
rect 9817 56489 9873 56545
rect 9959 56489 10015 56545
rect 10101 56489 10157 56545
rect 10243 56489 10299 56545
rect 10385 56489 10441 56545
rect 10527 56489 10583 56545
rect 10669 56489 10725 56545
rect 10811 56489 10867 56545
rect 10953 56489 11009 56545
rect 11095 56489 11151 56545
rect 11237 56489 11293 56545
rect 11379 56489 11435 56545
rect 11521 56489 11577 56545
rect 11663 56489 11719 56545
rect 11805 56489 11861 56545
rect 11947 56489 12003 56545
rect 12089 56489 12145 56545
rect 12231 56489 12287 56545
rect 12373 56489 12429 56545
rect 12515 56489 12571 56545
rect 12657 56489 12713 56545
rect 12799 56489 12855 56545
rect 12941 56489 12997 56545
rect 13083 56489 13139 56545
rect 13225 56489 13281 56545
rect 13367 56489 13423 56545
rect 13509 56489 13565 56545
rect 13651 56489 13707 56545
rect 13793 56489 13849 56545
rect 13935 56489 13991 56545
rect 14077 56489 14133 56545
rect 14219 56489 14275 56545
rect 14361 56489 14417 56545
rect 14503 56489 14559 56545
rect 14645 56489 14701 56545
rect 14787 56489 14843 56545
rect 161 56347 217 56403
rect 303 56347 359 56403
rect 445 56347 501 56403
rect 587 56347 643 56403
rect 729 56347 785 56403
rect 871 56347 927 56403
rect 1013 56347 1069 56403
rect 1155 56347 1211 56403
rect 1297 56347 1353 56403
rect 1439 56347 1495 56403
rect 1581 56347 1637 56403
rect 1723 56347 1779 56403
rect 1865 56347 1921 56403
rect 2007 56347 2063 56403
rect 2149 56347 2205 56403
rect 2291 56347 2347 56403
rect 2433 56347 2489 56403
rect 2575 56347 2631 56403
rect 2717 56347 2773 56403
rect 2859 56347 2915 56403
rect 3001 56347 3057 56403
rect 3143 56347 3199 56403
rect 3285 56347 3341 56403
rect 3427 56347 3483 56403
rect 3569 56347 3625 56403
rect 3711 56347 3767 56403
rect 3853 56347 3909 56403
rect 3995 56347 4051 56403
rect 4137 56347 4193 56403
rect 4279 56347 4335 56403
rect 4421 56347 4477 56403
rect 4563 56347 4619 56403
rect 4705 56347 4761 56403
rect 4847 56347 4903 56403
rect 4989 56347 5045 56403
rect 5131 56347 5187 56403
rect 5273 56347 5329 56403
rect 5415 56347 5471 56403
rect 5557 56347 5613 56403
rect 5699 56347 5755 56403
rect 5841 56347 5897 56403
rect 5983 56347 6039 56403
rect 6125 56347 6181 56403
rect 6267 56347 6323 56403
rect 6409 56347 6465 56403
rect 6551 56347 6607 56403
rect 6693 56347 6749 56403
rect 6835 56347 6891 56403
rect 6977 56347 7033 56403
rect 7119 56347 7175 56403
rect 7261 56347 7317 56403
rect 7403 56347 7459 56403
rect 7545 56347 7601 56403
rect 7687 56347 7743 56403
rect 7829 56347 7885 56403
rect 7971 56347 8027 56403
rect 8113 56347 8169 56403
rect 8255 56347 8311 56403
rect 8397 56347 8453 56403
rect 8539 56347 8595 56403
rect 8681 56347 8737 56403
rect 8823 56347 8879 56403
rect 8965 56347 9021 56403
rect 9107 56347 9163 56403
rect 9249 56347 9305 56403
rect 9391 56347 9447 56403
rect 9533 56347 9589 56403
rect 9675 56347 9731 56403
rect 9817 56347 9873 56403
rect 9959 56347 10015 56403
rect 10101 56347 10157 56403
rect 10243 56347 10299 56403
rect 10385 56347 10441 56403
rect 10527 56347 10583 56403
rect 10669 56347 10725 56403
rect 10811 56347 10867 56403
rect 10953 56347 11009 56403
rect 11095 56347 11151 56403
rect 11237 56347 11293 56403
rect 11379 56347 11435 56403
rect 11521 56347 11577 56403
rect 11663 56347 11719 56403
rect 11805 56347 11861 56403
rect 11947 56347 12003 56403
rect 12089 56347 12145 56403
rect 12231 56347 12287 56403
rect 12373 56347 12429 56403
rect 12515 56347 12571 56403
rect 12657 56347 12713 56403
rect 12799 56347 12855 56403
rect 12941 56347 12997 56403
rect 13083 56347 13139 56403
rect 13225 56347 13281 56403
rect 13367 56347 13423 56403
rect 13509 56347 13565 56403
rect 13651 56347 13707 56403
rect 13793 56347 13849 56403
rect 13935 56347 13991 56403
rect 14077 56347 14133 56403
rect 14219 56347 14275 56403
rect 14361 56347 14417 56403
rect 14503 56347 14559 56403
rect 14645 56347 14701 56403
rect 14787 56347 14843 56403
rect 161 56205 217 56261
rect 303 56205 359 56261
rect 445 56205 501 56261
rect 587 56205 643 56261
rect 729 56205 785 56261
rect 871 56205 927 56261
rect 1013 56205 1069 56261
rect 1155 56205 1211 56261
rect 1297 56205 1353 56261
rect 1439 56205 1495 56261
rect 1581 56205 1637 56261
rect 1723 56205 1779 56261
rect 1865 56205 1921 56261
rect 2007 56205 2063 56261
rect 2149 56205 2205 56261
rect 2291 56205 2347 56261
rect 2433 56205 2489 56261
rect 2575 56205 2631 56261
rect 2717 56205 2773 56261
rect 2859 56205 2915 56261
rect 3001 56205 3057 56261
rect 3143 56205 3199 56261
rect 3285 56205 3341 56261
rect 3427 56205 3483 56261
rect 3569 56205 3625 56261
rect 3711 56205 3767 56261
rect 3853 56205 3909 56261
rect 3995 56205 4051 56261
rect 4137 56205 4193 56261
rect 4279 56205 4335 56261
rect 4421 56205 4477 56261
rect 4563 56205 4619 56261
rect 4705 56205 4761 56261
rect 4847 56205 4903 56261
rect 4989 56205 5045 56261
rect 5131 56205 5187 56261
rect 5273 56205 5329 56261
rect 5415 56205 5471 56261
rect 5557 56205 5613 56261
rect 5699 56205 5755 56261
rect 5841 56205 5897 56261
rect 5983 56205 6039 56261
rect 6125 56205 6181 56261
rect 6267 56205 6323 56261
rect 6409 56205 6465 56261
rect 6551 56205 6607 56261
rect 6693 56205 6749 56261
rect 6835 56205 6891 56261
rect 6977 56205 7033 56261
rect 7119 56205 7175 56261
rect 7261 56205 7317 56261
rect 7403 56205 7459 56261
rect 7545 56205 7601 56261
rect 7687 56205 7743 56261
rect 7829 56205 7885 56261
rect 7971 56205 8027 56261
rect 8113 56205 8169 56261
rect 8255 56205 8311 56261
rect 8397 56205 8453 56261
rect 8539 56205 8595 56261
rect 8681 56205 8737 56261
rect 8823 56205 8879 56261
rect 8965 56205 9021 56261
rect 9107 56205 9163 56261
rect 9249 56205 9305 56261
rect 9391 56205 9447 56261
rect 9533 56205 9589 56261
rect 9675 56205 9731 56261
rect 9817 56205 9873 56261
rect 9959 56205 10015 56261
rect 10101 56205 10157 56261
rect 10243 56205 10299 56261
rect 10385 56205 10441 56261
rect 10527 56205 10583 56261
rect 10669 56205 10725 56261
rect 10811 56205 10867 56261
rect 10953 56205 11009 56261
rect 11095 56205 11151 56261
rect 11237 56205 11293 56261
rect 11379 56205 11435 56261
rect 11521 56205 11577 56261
rect 11663 56205 11719 56261
rect 11805 56205 11861 56261
rect 11947 56205 12003 56261
rect 12089 56205 12145 56261
rect 12231 56205 12287 56261
rect 12373 56205 12429 56261
rect 12515 56205 12571 56261
rect 12657 56205 12713 56261
rect 12799 56205 12855 56261
rect 12941 56205 12997 56261
rect 13083 56205 13139 56261
rect 13225 56205 13281 56261
rect 13367 56205 13423 56261
rect 13509 56205 13565 56261
rect 13651 56205 13707 56261
rect 13793 56205 13849 56261
rect 13935 56205 13991 56261
rect 14077 56205 14133 56261
rect 14219 56205 14275 56261
rect 14361 56205 14417 56261
rect 14503 56205 14559 56261
rect 14645 56205 14701 56261
rect 14787 56205 14843 56261
rect 161 56063 217 56119
rect 303 56063 359 56119
rect 445 56063 501 56119
rect 587 56063 643 56119
rect 729 56063 785 56119
rect 871 56063 927 56119
rect 1013 56063 1069 56119
rect 1155 56063 1211 56119
rect 1297 56063 1353 56119
rect 1439 56063 1495 56119
rect 1581 56063 1637 56119
rect 1723 56063 1779 56119
rect 1865 56063 1921 56119
rect 2007 56063 2063 56119
rect 2149 56063 2205 56119
rect 2291 56063 2347 56119
rect 2433 56063 2489 56119
rect 2575 56063 2631 56119
rect 2717 56063 2773 56119
rect 2859 56063 2915 56119
rect 3001 56063 3057 56119
rect 3143 56063 3199 56119
rect 3285 56063 3341 56119
rect 3427 56063 3483 56119
rect 3569 56063 3625 56119
rect 3711 56063 3767 56119
rect 3853 56063 3909 56119
rect 3995 56063 4051 56119
rect 4137 56063 4193 56119
rect 4279 56063 4335 56119
rect 4421 56063 4477 56119
rect 4563 56063 4619 56119
rect 4705 56063 4761 56119
rect 4847 56063 4903 56119
rect 4989 56063 5045 56119
rect 5131 56063 5187 56119
rect 5273 56063 5329 56119
rect 5415 56063 5471 56119
rect 5557 56063 5613 56119
rect 5699 56063 5755 56119
rect 5841 56063 5897 56119
rect 5983 56063 6039 56119
rect 6125 56063 6181 56119
rect 6267 56063 6323 56119
rect 6409 56063 6465 56119
rect 6551 56063 6607 56119
rect 6693 56063 6749 56119
rect 6835 56063 6891 56119
rect 6977 56063 7033 56119
rect 7119 56063 7175 56119
rect 7261 56063 7317 56119
rect 7403 56063 7459 56119
rect 7545 56063 7601 56119
rect 7687 56063 7743 56119
rect 7829 56063 7885 56119
rect 7971 56063 8027 56119
rect 8113 56063 8169 56119
rect 8255 56063 8311 56119
rect 8397 56063 8453 56119
rect 8539 56063 8595 56119
rect 8681 56063 8737 56119
rect 8823 56063 8879 56119
rect 8965 56063 9021 56119
rect 9107 56063 9163 56119
rect 9249 56063 9305 56119
rect 9391 56063 9447 56119
rect 9533 56063 9589 56119
rect 9675 56063 9731 56119
rect 9817 56063 9873 56119
rect 9959 56063 10015 56119
rect 10101 56063 10157 56119
rect 10243 56063 10299 56119
rect 10385 56063 10441 56119
rect 10527 56063 10583 56119
rect 10669 56063 10725 56119
rect 10811 56063 10867 56119
rect 10953 56063 11009 56119
rect 11095 56063 11151 56119
rect 11237 56063 11293 56119
rect 11379 56063 11435 56119
rect 11521 56063 11577 56119
rect 11663 56063 11719 56119
rect 11805 56063 11861 56119
rect 11947 56063 12003 56119
rect 12089 56063 12145 56119
rect 12231 56063 12287 56119
rect 12373 56063 12429 56119
rect 12515 56063 12571 56119
rect 12657 56063 12713 56119
rect 12799 56063 12855 56119
rect 12941 56063 12997 56119
rect 13083 56063 13139 56119
rect 13225 56063 13281 56119
rect 13367 56063 13423 56119
rect 13509 56063 13565 56119
rect 13651 56063 13707 56119
rect 13793 56063 13849 56119
rect 13935 56063 13991 56119
rect 14077 56063 14133 56119
rect 14219 56063 14275 56119
rect 14361 56063 14417 56119
rect 14503 56063 14559 56119
rect 14645 56063 14701 56119
rect 14787 56063 14843 56119
rect 161 55921 217 55977
rect 303 55921 359 55977
rect 445 55921 501 55977
rect 587 55921 643 55977
rect 729 55921 785 55977
rect 871 55921 927 55977
rect 1013 55921 1069 55977
rect 1155 55921 1211 55977
rect 1297 55921 1353 55977
rect 1439 55921 1495 55977
rect 1581 55921 1637 55977
rect 1723 55921 1779 55977
rect 1865 55921 1921 55977
rect 2007 55921 2063 55977
rect 2149 55921 2205 55977
rect 2291 55921 2347 55977
rect 2433 55921 2489 55977
rect 2575 55921 2631 55977
rect 2717 55921 2773 55977
rect 2859 55921 2915 55977
rect 3001 55921 3057 55977
rect 3143 55921 3199 55977
rect 3285 55921 3341 55977
rect 3427 55921 3483 55977
rect 3569 55921 3625 55977
rect 3711 55921 3767 55977
rect 3853 55921 3909 55977
rect 3995 55921 4051 55977
rect 4137 55921 4193 55977
rect 4279 55921 4335 55977
rect 4421 55921 4477 55977
rect 4563 55921 4619 55977
rect 4705 55921 4761 55977
rect 4847 55921 4903 55977
rect 4989 55921 5045 55977
rect 5131 55921 5187 55977
rect 5273 55921 5329 55977
rect 5415 55921 5471 55977
rect 5557 55921 5613 55977
rect 5699 55921 5755 55977
rect 5841 55921 5897 55977
rect 5983 55921 6039 55977
rect 6125 55921 6181 55977
rect 6267 55921 6323 55977
rect 6409 55921 6465 55977
rect 6551 55921 6607 55977
rect 6693 55921 6749 55977
rect 6835 55921 6891 55977
rect 6977 55921 7033 55977
rect 7119 55921 7175 55977
rect 7261 55921 7317 55977
rect 7403 55921 7459 55977
rect 7545 55921 7601 55977
rect 7687 55921 7743 55977
rect 7829 55921 7885 55977
rect 7971 55921 8027 55977
rect 8113 55921 8169 55977
rect 8255 55921 8311 55977
rect 8397 55921 8453 55977
rect 8539 55921 8595 55977
rect 8681 55921 8737 55977
rect 8823 55921 8879 55977
rect 8965 55921 9021 55977
rect 9107 55921 9163 55977
rect 9249 55921 9305 55977
rect 9391 55921 9447 55977
rect 9533 55921 9589 55977
rect 9675 55921 9731 55977
rect 9817 55921 9873 55977
rect 9959 55921 10015 55977
rect 10101 55921 10157 55977
rect 10243 55921 10299 55977
rect 10385 55921 10441 55977
rect 10527 55921 10583 55977
rect 10669 55921 10725 55977
rect 10811 55921 10867 55977
rect 10953 55921 11009 55977
rect 11095 55921 11151 55977
rect 11237 55921 11293 55977
rect 11379 55921 11435 55977
rect 11521 55921 11577 55977
rect 11663 55921 11719 55977
rect 11805 55921 11861 55977
rect 11947 55921 12003 55977
rect 12089 55921 12145 55977
rect 12231 55921 12287 55977
rect 12373 55921 12429 55977
rect 12515 55921 12571 55977
rect 12657 55921 12713 55977
rect 12799 55921 12855 55977
rect 12941 55921 12997 55977
rect 13083 55921 13139 55977
rect 13225 55921 13281 55977
rect 13367 55921 13423 55977
rect 13509 55921 13565 55977
rect 13651 55921 13707 55977
rect 13793 55921 13849 55977
rect 13935 55921 13991 55977
rect 14077 55921 14133 55977
rect 14219 55921 14275 55977
rect 14361 55921 14417 55977
rect 14503 55921 14559 55977
rect 14645 55921 14701 55977
rect 14787 55921 14843 55977
rect 161 55779 217 55835
rect 303 55779 359 55835
rect 445 55779 501 55835
rect 587 55779 643 55835
rect 729 55779 785 55835
rect 871 55779 927 55835
rect 1013 55779 1069 55835
rect 1155 55779 1211 55835
rect 1297 55779 1353 55835
rect 1439 55779 1495 55835
rect 1581 55779 1637 55835
rect 1723 55779 1779 55835
rect 1865 55779 1921 55835
rect 2007 55779 2063 55835
rect 2149 55779 2205 55835
rect 2291 55779 2347 55835
rect 2433 55779 2489 55835
rect 2575 55779 2631 55835
rect 2717 55779 2773 55835
rect 2859 55779 2915 55835
rect 3001 55779 3057 55835
rect 3143 55779 3199 55835
rect 3285 55779 3341 55835
rect 3427 55779 3483 55835
rect 3569 55779 3625 55835
rect 3711 55779 3767 55835
rect 3853 55779 3909 55835
rect 3995 55779 4051 55835
rect 4137 55779 4193 55835
rect 4279 55779 4335 55835
rect 4421 55779 4477 55835
rect 4563 55779 4619 55835
rect 4705 55779 4761 55835
rect 4847 55779 4903 55835
rect 4989 55779 5045 55835
rect 5131 55779 5187 55835
rect 5273 55779 5329 55835
rect 5415 55779 5471 55835
rect 5557 55779 5613 55835
rect 5699 55779 5755 55835
rect 5841 55779 5897 55835
rect 5983 55779 6039 55835
rect 6125 55779 6181 55835
rect 6267 55779 6323 55835
rect 6409 55779 6465 55835
rect 6551 55779 6607 55835
rect 6693 55779 6749 55835
rect 6835 55779 6891 55835
rect 6977 55779 7033 55835
rect 7119 55779 7175 55835
rect 7261 55779 7317 55835
rect 7403 55779 7459 55835
rect 7545 55779 7601 55835
rect 7687 55779 7743 55835
rect 7829 55779 7885 55835
rect 7971 55779 8027 55835
rect 8113 55779 8169 55835
rect 8255 55779 8311 55835
rect 8397 55779 8453 55835
rect 8539 55779 8595 55835
rect 8681 55779 8737 55835
rect 8823 55779 8879 55835
rect 8965 55779 9021 55835
rect 9107 55779 9163 55835
rect 9249 55779 9305 55835
rect 9391 55779 9447 55835
rect 9533 55779 9589 55835
rect 9675 55779 9731 55835
rect 9817 55779 9873 55835
rect 9959 55779 10015 55835
rect 10101 55779 10157 55835
rect 10243 55779 10299 55835
rect 10385 55779 10441 55835
rect 10527 55779 10583 55835
rect 10669 55779 10725 55835
rect 10811 55779 10867 55835
rect 10953 55779 11009 55835
rect 11095 55779 11151 55835
rect 11237 55779 11293 55835
rect 11379 55779 11435 55835
rect 11521 55779 11577 55835
rect 11663 55779 11719 55835
rect 11805 55779 11861 55835
rect 11947 55779 12003 55835
rect 12089 55779 12145 55835
rect 12231 55779 12287 55835
rect 12373 55779 12429 55835
rect 12515 55779 12571 55835
rect 12657 55779 12713 55835
rect 12799 55779 12855 55835
rect 12941 55779 12997 55835
rect 13083 55779 13139 55835
rect 13225 55779 13281 55835
rect 13367 55779 13423 55835
rect 13509 55779 13565 55835
rect 13651 55779 13707 55835
rect 13793 55779 13849 55835
rect 13935 55779 13991 55835
rect 14077 55779 14133 55835
rect 14219 55779 14275 55835
rect 14361 55779 14417 55835
rect 14503 55779 14559 55835
rect 14645 55779 14701 55835
rect 14787 55779 14843 55835
rect 161 55637 217 55693
rect 303 55637 359 55693
rect 445 55637 501 55693
rect 587 55637 643 55693
rect 729 55637 785 55693
rect 871 55637 927 55693
rect 1013 55637 1069 55693
rect 1155 55637 1211 55693
rect 1297 55637 1353 55693
rect 1439 55637 1495 55693
rect 1581 55637 1637 55693
rect 1723 55637 1779 55693
rect 1865 55637 1921 55693
rect 2007 55637 2063 55693
rect 2149 55637 2205 55693
rect 2291 55637 2347 55693
rect 2433 55637 2489 55693
rect 2575 55637 2631 55693
rect 2717 55637 2773 55693
rect 2859 55637 2915 55693
rect 3001 55637 3057 55693
rect 3143 55637 3199 55693
rect 3285 55637 3341 55693
rect 3427 55637 3483 55693
rect 3569 55637 3625 55693
rect 3711 55637 3767 55693
rect 3853 55637 3909 55693
rect 3995 55637 4051 55693
rect 4137 55637 4193 55693
rect 4279 55637 4335 55693
rect 4421 55637 4477 55693
rect 4563 55637 4619 55693
rect 4705 55637 4761 55693
rect 4847 55637 4903 55693
rect 4989 55637 5045 55693
rect 5131 55637 5187 55693
rect 5273 55637 5329 55693
rect 5415 55637 5471 55693
rect 5557 55637 5613 55693
rect 5699 55637 5755 55693
rect 5841 55637 5897 55693
rect 5983 55637 6039 55693
rect 6125 55637 6181 55693
rect 6267 55637 6323 55693
rect 6409 55637 6465 55693
rect 6551 55637 6607 55693
rect 6693 55637 6749 55693
rect 6835 55637 6891 55693
rect 6977 55637 7033 55693
rect 7119 55637 7175 55693
rect 7261 55637 7317 55693
rect 7403 55637 7459 55693
rect 7545 55637 7601 55693
rect 7687 55637 7743 55693
rect 7829 55637 7885 55693
rect 7971 55637 8027 55693
rect 8113 55637 8169 55693
rect 8255 55637 8311 55693
rect 8397 55637 8453 55693
rect 8539 55637 8595 55693
rect 8681 55637 8737 55693
rect 8823 55637 8879 55693
rect 8965 55637 9021 55693
rect 9107 55637 9163 55693
rect 9249 55637 9305 55693
rect 9391 55637 9447 55693
rect 9533 55637 9589 55693
rect 9675 55637 9731 55693
rect 9817 55637 9873 55693
rect 9959 55637 10015 55693
rect 10101 55637 10157 55693
rect 10243 55637 10299 55693
rect 10385 55637 10441 55693
rect 10527 55637 10583 55693
rect 10669 55637 10725 55693
rect 10811 55637 10867 55693
rect 10953 55637 11009 55693
rect 11095 55637 11151 55693
rect 11237 55637 11293 55693
rect 11379 55637 11435 55693
rect 11521 55637 11577 55693
rect 11663 55637 11719 55693
rect 11805 55637 11861 55693
rect 11947 55637 12003 55693
rect 12089 55637 12145 55693
rect 12231 55637 12287 55693
rect 12373 55637 12429 55693
rect 12515 55637 12571 55693
rect 12657 55637 12713 55693
rect 12799 55637 12855 55693
rect 12941 55637 12997 55693
rect 13083 55637 13139 55693
rect 13225 55637 13281 55693
rect 13367 55637 13423 55693
rect 13509 55637 13565 55693
rect 13651 55637 13707 55693
rect 13793 55637 13849 55693
rect 13935 55637 13991 55693
rect 14077 55637 14133 55693
rect 14219 55637 14275 55693
rect 14361 55637 14417 55693
rect 14503 55637 14559 55693
rect 14645 55637 14701 55693
rect 14787 55637 14843 55693
rect 161 55307 217 55363
rect 303 55307 359 55363
rect 445 55307 501 55363
rect 587 55307 643 55363
rect 729 55307 785 55363
rect 871 55307 927 55363
rect 1013 55307 1069 55363
rect 1155 55307 1211 55363
rect 1297 55307 1353 55363
rect 1439 55307 1495 55363
rect 1581 55307 1637 55363
rect 1723 55307 1779 55363
rect 1865 55307 1921 55363
rect 2007 55307 2063 55363
rect 2149 55307 2205 55363
rect 2291 55307 2347 55363
rect 2433 55307 2489 55363
rect 2575 55307 2631 55363
rect 2717 55307 2773 55363
rect 2859 55307 2915 55363
rect 3001 55307 3057 55363
rect 3143 55307 3199 55363
rect 3285 55307 3341 55363
rect 3427 55307 3483 55363
rect 3569 55307 3625 55363
rect 3711 55307 3767 55363
rect 3853 55307 3909 55363
rect 3995 55307 4051 55363
rect 4137 55307 4193 55363
rect 4279 55307 4335 55363
rect 4421 55307 4477 55363
rect 4563 55307 4619 55363
rect 4705 55307 4761 55363
rect 4847 55307 4903 55363
rect 4989 55307 5045 55363
rect 5131 55307 5187 55363
rect 5273 55307 5329 55363
rect 5415 55307 5471 55363
rect 5557 55307 5613 55363
rect 5699 55307 5755 55363
rect 5841 55307 5897 55363
rect 5983 55307 6039 55363
rect 6125 55307 6181 55363
rect 6267 55307 6323 55363
rect 6409 55307 6465 55363
rect 6551 55307 6607 55363
rect 6693 55307 6749 55363
rect 6835 55307 6891 55363
rect 6977 55307 7033 55363
rect 7119 55307 7175 55363
rect 7261 55307 7317 55363
rect 7403 55307 7459 55363
rect 7545 55307 7601 55363
rect 7687 55307 7743 55363
rect 7829 55307 7885 55363
rect 7971 55307 8027 55363
rect 8113 55307 8169 55363
rect 8255 55307 8311 55363
rect 8397 55307 8453 55363
rect 8539 55307 8595 55363
rect 8681 55307 8737 55363
rect 8823 55307 8879 55363
rect 8965 55307 9021 55363
rect 9107 55307 9163 55363
rect 9249 55307 9305 55363
rect 9391 55307 9447 55363
rect 9533 55307 9589 55363
rect 9675 55307 9731 55363
rect 9817 55307 9873 55363
rect 9959 55307 10015 55363
rect 10101 55307 10157 55363
rect 10243 55307 10299 55363
rect 10385 55307 10441 55363
rect 10527 55307 10583 55363
rect 10669 55307 10725 55363
rect 10811 55307 10867 55363
rect 10953 55307 11009 55363
rect 11095 55307 11151 55363
rect 11237 55307 11293 55363
rect 11379 55307 11435 55363
rect 11521 55307 11577 55363
rect 11663 55307 11719 55363
rect 11805 55307 11861 55363
rect 11947 55307 12003 55363
rect 12089 55307 12145 55363
rect 12231 55307 12287 55363
rect 12373 55307 12429 55363
rect 12515 55307 12571 55363
rect 12657 55307 12713 55363
rect 12799 55307 12855 55363
rect 12941 55307 12997 55363
rect 13083 55307 13139 55363
rect 13225 55307 13281 55363
rect 13367 55307 13423 55363
rect 13509 55307 13565 55363
rect 13651 55307 13707 55363
rect 13793 55307 13849 55363
rect 13935 55307 13991 55363
rect 14077 55307 14133 55363
rect 14219 55307 14275 55363
rect 14361 55307 14417 55363
rect 14503 55307 14559 55363
rect 14645 55307 14701 55363
rect 14787 55307 14843 55363
rect 161 55165 217 55221
rect 303 55165 359 55221
rect 445 55165 501 55221
rect 587 55165 643 55221
rect 729 55165 785 55221
rect 871 55165 927 55221
rect 1013 55165 1069 55221
rect 1155 55165 1211 55221
rect 1297 55165 1353 55221
rect 1439 55165 1495 55221
rect 1581 55165 1637 55221
rect 1723 55165 1779 55221
rect 1865 55165 1921 55221
rect 2007 55165 2063 55221
rect 2149 55165 2205 55221
rect 2291 55165 2347 55221
rect 2433 55165 2489 55221
rect 2575 55165 2631 55221
rect 2717 55165 2773 55221
rect 2859 55165 2915 55221
rect 3001 55165 3057 55221
rect 3143 55165 3199 55221
rect 3285 55165 3341 55221
rect 3427 55165 3483 55221
rect 3569 55165 3625 55221
rect 3711 55165 3767 55221
rect 3853 55165 3909 55221
rect 3995 55165 4051 55221
rect 4137 55165 4193 55221
rect 4279 55165 4335 55221
rect 4421 55165 4477 55221
rect 4563 55165 4619 55221
rect 4705 55165 4761 55221
rect 4847 55165 4903 55221
rect 4989 55165 5045 55221
rect 5131 55165 5187 55221
rect 5273 55165 5329 55221
rect 5415 55165 5471 55221
rect 5557 55165 5613 55221
rect 5699 55165 5755 55221
rect 5841 55165 5897 55221
rect 5983 55165 6039 55221
rect 6125 55165 6181 55221
rect 6267 55165 6323 55221
rect 6409 55165 6465 55221
rect 6551 55165 6607 55221
rect 6693 55165 6749 55221
rect 6835 55165 6891 55221
rect 6977 55165 7033 55221
rect 7119 55165 7175 55221
rect 7261 55165 7317 55221
rect 7403 55165 7459 55221
rect 7545 55165 7601 55221
rect 7687 55165 7743 55221
rect 7829 55165 7885 55221
rect 7971 55165 8027 55221
rect 8113 55165 8169 55221
rect 8255 55165 8311 55221
rect 8397 55165 8453 55221
rect 8539 55165 8595 55221
rect 8681 55165 8737 55221
rect 8823 55165 8879 55221
rect 8965 55165 9021 55221
rect 9107 55165 9163 55221
rect 9249 55165 9305 55221
rect 9391 55165 9447 55221
rect 9533 55165 9589 55221
rect 9675 55165 9731 55221
rect 9817 55165 9873 55221
rect 9959 55165 10015 55221
rect 10101 55165 10157 55221
rect 10243 55165 10299 55221
rect 10385 55165 10441 55221
rect 10527 55165 10583 55221
rect 10669 55165 10725 55221
rect 10811 55165 10867 55221
rect 10953 55165 11009 55221
rect 11095 55165 11151 55221
rect 11237 55165 11293 55221
rect 11379 55165 11435 55221
rect 11521 55165 11577 55221
rect 11663 55165 11719 55221
rect 11805 55165 11861 55221
rect 11947 55165 12003 55221
rect 12089 55165 12145 55221
rect 12231 55165 12287 55221
rect 12373 55165 12429 55221
rect 12515 55165 12571 55221
rect 12657 55165 12713 55221
rect 12799 55165 12855 55221
rect 12941 55165 12997 55221
rect 13083 55165 13139 55221
rect 13225 55165 13281 55221
rect 13367 55165 13423 55221
rect 13509 55165 13565 55221
rect 13651 55165 13707 55221
rect 13793 55165 13849 55221
rect 13935 55165 13991 55221
rect 14077 55165 14133 55221
rect 14219 55165 14275 55221
rect 14361 55165 14417 55221
rect 14503 55165 14559 55221
rect 14645 55165 14701 55221
rect 14787 55165 14843 55221
rect 161 55023 217 55079
rect 303 55023 359 55079
rect 445 55023 501 55079
rect 587 55023 643 55079
rect 729 55023 785 55079
rect 871 55023 927 55079
rect 1013 55023 1069 55079
rect 1155 55023 1211 55079
rect 1297 55023 1353 55079
rect 1439 55023 1495 55079
rect 1581 55023 1637 55079
rect 1723 55023 1779 55079
rect 1865 55023 1921 55079
rect 2007 55023 2063 55079
rect 2149 55023 2205 55079
rect 2291 55023 2347 55079
rect 2433 55023 2489 55079
rect 2575 55023 2631 55079
rect 2717 55023 2773 55079
rect 2859 55023 2915 55079
rect 3001 55023 3057 55079
rect 3143 55023 3199 55079
rect 3285 55023 3341 55079
rect 3427 55023 3483 55079
rect 3569 55023 3625 55079
rect 3711 55023 3767 55079
rect 3853 55023 3909 55079
rect 3995 55023 4051 55079
rect 4137 55023 4193 55079
rect 4279 55023 4335 55079
rect 4421 55023 4477 55079
rect 4563 55023 4619 55079
rect 4705 55023 4761 55079
rect 4847 55023 4903 55079
rect 4989 55023 5045 55079
rect 5131 55023 5187 55079
rect 5273 55023 5329 55079
rect 5415 55023 5471 55079
rect 5557 55023 5613 55079
rect 5699 55023 5755 55079
rect 5841 55023 5897 55079
rect 5983 55023 6039 55079
rect 6125 55023 6181 55079
rect 6267 55023 6323 55079
rect 6409 55023 6465 55079
rect 6551 55023 6607 55079
rect 6693 55023 6749 55079
rect 6835 55023 6891 55079
rect 6977 55023 7033 55079
rect 7119 55023 7175 55079
rect 7261 55023 7317 55079
rect 7403 55023 7459 55079
rect 7545 55023 7601 55079
rect 7687 55023 7743 55079
rect 7829 55023 7885 55079
rect 7971 55023 8027 55079
rect 8113 55023 8169 55079
rect 8255 55023 8311 55079
rect 8397 55023 8453 55079
rect 8539 55023 8595 55079
rect 8681 55023 8737 55079
rect 8823 55023 8879 55079
rect 8965 55023 9021 55079
rect 9107 55023 9163 55079
rect 9249 55023 9305 55079
rect 9391 55023 9447 55079
rect 9533 55023 9589 55079
rect 9675 55023 9731 55079
rect 9817 55023 9873 55079
rect 9959 55023 10015 55079
rect 10101 55023 10157 55079
rect 10243 55023 10299 55079
rect 10385 55023 10441 55079
rect 10527 55023 10583 55079
rect 10669 55023 10725 55079
rect 10811 55023 10867 55079
rect 10953 55023 11009 55079
rect 11095 55023 11151 55079
rect 11237 55023 11293 55079
rect 11379 55023 11435 55079
rect 11521 55023 11577 55079
rect 11663 55023 11719 55079
rect 11805 55023 11861 55079
rect 11947 55023 12003 55079
rect 12089 55023 12145 55079
rect 12231 55023 12287 55079
rect 12373 55023 12429 55079
rect 12515 55023 12571 55079
rect 12657 55023 12713 55079
rect 12799 55023 12855 55079
rect 12941 55023 12997 55079
rect 13083 55023 13139 55079
rect 13225 55023 13281 55079
rect 13367 55023 13423 55079
rect 13509 55023 13565 55079
rect 13651 55023 13707 55079
rect 13793 55023 13849 55079
rect 13935 55023 13991 55079
rect 14077 55023 14133 55079
rect 14219 55023 14275 55079
rect 14361 55023 14417 55079
rect 14503 55023 14559 55079
rect 14645 55023 14701 55079
rect 14787 55023 14843 55079
rect 161 54881 217 54937
rect 303 54881 359 54937
rect 445 54881 501 54937
rect 587 54881 643 54937
rect 729 54881 785 54937
rect 871 54881 927 54937
rect 1013 54881 1069 54937
rect 1155 54881 1211 54937
rect 1297 54881 1353 54937
rect 1439 54881 1495 54937
rect 1581 54881 1637 54937
rect 1723 54881 1779 54937
rect 1865 54881 1921 54937
rect 2007 54881 2063 54937
rect 2149 54881 2205 54937
rect 2291 54881 2347 54937
rect 2433 54881 2489 54937
rect 2575 54881 2631 54937
rect 2717 54881 2773 54937
rect 2859 54881 2915 54937
rect 3001 54881 3057 54937
rect 3143 54881 3199 54937
rect 3285 54881 3341 54937
rect 3427 54881 3483 54937
rect 3569 54881 3625 54937
rect 3711 54881 3767 54937
rect 3853 54881 3909 54937
rect 3995 54881 4051 54937
rect 4137 54881 4193 54937
rect 4279 54881 4335 54937
rect 4421 54881 4477 54937
rect 4563 54881 4619 54937
rect 4705 54881 4761 54937
rect 4847 54881 4903 54937
rect 4989 54881 5045 54937
rect 5131 54881 5187 54937
rect 5273 54881 5329 54937
rect 5415 54881 5471 54937
rect 5557 54881 5613 54937
rect 5699 54881 5755 54937
rect 5841 54881 5897 54937
rect 5983 54881 6039 54937
rect 6125 54881 6181 54937
rect 6267 54881 6323 54937
rect 6409 54881 6465 54937
rect 6551 54881 6607 54937
rect 6693 54881 6749 54937
rect 6835 54881 6891 54937
rect 6977 54881 7033 54937
rect 7119 54881 7175 54937
rect 7261 54881 7317 54937
rect 7403 54881 7459 54937
rect 7545 54881 7601 54937
rect 7687 54881 7743 54937
rect 7829 54881 7885 54937
rect 7971 54881 8027 54937
rect 8113 54881 8169 54937
rect 8255 54881 8311 54937
rect 8397 54881 8453 54937
rect 8539 54881 8595 54937
rect 8681 54881 8737 54937
rect 8823 54881 8879 54937
rect 8965 54881 9021 54937
rect 9107 54881 9163 54937
rect 9249 54881 9305 54937
rect 9391 54881 9447 54937
rect 9533 54881 9589 54937
rect 9675 54881 9731 54937
rect 9817 54881 9873 54937
rect 9959 54881 10015 54937
rect 10101 54881 10157 54937
rect 10243 54881 10299 54937
rect 10385 54881 10441 54937
rect 10527 54881 10583 54937
rect 10669 54881 10725 54937
rect 10811 54881 10867 54937
rect 10953 54881 11009 54937
rect 11095 54881 11151 54937
rect 11237 54881 11293 54937
rect 11379 54881 11435 54937
rect 11521 54881 11577 54937
rect 11663 54881 11719 54937
rect 11805 54881 11861 54937
rect 11947 54881 12003 54937
rect 12089 54881 12145 54937
rect 12231 54881 12287 54937
rect 12373 54881 12429 54937
rect 12515 54881 12571 54937
rect 12657 54881 12713 54937
rect 12799 54881 12855 54937
rect 12941 54881 12997 54937
rect 13083 54881 13139 54937
rect 13225 54881 13281 54937
rect 13367 54881 13423 54937
rect 13509 54881 13565 54937
rect 13651 54881 13707 54937
rect 13793 54881 13849 54937
rect 13935 54881 13991 54937
rect 14077 54881 14133 54937
rect 14219 54881 14275 54937
rect 14361 54881 14417 54937
rect 14503 54881 14559 54937
rect 14645 54881 14701 54937
rect 14787 54881 14843 54937
rect 161 54739 217 54795
rect 303 54739 359 54795
rect 445 54739 501 54795
rect 587 54739 643 54795
rect 729 54739 785 54795
rect 871 54739 927 54795
rect 1013 54739 1069 54795
rect 1155 54739 1211 54795
rect 1297 54739 1353 54795
rect 1439 54739 1495 54795
rect 1581 54739 1637 54795
rect 1723 54739 1779 54795
rect 1865 54739 1921 54795
rect 2007 54739 2063 54795
rect 2149 54739 2205 54795
rect 2291 54739 2347 54795
rect 2433 54739 2489 54795
rect 2575 54739 2631 54795
rect 2717 54739 2773 54795
rect 2859 54739 2915 54795
rect 3001 54739 3057 54795
rect 3143 54739 3199 54795
rect 3285 54739 3341 54795
rect 3427 54739 3483 54795
rect 3569 54739 3625 54795
rect 3711 54739 3767 54795
rect 3853 54739 3909 54795
rect 3995 54739 4051 54795
rect 4137 54739 4193 54795
rect 4279 54739 4335 54795
rect 4421 54739 4477 54795
rect 4563 54739 4619 54795
rect 4705 54739 4761 54795
rect 4847 54739 4903 54795
rect 4989 54739 5045 54795
rect 5131 54739 5187 54795
rect 5273 54739 5329 54795
rect 5415 54739 5471 54795
rect 5557 54739 5613 54795
rect 5699 54739 5755 54795
rect 5841 54739 5897 54795
rect 5983 54739 6039 54795
rect 6125 54739 6181 54795
rect 6267 54739 6323 54795
rect 6409 54739 6465 54795
rect 6551 54739 6607 54795
rect 6693 54739 6749 54795
rect 6835 54739 6891 54795
rect 6977 54739 7033 54795
rect 7119 54739 7175 54795
rect 7261 54739 7317 54795
rect 7403 54739 7459 54795
rect 7545 54739 7601 54795
rect 7687 54739 7743 54795
rect 7829 54739 7885 54795
rect 7971 54739 8027 54795
rect 8113 54739 8169 54795
rect 8255 54739 8311 54795
rect 8397 54739 8453 54795
rect 8539 54739 8595 54795
rect 8681 54739 8737 54795
rect 8823 54739 8879 54795
rect 8965 54739 9021 54795
rect 9107 54739 9163 54795
rect 9249 54739 9305 54795
rect 9391 54739 9447 54795
rect 9533 54739 9589 54795
rect 9675 54739 9731 54795
rect 9817 54739 9873 54795
rect 9959 54739 10015 54795
rect 10101 54739 10157 54795
rect 10243 54739 10299 54795
rect 10385 54739 10441 54795
rect 10527 54739 10583 54795
rect 10669 54739 10725 54795
rect 10811 54739 10867 54795
rect 10953 54739 11009 54795
rect 11095 54739 11151 54795
rect 11237 54739 11293 54795
rect 11379 54739 11435 54795
rect 11521 54739 11577 54795
rect 11663 54739 11719 54795
rect 11805 54739 11861 54795
rect 11947 54739 12003 54795
rect 12089 54739 12145 54795
rect 12231 54739 12287 54795
rect 12373 54739 12429 54795
rect 12515 54739 12571 54795
rect 12657 54739 12713 54795
rect 12799 54739 12855 54795
rect 12941 54739 12997 54795
rect 13083 54739 13139 54795
rect 13225 54739 13281 54795
rect 13367 54739 13423 54795
rect 13509 54739 13565 54795
rect 13651 54739 13707 54795
rect 13793 54739 13849 54795
rect 13935 54739 13991 54795
rect 14077 54739 14133 54795
rect 14219 54739 14275 54795
rect 14361 54739 14417 54795
rect 14503 54739 14559 54795
rect 14645 54739 14701 54795
rect 14787 54739 14843 54795
rect 161 54597 217 54653
rect 303 54597 359 54653
rect 445 54597 501 54653
rect 587 54597 643 54653
rect 729 54597 785 54653
rect 871 54597 927 54653
rect 1013 54597 1069 54653
rect 1155 54597 1211 54653
rect 1297 54597 1353 54653
rect 1439 54597 1495 54653
rect 1581 54597 1637 54653
rect 1723 54597 1779 54653
rect 1865 54597 1921 54653
rect 2007 54597 2063 54653
rect 2149 54597 2205 54653
rect 2291 54597 2347 54653
rect 2433 54597 2489 54653
rect 2575 54597 2631 54653
rect 2717 54597 2773 54653
rect 2859 54597 2915 54653
rect 3001 54597 3057 54653
rect 3143 54597 3199 54653
rect 3285 54597 3341 54653
rect 3427 54597 3483 54653
rect 3569 54597 3625 54653
rect 3711 54597 3767 54653
rect 3853 54597 3909 54653
rect 3995 54597 4051 54653
rect 4137 54597 4193 54653
rect 4279 54597 4335 54653
rect 4421 54597 4477 54653
rect 4563 54597 4619 54653
rect 4705 54597 4761 54653
rect 4847 54597 4903 54653
rect 4989 54597 5045 54653
rect 5131 54597 5187 54653
rect 5273 54597 5329 54653
rect 5415 54597 5471 54653
rect 5557 54597 5613 54653
rect 5699 54597 5755 54653
rect 5841 54597 5897 54653
rect 5983 54597 6039 54653
rect 6125 54597 6181 54653
rect 6267 54597 6323 54653
rect 6409 54597 6465 54653
rect 6551 54597 6607 54653
rect 6693 54597 6749 54653
rect 6835 54597 6891 54653
rect 6977 54597 7033 54653
rect 7119 54597 7175 54653
rect 7261 54597 7317 54653
rect 7403 54597 7459 54653
rect 7545 54597 7601 54653
rect 7687 54597 7743 54653
rect 7829 54597 7885 54653
rect 7971 54597 8027 54653
rect 8113 54597 8169 54653
rect 8255 54597 8311 54653
rect 8397 54597 8453 54653
rect 8539 54597 8595 54653
rect 8681 54597 8737 54653
rect 8823 54597 8879 54653
rect 8965 54597 9021 54653
rect 9107 54597 9163 54653
rect 9249 54597 9305 54653
rect 9391 54597 9447 54653
rect 9533 54597 9589 54653
rect 9675 54597 9731 54653
rect 9817 54597 9873 54653
rect 9959 54597 10015 54653
rect 10101 54597 10157 54653
rect 10243 54597 10299 54653
rect 10385 54597 10441 54653
rect 10527 54597 10583 54653
rect 10669 54597 10725 54653
rect 10811 54597 10867 54653
rect 10953 54597 11009 54653
rect 11095 54597 11151 54653
rect 11237 54597 11293 54653
rect 11379 54597 11435 54653
rect 11521 54597 11577 54653
rect 11663 54597 11719 54653
rect 11805 54597 11861 54653
rect 11947 54597 12003 54653
rect 12089 54597 12145 54653
rect 12231 54597 12287 54653
rect 12373 54597 12429 54653
rect 12515 54597 12571 54653
rect 12657 54597 12713 54653
rect 12799 54597 12855 54653
rect 12941 54597 12997 54653
rect 13083 54597 13139 54653
rect 13225 54597 13281 54653
rect 13367 54597 13423 54653
rect 13509 54597 13565 54653
rect 13651 54597 13707 54653
rect 13793 54597 13849 54653
rect 13935 54597 13991 54653
rect 14077 54597 14133 54653
rect 14219 54597 14275 54653
rect 14361 54597 14417 54653
rect 14503 54597 14559 54653
rect 14645 54597 14701 54653
rect 14787 54597 14843 54653
rect 161 54455 217 54511
rect 303 54455 359 54511
rect 445 54455 501 54511
rect 587 54455 643 54511
rect 729 54455 785 54511
rect 871 54455 927 54511
rect 1013 54455 1069 54511
rect 1155 54455 1211 54511
rect 1297 54455 1353 54511
rect 1439 54455 1495 54511
rect 1581 54455 1637 54511
rect 1723 54455 1779 54511
rect 1865 54455 1921 54511
rect 2007 54455 2063 54511
rect 2149 54455 2205 54511
rect 2291 54455 2347 54511
rect 2433 54455 2489 54511
rect 2575 54455 2631 54511
rect 2717 54455 2773 54511
rect 2859 54455 2915 54511
rect 3001 54455 3057 54511
rect 3143 54455 3199 54511
rect 3285 54455 3341 54511
rect 3427 54455 3483 54511
rect 3569 54455 3625 54511
rect 3711 54455 3767 54511
rect 3853 54455 3909 54511
rect 3995 54455 4051 54511
rect 4137 54455 4193 54511
rect 4279 54455 4335 54511
rect 4421 54455 4477 54511
rect 4563 54455 4619 54511
rect 4705 54455 4761 54511
rect 4847 54455 4903 54511
rect 4989 54455 5045 54511
rect 5131 54455 5187 54511
rect 5273 54455 5329 54511
rect 5415 54455 5471 54511
rect 5557 54455 5613 54511
rect 5699 54455 5755 54511
rect 5841 54455 5897 54511
rect 5983 54455 6039 54511
rect 6125 54455 6181 54511
rect 6267 54455 6323 54511
rect 6409 54455 6465 54511
rect 6551 54455 6607 54511
rect 6693 54455 6749 54511
rect 6835 54455 6891 54511
rect 6977 54455 7033 54511
rect 7119 54455 7175 54511
rect 7261 54455 7317 54511
rect 7403 54455 7459 54511
rect 7545 54455 7601 54511
rect 7687 54455 7743 54511
rect 7829 54455 7885 54511
rect 7971 54455 8027 54511
rect 8113 54455 8169 54511
rect 8255 54455 8311 54511
rect 8397 54455 8453 54511
rect 8539 54455 8595 54511
rect 8681 54455 8737 54511
rect 8823 54455 8879 54511
rect 8965 54455 9021 54511
rect 9107 54455 9163 54511
rect 9249 54455 9305 54511
rect 9391 54455 9447 54511
rect 9533 54455 9589 54511
rect 9675 54455 9731 54511
rect 9817 54455 9873 54511
rect 9959 54455 10015 54511
rect 10101 54455 10157 54511
rect 10243 54455 10299 54511
rect 10385 54455 10441 54511
rect 10527 54455 10583 54511
rect 10669 54455 10725 54511
rect 10811 54455 10867 54511
rect 10953 54455 11009 54511
rect 11095 54455 11151 54511
rect 11237 54455 11293 54511
rect 11379 54455 11435 54511
rect 11521 54455 11577 54511
rect 11663 54455 11719 54511
rect 11805 54455 11861 54511
rect 11947 54455 12003 54511
rect 12089 54455 12145 54511
rect 12231 54455 12287 54511
rect 12373 54455 12429 54511
rect 12515 54455 12571 54511
rect 12657 54455 12713 54511
rect 12799 54455 12855 54511
rect 12941 54455 12997 54511
rect 13083 54455 13139 54511
rect 13225 54455 13281 54511
rect 13367 54455 13423 54511
rect 13509 54455 13565 54511
rect 13651 54455 13707 54511
rect 13793 54455 13849 54511
rect 13935 54455 13991 54511
rect 14077 54455 14133 54511
rect 14219 54455 14275 54511
rect 14361 54455 14417 54511
rect 14503 54455 14559 54511
rect 14645 54455 14701 54511
rect 14787 54455 14843 54511
rect 161 54313 217 54369
rect 303 54313 359 54369
rect 445 54313 501 54369
rect 587 54313 643 54369
rect 729 54313 785 54369
rect 871 54313 927 54369
rect 1013 54313 1069 54369
rect 1155 54313 1211 54369
rect 1297 54313 1353 54369
rect 1439 54313 1495 54369
rect 1581 54313 1637 54369
rect 1723 54313 1779 54369
rect 1865 54313 1921 54369
rect 2007 54313 2063 54369
rect 2149 54313 2205 54369
rect 2291 54313 2347 54369
rect 2433 54313 2489 54369
rect 2575 54313 2631 54369
rect 2717 54313 2773 54369
rect 2859 54313 2915 54369
rect 3001 54313 3057 54369
rect 3143 54313 3199 54369
rect 3285 54313 3341 54369
rect 3427 54313 3483 54369
rect 3569 54313 3625 54369
rect 3711 54313 3767 54369
rect 3853 54313 3909 54369
rect 3995 54313 4051 54369
rect 4137 54313 4193 54369
rect 4279 54313 4335 54369
rect 4421 54313 4477 54369
rect 4563 54313 4619 54369
rect 4705 54313 4761 54369
rect 4847 54313 4903 54369
rect 4989 54313 5045 54369
rect 5131 54313 5187 54369
rect 5273 54313 5329 54369
rect 5415 54313 5471 54369
rect 5557 54313 5613 54369
rect 5699 54313 5755 54369
rect 5841 54313 5897 54369
rect 5983 54313 6039 54369
rect 6125 54313 6181 54369
rect 6267 54313 6323 54369
rect 6409 54313 6465 54369
rect 6551 54313 6607 54369
rect 6693 54313 6749 54369
rect 6835 54313 6891 54369
rect 6977 54313 7033 54369
rect 7119 54313 7175 54369
rect 7261 54313 7317 54369
rect 7403 54313 7459 54369
rect 7545 54313 7601 54369
rect 7687 54313 7743 54369
rect 7829 54313 7885 54369
rect 7971 54313 8027 54369
rect 8113 54313 8169 54369
rect 8255 54313 8311 54369
rect 8397 54313 8453 54369
rect 8539 54313 8595 54369
rect 8681 54313 8737 54369
rect 8823 54313 8879 54369
rect 8965 54313 9021 54369
rect 9107 54313 9163 54369
rect 9249 54313 9305 54369
rect 9391 54313 9447 54369
rect 9533 54313 9589 54369
rect 9675 54313 9731 54369
rect 9817 54313 9873 54369
rect 9959 54313 10015 54369
rect 10101 54313 10157 54369
rect 10243 54313 10299 54369
rect 10385 54313 10441 54369
rect 10527 54313 10583 54369
rect 10669 54313 10725 54369
rect 10811 54313 10867 54369
rect 10953 54313 11009 54369
rect 11095 54313 11151 54369
rect 11237 54313 11293 54369
rect 11379 54313 11435 54369
rect 11521 54313 11577 54369
rect 11663 54313 11719 54369
rect 11805 54313 11861 54369
rect 11947 54313 12003 54369
rect 12089 54313 12145 54369
rect 12231 54313 12287 54369
rect 12373 54313 12429 54369
rect 12515 54313 12571 54369
rect 12657 54313 12713 54369
rect 12799 54313 12855 54369
rect 12941 54313 12997 54369
rect 13083 54313 13139 54369
rect 13225 54313 13281 54369
rect 13367 54313 13423 54369
rect 13509 54313 13565 54369
rect 13651 54313 13707 54369
rect 13793 54313 13849 54369
rect 13935 54313 13991 54369
rect 14077 54313 14133 54369
rect 14219 54313 14275 54369
rect 14361 54313 14417 54369
rect 14503 54313 14559 54369
rect 14645 54313 14701 54369
rect 14787 54313 14843 54369
rect 161 54171 217 54227
rect 303 54171 359 54227
rect 445 54171 501 54227
rect 587 54171 643 54227
rect 729 54171 785 54227
rect 871 54171 927 54227
rect 1013 54171 1069 54227
rect 1155 54171 1211 54227
rect 1297 54171 1353 54227
rect 1439 54171 1495 54227
rect 1581 54171 1637 54227
rect 1723 54171 1779 54227
rect 1865 54171 1921 54227
rect 2007 54171 2063 54227
rect 2149 54171 2205 54227
rect 2291 54171 2347 54227
rect 2433 54171 2489 54227
rect 2575 54171 2631 54227
rect 2717 54171 2773 54227
rect 2859 54171 2915 54227
rect 3001 54171 3057 54227
rect 3143 54171 3199 54227
rect 3285 54171 3341 54227
rect 3427 54171 3483 54227
rect 3569 54171 3625 54227
rect 3711 54171 3767 54227
rect 3853 54171 3909 54227
rect 3995 54171 4051 54227
rect 4137 54171 4193 54227
rect 4279 54171 4335 54227
rect 4421 54171 4477 54227
rect 4563 54171 4619 54227
rect 4705 54171 4761 54227
rect 4847 54171 4903 54227
rect 4989 54171 5045 54227
rect 5131 54171 5187 54227
rect 5273 54171 5329 54227
rect 5415 54171 5471 54227
rect 5557 54171 5613 54227
rect 5699 54171 5755 54227
rect 5841 54171 5897 54227
rect 5983 54171 6039 54227
rect 6125 54171 6181 54227
rect 6267 54171 6323 54227
rect 6409 54171 6465 54227
rect 6551 54171 6607 54227
rect 6693 54171 6749 54227
rect 6835 54171 6891 54227
rect 6977 54171 7033 54227
rect 7119 54171 7175 54227
rect 7261 54171 7317 54227
rect 7403 54171 7459 54227
rect 7545 54171 7601 54227
rect 7687 54171 7743 54227
rect 7829 54171 7885 54227
rect 7971 54171 8027 54227
rect 8113 54171 8169 54227
rect 8255 54171 8311 54227
rect 8397 54171 8453 54227
rect 8539 54171 8595 54227
rect 8681 54171 8737 54227
rect 8823 54171 8879 54227
rect 8965 54171 9021 54227
rect 9107 54171 9163 54227
rect 9249 54171 9305 54227
rect 9391 54171 9447 54227
rect 9533 54171 9589 54227
rect 9675 54171 9731 54227
rect 9817 54171 9873 54227
rect 9959 54171 10015 54227
rect 10101 54171 10157 54227
rect 10243 54171 10299 54227
rect 10385 54171 10441 54227
rect 10527 54171 10583 54227
rect 10669 54171 10725 54227
rect 10811 54171 10867 54227
rect 10953 54171 11009 54227
rect 11095 54171 11151 54227
rect 11237 54171 11293 54227
rect 11379 54171 11435 54227
rect 11521 54171 11577 54227
rect 11663 54171 11719 54227
rect 11805 54171 11861 54227
rect 11947 54171 12003 54227
rect 12089 54171 12145 54227
rect 12231 54171 12287 54227
rect 12373 54171 12429 54227
rect 12515 54171 12571 54227
rect 12657 54171 12713 54227
rect 12799 54171 12855 54227
rect 12941 54171 12997 54227
rect 13083 54171 13139 54227
rect 13225 54171 13281 54227
rect 13367 54171 13423 54227
rect 13509 54171 13565 54227
rect 13651 54171 13707 54227
rect 13793 54171 13849 54227
rect 13935 54171 13991 54227
rect 14077 54171 14133 54227
rect 14219 54171 14275 54227
rect 14361 54171 14417 54227
rect 14503 54171 14559 54227
rect 14645 54171 14701 54227
rect 14787 54171 14843 54227
rect 161 54029 217 54085
rect 303 54029 359 54085
rect 445 54029 501 54085
rect 587 54029 643 54085
rect 729 54029 785 54085
rect 871 54029 927 54085
rect 1013 54029 1069 54085
rect 1155 54029 1211 54085
rect 1297 54029 1353 54085
rect 1439 54029 1495 54085
rect 1581 54029 1637 54085
rect 1723 54029 1779 54085
rect 1865 54029 1921 54085
rect 2007 54029 2063 54085
rect 2149 54029 2205 54085
rect 2291 54029 2347 54085
rect 2433 54029 2489 54085
rect 2575 54029 2631 54085
rect 2717 54029 2773 54085
rect 2859 54029 2915 54085
rect 3001 54029 3057 54085
rect 3143 54029 3199 54085
rect 3285 54029 3341 54085
rect 3427 54029 3483 54085
rect 3569 54029 3625 54085
rect 3711 54029 3767 54085
rect 3853 54029 3909 54085
rect 3995 54029 4051 54085
rect 4137 54029 4193 54085
rect 4279 54029 4335 54085
rect 4421 54029 4477 54085
rect 4563 54029 4619 54085
rect 4705 54029 4761 54085
rect 4847 54029 4903 54085
rect 4989 54029 5045 54085
rect 5131 54029 5187 54085
rect 5273 54029 5329 54085
rect 5415 54029 5471 54085
rect 5557 54029 5613 54085
rect 5699 54029 5755 54085
rect 5841 54029 5897 54085
rect 5983 54029 6039 54085
rect 6125 54029 6181 54085
rect 6267 54029 6323 54085
rect 6409 54029 6465 54085
rect 6551 54029 6607 54085
rect 6693 54029 6749 54085
rect 6835 54029 6891 54085
rect 6977 54029 7033 54085
rect 7119 54029 7175 54085
rect 7261 54029 7317 54085
rect 7403 54029 7459 54085
rect 7545 54029 7601 54085
rect 7687 54029 7743 54085
rect 7829 54029 7885 54085
rect 7971 54029 8027 54085
rect 8113 54029 8169 54085
rect 8255 54029 8311 54085
rect 8397 54029 8453 54085
rect 8539 54029 8595 54085
rect 8681 54029 8737 54085
rect 8823 54029 8879 54085
rect 8965 54029 9021 54085
rect 9107 54029 9163 54085
rect 9249 54029 9305 54085
rect 9391 54029 9447 54085
rect 9533 54029 9589 54085
rect 9675 54029 9731 54085
rect 9817 54029 9873 54085
rect 9959 54029 10015 54085
rect 10101 54029 10157 54085
rect 10243 54029 10299 54085
rect 10385 54029 10441 54085
rect 10527 54029 10583 54085
rect 10669 54029 10725 54085
rect 10811 54029 10867 54085
rect 10953 54029 11009 54085
rect 11095 54029 11151 54085
rect 11237 54029 11293 54085
rect 11379 54029 11435 54085
rect 11521 54029 11577 54085
rect 11663 54029 11719 54085
rect 11805 54029 11861 54085
rect 11947 54029 12003 54085
rect 12089 54029 12145 54085
rect 12231 54029 12287 54085
rect 12373 54029 12429 54085
rect 12515 54029 12571 54085
rect 12657 54029 12713 54085
rect 12799 54029 12855 54085
rect 12941 54029 12997 54085
rect 13083 54029 13139 54085
rect 13225 54029 13281 54085
rect 13367 54029 13423 54085
rect 13509 54029 13565 54085
rect 13651 54029 13707 54085
rect 13793 54029 13849 54085
rect 13935 54029 13991 54085
rect 14077 54029 14133 54085
rect 14219 54029 14275 54085
rect 14361 54029 14417 54085
rect 14503 54029 14559 54085
rect 14645 54029 14701 54085
rect 14787 54029 14843 54085
rect 161 53715 217 53771
rect 303 53715 359 53771
rect 445 53715 501 53771
rect 587 53715 643 53771
rect 729 53715 785 53771
rect 871 53715 927 53771
rect 1013 53715 1069 53771
rect 1155 53715 1211 53771
rect 1297 53715 1353 53771
rect 1439 53715 1495 53771
rect 1581 53715 1637 53771
rect 1723 53715 1779 53771
rect 1865 53715 1921 53771
rect 2007 53715 2063 53771
rect 2149 53715 2205 53771
rect 2291 53715 2347 53771
rect 2433 53715 2489 53771
rect 2575 53715 2631 53771
rect 2717 53715 2773 53771
rect 2859 53715 2915 53771
rect 3001 53715 3057 53771
rect 3143 53715 3199 53771
rect 3285 53715 3341 53771
rect 3427 53715 3483 53771
rect 3569 53715 3625 53771
rect 3711 53715 3767 53771
rect 3853 53715 3909 53771
rect 3995 53715 4051 53771
rect 4137 53715 4193 53771
rect 4279 53715 4335 53771
rect 4421 53715 4477 53771
rect 4563 53715 4619 53771
rect 4705 53715 4761 53771
rect 4847 53715 4903 53771
rect 4989 53715 5045 53771
rect 5131 53715 5187 53771
rect 5273 53715 5329 53771
rect 5415 53715 5471 53771
rect 5557 53715 5613 53771
rect 5699 53715 5755 53771
rect 5841 53715 5897 53771
rect 5983 53715 6039 53771
rect 6125 53715 6181 53771
rect 6267 53715 6323 53771
rect 6409 53715 6465 53771
rect 6551 53715 6607 53771
rect 6693 53715 6749 53771
rect 6835 53715 6891 53771
rect 6977 53715 7033 53771
rect 7119 53715 7175 53771
rect 7261 53715 7317 53771
rect 7403 53715 7459 53771
rect 7545 53715 7601 53771
rect 7687 53715 7743 53771
rect 7829 53715 7885 53771
rect 7971 53715 8027 53771
rect 8113 53715 8169 53771
rect 8255 53715 8311 53771
rect 8397 53715 8453 53771
rect 8539 53715 8595 53771
rect 8681 53715 8737 53771
rect 8823 53715 8879 53771
rect 8965 53715 9021 53771
rect 9107 53715 9163 53771
rect 9249 53715 9305 53771
rect 9391 53715 9447 53771
rect 9533 53715 9589 53771
rect 9675 53715 9731 53771
rect 9817 53715 9873 53771
rect 9959 53715 10015 53771
rect 10101 53715 10157 53771
rect 10243 53715 10299 53771
rect 10385 53715 10441 53771
rect 10527 53715 10583 53771
rect 10669 53715 10725 53771
rect 10811 53715 10867 53771
rect 10953 53715 11009 53771
rect 11095 53715 11151 53771
rect 11237 53715 11293 53771
rect 11379 53715 11435 53771
rect 11521 53715 11577 53771
rect 11663 53715 11719 53771
rect 11805 53715 11861 53771
rect 11947 53715 12003 53771
rect 12089 53715 12145 53771
rect 12231 53715 12287 53771
rect 12373 53715 12429 53771
rect 12515 53715 12571 53771
rect 12657 53715 12713 53771
rect 12799 53715 12855 53771
rect 12941 53715 12997 53771
rect 13083 53715 13139 53771
rect 13225 53715 13281 53771
rect 13367 53715 13423 53771
rect 13509 53715 13565 53771
rect 13651 53715 13707 53771
rect 13793 53715 13849 53771
rect 13935 53715 13991 53771
rect 14077 53715 14133 53771
rect 14219 53715 14275 53771
rect 14361 53715 14417 53771
rect 14503 53715 14559 53771
rect 14645 53715 14701 53771
rect 14787 53715 14843 53771
rect 161 53573 217 53629
rect 303 53573 359 53629
rect 445 53573 501 53629
rect 587 53573 643 53629
rect 729 53573 785 53629
rect 871 53573 927 53629
rect 1013 53573 1069 53629
rect 1155 53573 1211 53629
rect 1297 53573 1353 53629
rect 1439 53573 1495 53629
rect 1581 53573 1637 53629
rect 1723 53573 1779 53629
rect 1865 53573 1921 53629
rect 2007 53573 2063 53629
rect 2149 53573 2205 53629
rect 2291 53573 2347 53629
rect 2433 53573 2489 53629
rect 2575 53573 2631 53629
rect 2717 53573 2773 53629
rect 2859 53573 2915 53629
rect 3001 53573 3057 53629
rect 3143 53573 3199 53629
rect 3285 53573 3341 53629
rect 3427 53573 3483 53629
rect 3569 53573 3625 53629
rect 3711 53573 3767 53629
rect 3853 53573 3909 53629
rect 3995 53573 4051 53629
rect 4137 53573 4193 53629
rect 4279 53573 4335 53629
rect 4421 53573 4477 53629
rect 4563 53573 4619 53629
rect 4705 53573 4761 53629
rect 4847 53573 4903 53629
rect 4989 53573 5045 53629
rect 5131 53573 5187 53629
rect 5273 53573 5329 53629
rect 5415 53573 5471 53629
rect 5557 53573 5613 53629
rect 5699 53573 5755 53629
rect 5841 53573 5897 53629
rect 5983 53573 6039 53629
rect 6125 53573 6181 53629
rect 6267 53573 6323 53629
rect 6409 53573 6465 53629
rect 6551 53573 6607 53629
rect 6693 53573 6749 53629
rect 6835 53573 6891 53629
rect 6977 53573 7033 53629
rect 7119 53573 7175 53629
rect 7261 53573 7317 53629
rect 7403 53573 7459 53629
rect 7545 53573 7601 53629
rect 7687 53573 7743 53629
rect 7829 53573 7885 53629
rect 7971 53573 8027 53629
rect 8113 53573 8169 53629
rect 8255 53573 8311 53629
rect 8397 53573 8453 53629
rect 8539 53573 8595 53629
rect 8681 53573 8737 53629
rect 8823 53573 8879 53629
rect 8965 53573 9021 53629
rect 9107 53573 9163 53629
rect 9249 53573 9305 53629
rect 9391 53573 9447 53629
rect 9533 53573 9589 53629
rect 9675 53573 9731 53629
rect 9817 53573 9873 53629
rect 9959 53573 10015 53629
rect 10101 53573 10157 53629
rect 10243 53573 10299 53629
rect 10385 53573 10441 53629
rect 10527 53573 10583 53629
rect 10669 53573 10725 53629
rect 10811 53573 10867 53629
rect 10953 53573 11009 53629
rect 11095 53573 11151 53629
rect 11237 53573 11293 53629
rect 11379 53573 11435 53629
rect 11521 53573 11577 53629
rect 11663 53573 11719 53629
rect 11805 53573 11861 53629
rect 11947 53573 12003 53629
rect 12089 53573 12145 53629
rect 12231 53573 12287 53629
rect 12373 53573 12429 53629
rect 12515 53573 12571 53629
rect 12657 53573 12713 53629
rect 12799 53573 12855 53629
rect 12941 53573 12997 53629
rect 13083 53573 13139 53629
rect 13225 53573 13281 53629
rect 13367 53573 13423 53629
rect 13509 53573 13565 53629
rect 13651 53573 13707 53629
rect 13793 53573 13849 53629
rect 13935 53573 13991 53629
rect 14077 53573 14133 53629
rect 14219 53573 14275 53629
rect 14361 53573 14417 53629
rect 14503 53573 14559 53629
rect 14645 53573 14701 53629
rect 14787 53573 14843 53629
rect 161 53431 217 53487
rect 303 53431 359 53487
rect 445 53431 501 53487
rect 587 53431 643 53487
rect 729 53431 785 53487
rect 871 53431 927 53487
rect 1013 53431 1069 53487
rect 1155 53431 1211 53487
rect 1297 53431 1353 53487
rect 1439 53431 1495 53487
rect 1581 53431 1637 53487
rect 1723 53431 1779 53487
rect 1865 53431 1921 53487
rect 2007 53431 2063 53487
rect 2149 53431 2205 53487
rect 2291 53431 2347 53487
rect 2433 53431 2489 53487
rect 2575 53431 2631 53487
rect 2717 53431 2773 53487
rect 2859 53431 2915 53487
rect 3001 53431 3057 53487
rect 3143 53431 3199 53487
rect 3285 53431 3341 53487
rect 3427 53431 3483 53487
rect 3569 53431 3625 53487
rect 3711 53431 3767 53487
rect 3853 53431 3909 53487
rect 3995 53431 4051 53487
rect 4137 53431 4193 53487
rect 4279 53431 4335 53487
rect 4421 53431 4477 53487
rect 4563 53431 4619 53487
rect 4705 53431 4761 53487
rect 4847 53431 4903 53487
rect 4989 53431 5045 53487
rect 5131 53431 5187 53487
rect 5273 53431 5329 53487
rect 5415 53431 5471 53487
rect 5557 53431 5613 53487
rect 5699 53431 5755 53487
rect 5841 53431 5897 53487
rect 5983 53431 6039 53487
rect 6125 53431 6181 53487
rect 6267 53431 6323 53487
rect 6409 53431 6465 53487
rect 6551 53431 6607 53487
rect 6693 53431 6749 53487
rect 6835 53431 6891 53487
rect 6977 53431 7033 53487
rect 7119 53431 7175 53487
rect 7261 53431 7317 53487
rect 7403 53431 7459 53487
rect 7545 53431 7601 53487
rect 7687 53431 7743 53487
rect 7829 53431 7885 53487
rect 7971 53431 8027 53487
rect 8113 53431 8169 53487
rect 8255 53431 8311 53487
rect 8397 53431 8453 53487
rect 8539 53431 8595 53487
rect 8681 53431 8737 53487
rect 8823 53431 8879 53487
rect 8965 53431 9021 53487
rect 9107 53431 9163 53487
rect 9249 53431 9305 53487
rect 9391 53431 9447 53487
rect 9533 53431 9589 53487
rect 9675 53431 9731 53487
rect 9817 53431 9873 53487
rect 9959 53431 10015 53487
rect 10101 53431 10157 53487
rect 10243 53431 10299 53487
rect 10385 53431 10441 53487
rect 10527 53431 10583 53487
rect 10669 53431 10725 53487
rect 10811 53431 10867 53487
rect 10953 53431 11009 53487
rect 11095 53431 11151 53487
rect 11237 53431 11293 53487
rect 11379 53431 11435 53487
rect 11521 53431 11577 53487
rect 11663 53431 11719 53487
rect 11805 53431 11861 53487
rect 11947 53431 12003 53487
rect 12089 53431 12145 53487
rect 12231 53431 12287 53487
rect 12373 53431 12429 53487
rect 12515 53431 12571 53487
rect 12657 53431 12713 53487
rect 12799 53431 12855 53487
rect 12941 53431 12997 53487
rect 13083 53431 13139 53487
rect 13225 53431 13281 53487
rect 13367 53431 13423 53487
rect 13509 53431 13565 53487
rect 13651 53431 13707 53487
rect 13793 53431 13849 53487
rect 13935 53431 13991 53487
rect 14077 53431 14133 53487
rect 14219 53431 14275 53487
rect 14361 53431 14417 53487
rect 14503 53431 14559 53487
rect 14645 53431 14701 53487
rect 14787 53431 14843 53487
rect 161 53289 217 53345
rect 303 53289 359 53345
rect 445 53289 501 53345
rect 587 53289 643 53345
rect 729 53289 785 53345
rect 871 53289 927 53345
rect 1013 53289 1069 53345
rect 1155 53289 1211 53345
rect 1297 53289 1353 53345
rect 1439 53289 1495 53345
rect 1581 53289 1637 53345
rect 1723 53289 1779 53345
rect 1865 53289 1921 53345
rect 2007 53289 2063 53345
rect 2149 53289 2205 53345
rect 2291 53289 2347 53345
rect 2433 53289 2489 53345
rect 2575 53289 2631 53345
rect 2717 53289 2773 53345
rect 2859 53289 2915 53345
rect 3001 53289 3057 53345
rect 3143 53289 3199 53345
rect 3285 53289 3341 53345
rect 3427 53289 3483 53345
rect 3569 53289 3625 53345
rect 3711 53289 3767 53345
rect 3853 53289 3909 53345
rect 3995 53289 4051 53345
rect 4137 53289 4193 53345
rect 4279 53289 4335 53345
rect 4421 53289 4477 53345
rect 4563 53289 4619 53345
rect 4705 53289 4761 53345
rect 4847 53289 4903 53345
rect 4989 53289 5045 53345
rect 5131 53289 5187 53345
rect 5273 53289 5329 53345
rect 5415 53289 5471 53345
rect 5557 53289 5613 53345
rect 5699 53289 5755 53345
rect 5841 53289 5897 53345
rect 5983 53289 6039 53345
rect 6125 53289 6181 53345
rect 6267 53289 6323 53345
rect 6409 53289 6465 53345
rect 6551 53289 6607 53345
rect 6693 53289 6749 53345
rect 6835 53289 6891 53345
rect 6977 53289 7033 53345
rect 7119 53289 7175 53345
rect 7261 53289 7317 53345
rect 7403 53289 7459 53345
rect 7545 53289 7601 53345
rect 7687 53289 7743 53345
rect 7829 53289 7885 53345
rect 7971 53289 8027 53345
rect 8113 53289 8169 53345
rect 8255 53289 8311 53345
rect 8397 53289 8453 53345
rect 8539 53289 8595 53345
rect 8681 53289 8737 53345
rect 8823 53289 8879 53345
rect 8965 53289 9021 53345
rect 9107 53289 9163 53345
rect 9249 53289 9305 53345
rect 9391 53289 9447 53345
rect 9533 53289 9589 53345
rect 9675 53289 9731 53345
rect 9817 53289 9873 53345
rect 9959 53289 10015 53345
rect 10101 53289 10157 53345
rect 10243 53289 10299 53345
rect 10385 53289 10441 53345
rect 10527 53289 10583 53345
rect 10669 53289 10725 53345
rect 10811 53289 10867 53345
rect 10953 53289 11009 53345
rect 11095 53289 11151 53345
rect 11237 53289 11293 53345
rect 11379 53289 11435 53345
rect 11521 53289 11577 53345
rect 11663 53289 11719 53345
rect 11805 53289 11861 53345
rect 11947 53289 12003 53345
rect 12089 53289 12145 53345
rect 12231 53289 12287 53345
rect 12373 53289 12429 53345
rect 12515 53289 12571 53345
rect 12657 53289 12713 53345
rect 12799 53289 12855 53345
rect 12941 53289 12997 53345
rect 13083 53289 13139 53345
rect 13225 53289 13281 53345
rect 13367 53289 13423 53345
rect 13509 53289 13565 53345
rect 13651 53289 13707 53345
rect 13793 53289 13849 53345
rect 13935 53289 13991 53345
rect 14077 53289 14133 53345
rect 14219 53289 14275 53345
rect 14361 53289 14417 53345
rect 14503 53289 14559 53345
rect 14645 53289 14701 53345
rect 14787 53289 14843 53345
rect 161 53147 217 53203
rect 303 53147 359 53203
rect 445 53147 501 53203
rect 587 53147 643 53203
rect 729 53147 785 53203
rect 871 53147 927 53203
rect 1013 53147 1069 53203
rect 1155 53147 1211 53203
rect 1297 53147 1353 53203
rect 1439 53147 1495 53203
rect 1581 53147 1637 53203
rect 1723 53147 1779 53203
rect 1865 53147 1921 53203
rect 2007 53147 2063 53203
rect 2149 53147 2205 53203
rect 2291 53147 2347 53203
rect 2433 53147 2489 53203
rect 2575 53147 2631 53203
rect 2717 53147 2773 53203
rect 2859 53147 2915 53203
rect 3001 53147 3057 53203
rect 3143 53147 3199 53203
rect 3285 53147 3341 53203
rect 3427 53147 3483 53203
rect 3569 53147 3625 53203
rect 3711 53147 3767 53203
rect 3853 53147 3909 53203
rect 3995 53147 4051 53203
rect 4137 53147 4193 53203
rect 4279 53147 4335 53203
rect 4421 53147 4477 53203
rect 4563 53147 4619 53203
rect 4705 53147 4761 53203
rect 4847 53147 4903 53203
rect 4989 53147 5045 53203
rect 5131 53147 5187 53203
rect 5273 53147 5329 53203
rect 5415 53147 5471 53203
rect 5557 53147 5613 53203
rect 5699 53147 5755 53203
rect 5841 53147 5897 53203
rect 5983 53147 6039 53203
rect 6125 53147 6181 53203
rect 6267 53147 6323 53203
rect 6409 53147 6465 53203
rect 6551 53147 6607 53203
rect 6693 53147 6749 53203
rect 6835 53147 6891 53203
rect 6977 53147 7033 53203
rect 7119 53147 7175 53203
rect 7261 53147 7317 53203
rect 7403 53147 7459 53203
rect 7545 53147 7601 53203
rect 7687 53147 7743 53203
rect 7829 53147 7885 53203
rect 7971 53147 8027 53203
rect 8113 53147 8169 53203
rect 8255 53147 8311 53203
rect 8397 53147 8453 53203
rect 8539 53147 8595 53203
rect 8681 53147 8737 53203
rect 8823 53147 8879 53203
rect 8965 53147 9021 53203
rect 9107 53147 9163 53203
rect 9249 53147 9305 53203
rect 9391 53147 9447 53203
rect 9533 53147 9589 53203
rect 9675 53147 9731 53203
rect 9817 53147 9873 53203
rect 9959 53147 10015 53203
rect 10101 53147 10157 53203
rect 10243 53147 10299 53203
rect 10385 53147 10441 53203
rect 10527 53147 10583 53203
rect 10669 53147 10725 53203
rect 10811 53147 10867 53203
rect 10953 53147 11009 53203
rect 11095 53147 11151 53203
rect 11237 53147 11293 53203
rect 11379 53147 11435 53203
rect 11521 53147 11577 53203
rect 11663 53147 11719 53203
rect 11805 53147 11861 53203
rect 11947 53147 12003 53203
rect 12089 53147 12145 53203
rect 12231 53147 12287 53203
rect 12373 53147 12429 53203
rect 12515 53147 12571 53203
rect 12657 53147 12713 53203
rect 12799 53147 12855 53203
rect 12941 53147 12997 53203
rect 13083 53147 13139 53203
rect 13225 53147 13281 53203
rect 13367 53147 13423 53203
rect 13509 53147 13565 53203
rect 13651 53147 13707 53203
rect 13793 53147 13849 53203
rect 13935 53147 13991 53203
rect 14077 53147 14133 53203
rect 14219 53147 14275 53203
rect 14361 53147 14417 53203
rect 14503 53147 14559 53203
rect 14645 53147 14701 53203
rect 14787 53147 14843 53203
rect 161 53005 217 53061
rect 303 53005 359 53061
rect 445 53005 501 53061
rect 587 53005 643 53061
rect 729 53005 785 53061
rect 871 53005 927 53061
rect 1013 53005 1069 53061
rect 1155 53005 1211 53061
rect 1297 53005 1353 53061
rect 1439 53005 1495 53061
rect 1581 53005 1637 53061
rect 1723 53005 1779 53061
rect 1865 53005 1921 53061
rect 2007 53005 2063 53061
rect 2149 53005 2205 53061
rect 2291 53005 2347 53061
rect 2433 53005 2489 53061
rect 2575 53005 2631 53061
rect 2717 53005 2773 53061
rect 2859 53005 2915 53061
rect 3001 53005 3057 53061
rect 3143 53005 3199 53061
rect 3285 53005 3341 53061
rect 3427 53005 3483 53061
rect 3569 53005 3625 53061
rect 3711 53005 3767 53061
rect 3853 53005 3909 53061
rect 3995 53005 4051 53061
rect 4137 53005 4193 53061
rect 4279 53005 4335 53061
rect 4421 53005 4477 53061
rect 4563 53005 4619 53061
rect 4705 53005 4761 53061
rect 4847 53005 4903 53061
rect 4989 53005 5045 53061
rect 5131 53005 5187 53061
rect 5273 53005 5329 53061
rect 5415 53005 5471 53061
rect 5557 53005 5613 53061
rect 5699 53005 5755 53061
rect 5841 53005 5897 53061
rect 5983 53005 6039 53061
rect 6125 53005 6181 53061
rect 6267 53005 6323 53061
rect 6409 53005 6465 53061
rect 6551 53005 6607 53061
rect 6693 53005 6749 53061
rect 6835 53005 6891 53061
rect 6977 53005 7033 53061
rect 7119 53005 7175 53061
rect 7261 53005 7317 53061
rect 7403 53005 7459 53061
rect 7545 53005 7601 53061
rect 7687 53005 7743 53061
rect 7829 53005 7885 53061
rect 7971 53005 8027 53061
rect 8113 53005 8169 53061
rect 8255 53005 8311 53061
rect 8397 53005 8453 53061
rect 8539 53005 8595 53061
rect 8681 53005 8737 53061
rect 8823 53005 8879 53061
rect 8965 53005 9021 53061
rect 9107 53005 9163 53061
rect 9249 53005 9305 53061
rect 9391 53005 9447 53061
rect 9533 53005 9589 53061
rect 9675 53005 9731 53061
rect 9817 53005 9873 53061
rect 9959 53005 10015 53061
rect 10101 53005 10157 53061
rect 10243 53005 10299 53061
rect 10385 53005 10441 53061
rect 10527 53005 10583 53061
rect 10669 53005 10725 53061
rect 10811 53005 10867 53061
rect 10953 53005 11009 53061
rect 11095 53005 11151 53061
rect 11237 53005 11293 53061
rect 11379 53005 11435 53061
rect 11521 53005 11577 53061
rect 11663 53005 11719 53061
rect 11805 53005 11861 53061
rect 11947 53005 12003 53061
rect 12089 53005 12145 53061
rect 12231 53005 12287 53061
rect 12373 53005 12429 53061
rect 12515 53005 12571 53061
rect 12657 53005 12713 53061
rect 12799 53005 12855 53061
rect 12941 53005 12997 53061
rect 13083 53005 13139 53061
rect 13225 53005 13281 53061
rect 13367 53005 13423 53061
rect 13509 53005 13565 53061
rect 13651 53005 13707 53061
rect 13793 53005 13849 53061
rect 13935 53005 13991 53061
rect 14077 53005 14133 53061
rect 14219 53005 14275 53061
rect 14361 53005 14417 53061
rect 14503 53005 14559 53061
rect 14645 53005 14701 53061
rect 14787 53005 14843 53061
rect 161 52863 217 52919
rect 303 52863 359 52919
rect 445 52863 501 52919
rect 587 52863 643 52919
rect 729 52863 785 52919
rect 871 52863 927 52919
rect 1013 52863 1069 52919
rect 1155 52863 1211 52919
rect 1297 52863 1353 52919
rect 1439 52863 1495 52919
rect 1581 52863 1637 52919
rect 1723 52863 1779 52919
rect 1865 52863 1921 52919
rect 2007 52863 2063 52919
rect 2149 52863 2205 52919
rect 2291 52863 2347 52919
rect 2433 52863 2489 52919
rect 2575 52863 2631 52919
rect 2717 52863 2773 52919
rect 2859 52863 2915 52919
rect 3001 52863 3057 52919
rect 3143 52863 3199 52919
rect 3285 52863 3341 52919
rect 3427 52863 3483 52919
rect 3569 52863 3625 52919
rect 3711 52863 3767 52919
rect 3853 52863 3909 52919
rect 3995 52863 4051 52919
rect 4137 52863 4193 52919
rect 4279 52863 4335 52919
rect 4421 52863 4477 52919
rect 4563 52863 4619 52919
rect 4705 52863 4761 52919
rect 4847 52863 4903 52919
rect 4989 52863 5045 52919
rect 5131 52863 5187 52919
rect 5273 52863 5329 52919
rect 5415 52863 5471 52919
rect 5557 52863 5613 52919
rect 5699 52863 5755 52919
rect 5841 52863 5897 52919
rect 5983 52863 6039 52919
rect 6125 52863 6181 52919
rect 6267 52863 6323 52919
rect 6409 52863 6465 52919
rect 6551 52863 6607 52919
rect 6693 52863 6749 52919
rect 6835 52863 6891 52919
rect 6977 52863 7033 52919
rect 7119 52863 7175 52919
rect 7261 52863 7317 52919
rect 7403 52863 7459 52919
rect 7545 52863 7601 52919
rect 7687 52863 7743 52919
rect 7829 52863 7885 52919
rect 7971 52863 8027 52919
rect 8113 52863 8169 52919
rect 8255 52863 8311 52919
rect 8397 52863 8453 52919
rect 8539 52863 8595 52919
rect 8681 52863 8737 52919
rect 8823 52863 8879 52919
rect 8965 52863 9021 52919
rect 9107 52863 9163 52919
rect 9249 52863 9305 52919
rect 9391 52863 9447 52919
rect 9533 52863 9589 52919
rect 9675 52863 9731 52919
rect 9817 52863 9873 52919
rect 9959 52863 10015 52919
rect 10101 52863 10157 52919
rect 10243 52863 10299 52919
rect 10385 52863 10441 52919
rect 10527 52863 10583 52919
rect 10669 52863 10725 52919
rect 10811 52863 10867 52919
rect 10953 52863 11009 52919
rect 11095 52863 11151 52919
rect 11237 52863 11293 52919
rect 11379 52863 11435 52919
rect 11521 52863 11577 52919
rect 11663 52863 11719 52919
rect 11805 52863 11861 52919
rect 11947 52863 12003 52919
rect 12089 52863 12145 52919
rect 12231 52863 12287 52919
rect 12373 52863 12429 52919
rect 12515 52863 12571 52919
rect 12657 52863 12713 52919
rect 12799 52863 12855 52919
rect 12941 52863 12997 52919
rect 13083 52863 13139 52919
rect 13225 52863 13281 52919
rect 13367 52863 13423 52919
rect 13509 52863 13565 52919
rect 13651 52863 13707 52919
rect 13793 52863 13849 52919
rect 13935 52863 13991 52919
rect 14077 52863 14133 52919
rect 14219 52863 14275 52919
rect 14361 52863 14417 52919
rect 14503 52863 14559 52919
rect 14645 52863 14701 52919
rect 14787 52863 14843 52919
rect 161 52721 217 52777
rect 303 52721 359 52777
rect 445 52721 501 52777
rect 587 52721 643 52777
rect 729 52721 785 52777
rect 871 52721 927 52777
rect 1013 52721 1069 52777
rect 1155 52721 1211 52777
rect 1297 52721 1353 52777
rect 1439 52721 1495 52777
rect 1581 52721 1637 52777
rect 1723 52721 1779 52777
rect 1865 52721 1921 52777
rect 2007 52721 2063 52777
rect 2149 52721 2205 52777
rect 2291 52721 2347 52777
rect 2433 52721 2489 52777
rect 2575 52721 2631 52777
rect 2717 52721 2773 52777
rect 2859 52721 2915 52777
rect 3001 52721 3057 52777
rect 3143 52721 3199 52777
rect 3285 52721 3341 52777
rect 3427 52721 3483 52777
rect 3569 52721 3625 52777
rect 3711 52721 3767 52777
rect 3853 52721 3909 52777
rect 3995 52721 4051 52777
rect 4137 52721 4193 52777
rect 4279 52721 4335 52777
rect 4421 52721 4477 52777
rect 4563 52721 4619 52777
rect 4705 52721 4761 52777
rect 4847 52721 4903 52777
rect 4989 52721 5045 52777
rect 5131 52721 5187 52777
rect 5273 52721 5329 52777
rect 5415 52721 5471 52777
rect 5557 52721 5613 52777
rect 5699 52721 5755 52777
rect 5841 52721 5897 52777
rect 5983 52721 6039 52777
rect 6125 52721 6181 52777
rect 6267 52721 6323 52777
rect 6409 52721 6465 52777
rect 6551 52721 6607 52777
rect 6693 52721 6749 52777
rect 6835 52721 6891 52777
rect 6977 52721 7033 52777
rect 7119 52721 7175 52777
rect 7261 52721 7317 52777
rect 7403 52721 7459 52777
rect 7545 52721 7601 52777
rect 7687 52721 7743 52777
rect 7829 52721 7885 52777
rect 7971 52721 8027 52777
rect 8113 52721 8169 52777
rect 8255 52721 8311 52777
rect 8397 52721 8453 52777
rect 8539 52721 8595 52777
rect 8681 52721 8737 52777
rect 8823 52721 8879 52777
rect 8965 52721 9021 52777
rect 9107 52721 9163 52777
rect 9249 52721 9305 52777
rect 9391 52721 9447 52777
rect 9533 52721 9589 52777
rect 9675 52721 9731 52777
rect 9817 52721 9873 52777
rect 9959 52721 10015 52777
rect 10101 52721 10157 52777
rect 10243 52721 10299 52777
rect 10385 52721 10441 52777
rect 10527 52721 10583 52777
rect 10669 52721 10725 52777
rect 10811 52721 10867 52777
rect 10953 52721 11009 52777
rect 11095 52721 11151 52777
rect 11237 52721 11293 52777
rect 11379 52721 11435 52777
rect 11521 52721 11577 52777
rect 11663 52721 11719 52777
rect 11805 52721 11861 52777
rect 11947 52721 12003 52777
rect 12089 52721 12145 52777
rect 12231 52721 12287 52777
rect 12373 52721 12429 52777
rect 12515 52721 12571 52777
rect 12657 52721 12713 52777
rect 12799 52721 12855 52777
rect 12941 52721 12997 52777
rect 13083 52721 13139 52777
rect 13225 52721 13281 52777
rect 13367 52721 13423 52777
rect 13509 52721 13565 52777
rect 13651 52721 13707 52777
rect 13793 52721 13849 52777
rect 13935 52721 13991 52777
rect 14077 52721 14133 52777
rect 14219 52721 14275 52777
rect 14361 52721 14417 52777
rect 14503 52721 14559 52777
rect 14645 52721 14701 52777
rect 14787 52721 14843 52777
rect 161 52579 217 52635
rect 303 52579 359 52635
rect 445 52579 501 52635
rect 587 52579 643 52635
rect 729 52579 785 52635
rect 871 52579 927 52635
rect 1013 52579 1069 52635
rect 1155 52579 1211 52635
rect 1297 52579 1353 52635
rect 1439 52579 1495 52635
rect 1581 52579 1637 52635
rect 1723 52579 1779 52635
rect 1865 52579 1921 52635
rect 2007 52579 2063 52635
rect 2149 52579 2205 52635
rect 2291 52579 2347 52635
rect 2433 52579 2489 52635
rect 2575 52579 2631 52635
rect 2717 52579 2773 52635
rect 2859 52579 2915 52635
rect 3001 52579 3057 52635
rect 3143 52579 3199 52635
rect 3285 52579 3341 52635
rect 3427 52579 3483 52635
rect 3569 52579 3625 52635
rect 3711 52579 3767 52635
rect 3853 52579 3909 52635
rect 3995 52579 4051 52635
rect 4137 52579 4193 52635
rect 4279 52579 4335 52635
rect 4421 52579 4477 52635
rect 4563 52579 4619 52635
rect 4705 52579 4761 52635
rect 4847 52579 4903 52635
rect 4989 52579 5045 52635
rect 5131 52579 5187 52635
rect 5273 52579 5329 52635
rect 5415 52579 5471 52635
rect 5557 52579 5613 52635
rect 5699 52579 5755 52635
rect 5841 52579 5897 52635
rect 5983 52579 6039 52635
rect 6125 52579 6181 52635
rect 6267 52579 6323 52635
rect 6409 52579 6465 52635
rect 6551 52579 6607 52635
rect 6693 52579 6749 52635
rect 6835 52579 6891 52635
rect 6977 52579 7033 52635
rect 7119 52579 7175 52635
rect 7261 52579 7317 52635
rect 7403 52579 7459 52635
rect 7545 52579 7601 52635
rect 7687 52579 7743 52635
rect 7829 52579 7885 52635
rect 7971 52579 8027 52635
rect 8113 52579 8169 52635
rect 8255 52579 8311 52635
rect 8397 52579 8453 52635
rect 8539 52579 8595 52635
rect 8681 52579 8737 52635
rect 8823 52579 8879 52635
rect 8965 52579 9021 52635
rect 9107 52579 9163 52635
rect 9249 52579 9305 52635
rect 9391 52579 9447 52635
rect 9533 52579 9589 52635
rect 9675 52579 9731 52635
rect 9817 52579 9873 52635
rect 9959 52579 10015 52635
rect 10101 52579 10157 52635
rect 10243 52579 10299 52635
rect 10385 52579 10441 52635
rect 10527 52579 10583 52635
rect 10669 52579 10725 52635
rect 10811 52579 10867 52635
rect 10953 52579 11009 52635
rect 11095 52579 11151 52635
rect 11237 52579 11293 52635
rect 11379 52579 11435 52635
rect 11521 52579 11577 52635
rect 11663 52579 11719 52635
rect 11805 52579 11861 52635
rect 11947 52579 12003 52635
rect 12089 52579 12145 52635
rect 12231 52579 12287 52635
rect 12373 52579 12429 52635
rect 12515 52579 12571 52635
rect 12657 52579 12713 52635
rect 12799 52579 12855 52635
rect 12941 52579 12997 52635
rect 13083 52579 13139 52635
rect 13225 52579 13281 52635
rect 13367 52579 13423 52635
rect 13509 52579 13565 52635
rect 13651 52579 13707 52635
rect 13793 52579 13849 52635
rect 13935 52579 13991 52635
rect 14077 52579 14133 52635
rect 14219 52579 14275 52635
rect 14361 52579 14417 52635
rect 14503 52579 14559 52635
rect 14645 52579 14701 52635
rect 14787 52579 14843 52635
rect 161 52437 217 52493
rect 303 52437 359 52493
rect 445 52437 501 52493
rect 587 52437 643 52493
rect 729 52437 785 52493
rect 871 52437 927 52493
rect 1013 52437 1069 52493
rect 1155 52437 1211 52493
rect 1297 52437 1353 52493
rect 1439 52437 1495 52493
rect 1581 52437 1637 52493
rect 1723 52437 1779 52493
rect 1865 52437 1921 52493
rect 2007 52437 2063 52493
rect 2149 52437 2205 52493
rect 2291 52437 2347 52493
rect 2433 52437 2489 52493
rect 2575 52437 2631 52493
rect 2717 52437 2773 52493
rect 2859 52437 2915 52493
rect 3001 52437 3057 52493
rect 3143 52437 3199 52493
rect 3285 52437 3341 52493
rect 3427 52437 3483 52493
rect 3569 52437 3625 52493
rect 3711 52437 3767 52493
rect 3853 52437 3909 52493
rect 3995 52437 4051 52493
rect 4137 52437 4193 52493
rect 4279 52437 4335 52493
rect 4421 52437 4477 52493
rect 4563 52437 4619 52493
rect 4705 52437 4761 52493
rect 4847 52437 4903 52493
rect 4989 52437 5045 52493
rect 5131 52437 5187 52493
rect 5273 52437 5329 52493
rect 5415 52437 5471 52493
rect 5557 52437 5613 52493
rect 5699 52437 5755 52493
rect 5841 52437 5897 52493
rect 5983 52437 6039 52493
rect 6125 52437 6181 52493
rect 6267 52437 6323 52493
rect 6409 52437 6465 52493
rect 6551 52437 6607 52493
rect 6693 52437 6749 52493
rect 6835 52437 6891 52493
rect 6977 52437 7033 52493
rect 7119 52437 7175 52493
rect 7261 52437 7317 52493
rect 7403 52437 7459 52493
rect 7545 52437 7601 52493
rect 7687 52437 7743 52493
rect 7829 52437 7885 52493
rect 7971 52437 8027 52493
rect 8113 52437 8169 52493
rect 8255 52437 8311 52493
rect 8397 52437 8453 52493
rect 8539 52437 8595 52493
rect 8681 52437 8737 52493
rect 8823 52437 8879 52493
rect 8965 52437 9021 52493
rect 9107 52437 9163 52493
rect 9249 52437 9305 52493
rect 9391 52437 9447 52493
rect 9533 52437 9589 52493
rect 9675 52437 9731 52493
rect 9817 52437 9873 52493
rect 9959 52437 10015 52493
rect 10101 52437 10157 52493
rect 10243 52437 10299 52493
rect 10385 52437 10441 52493
rect 10527 52437 10583 52493
rect 10669 52437 10725 52493
rect 10811 52437 10867 52493
rect 10953 52437 11009 52493
rect 11095 52437 11151 52493
rect 11237 52437 11293 52493
rect 11379 52437 11435 52493
rect 11521 52437 11577 52493
rect 11663 52437 11719 52493
rect 11805 52437 11861 52493
rect 11947 52437 12003 52493
rect 12089 52437 12145 52493
rect 12231 52437 12287 52493
rect 12373 52437 12429 52493
rect 12515 52437 12571 52493
rect 12657 52437 12713 52493
rect 12799 52437 12855 52493
rect 12941 52437 12997 52493
rect 13083 52437 13139 52493
rect 13225 52437 13281 52493
rect 13367 52437 13423 52493
rect 13509 52437 13565 52493
rect 13651 52437 13707 52493
rect 13793 52437 13849 52493
rect 13935 52437 13991 52493
rect 14077 52437 14133 52493
rect 14219 52437 14275 52493
rect 14361 52437 14417 52493
rect 14503 52437 14559 52493
rect 14645 52437 14701 52493
rect 14787 52437 14843 52493
rect 161 52107 217 52163
rect 303 52107 359 52163
rect 445 52107 501 52163
rect 587 52107 643 52163
rect 729 52107 785 52163
rect 871 52107 927 52163
rect 1013 52107 1069 52163
rect 1155 52107 1211 52163
rect 1297 52107 1353 52163
rect 1439 52107 1495 52163
rect 1581 52107 1637 52163
rect 1723 52107 1779 52163
rect 1865 52107 1921 52163
rect 2007 52107 2063 52163
rect 2149 52107 2205 52163
rect 2291 52107 2347 52163
rect 2433 52107 2489 52163
rect 2575 52107 2631 52163
rect 2717 52107 2773 52163
rect 2859 52107 2915 52163
rect 3001 52107 3057 52163
rect 3143 52107 3199 52163
rect 3285 52107 3341 52163
rect 3427 52107 3483 52163
rect 3569 52107 3625 52163
rect 3711 52107 3767 52163
rect 3853 52107 3909 52163
rect 3995 52107 4051 52163
rect 4137 52107 4193 52163
rect 4279 52107 4335 52163
rect 4421 52107 4477 52163
rect 4563 52107 4619 52163
rect 4705 52107 4761 52163
rect 4847 52107 4903 52163
rect 4989 52107 5045 52163
rect 5131 52107 5187 52163
rect 5273 52107 5329 52163
rect 5415 52107 5471 52163
rect 5557 52107 5613 52163
rect 5699 52107 5755 52163
rect 5841 52107 5897 52163
rect 5983 52107 6039 52163
rect 6125 52107 6181 52163
rect 6267 52107 6323 52163
rect 6409 52107 6465 52163
rect 6551 52107 6607 52163
rect 6693 52107 6749 52163
rect 6835 52107 6891 52163
rect 6977 52107 7033 52163
rect 7119 52107 7175 52163
rect 7261 52107 7317 52163
rect 7403 52107 7459 52163
rect 7545 52107 7601 52163
rect 7687 52107 7743 52163
rect 7829 52107 7885 52163
rect 7971 52107 8027 52163
rect 8113 52107 8169 52163
rect 8255 52107 8311 52163
rect 8397 52107 8453 52163
rect 8539 52107 8595 52163
rect 8681 52107 8737 52163
rect 8823 52107 8879 52163
rect 8965 52107 9021 52163
rect 9107 52107 9163 52163
rect 9249 52107 9305 52163
rect 9391 52107 9447 52163
rect 9533 52107 9589 52163
rect 9675 52107 9731 52163
rect 9817 52107 9873 52163
rect 9959 52107 10015 52163
rect 10101 52107 10157 52163
rect 10243 52107 10299 52163
rect 10385 52107 10441 52163
rect 10527 52107 10583 52163
rect 10669 52107 10725 52163
rect 10811 52107 10867 52163
rect 10953 52107 11009 52163
rect 11095 52107 11151 52163
rect 11237 52107 11293 52163
rect 11379 52107 11435 52163
rect 11521 52107 11577 52163
rect 11663 52107 11719 52163
rect 11805 52107 11861 52163
rect 11947 52107 12003 52163
rect 12089 52107 12145 52163
rect 12231 52107 12287 52163
rect 12373 52107 12429 52163
rect 12515 52107 12571 52163
rect 12657 52107 12713 52163
rect 12799 52107 12855 52163
rect 12941 52107 12997 52163
rect 13083 52107 13139 52163
rect 13225 52107 13281 52163
rect 13367 52107 13423 52163
rect 13509 52107 13565 52163
rect 13651 52107 13707 52163
rect 13793 52107 13849 52163
rect 13935 52107 13991 52163
rect 14077 52107 14133 52163
rect 14219 52107 14275 52163
rect 14361 52107 14417 52163
rect 14503 52107 14559 52163
rect 14645 52107 14701 52163
rect 14787 52107 14843 52163
rect 161 51965 217 52021
rect 303 51965 359 52021
rect 445 51965 501 52021
rect 587 51965 643 52021
rect 729 51965 785 52021
rect 871 51965 927 52021
rect 1013 51965 1069 52021
rect 1155 51965 1211 52021
rect 1297 51965 1353 52021
rect 1439 51965 1495 52021
rect 1581 51965 1637 52021
rect 1723 51965 1779 52021
rect 1865 51965 1921 52021
rect 2007 51965 2063 52021
rect 2149 51965 2205 52021
rect 2291 51965 2347 52021
rect 2433 51965 2489 52021
rect 2575 51965 2631 52021
rect 2717 51965 2773 52021
rect 2859 51965 2915 52021
rect 3001 51965 3057 52021
rect 3143 51965 3199 52021
rect 3285 51965 3341 52021
rect 3427 51965 3483 52021
rect 3569 51965 3625 52021
rect 3711 51965 3767 52021
rect 3853 51965 3909 52021
rect 3995 51965 4051 52021
rect 4137 51965 4193 52021
rect 4279 51965 4335 52021
rect 4421 51965 4477 52021
rect 4563 51965 4619 52021
rect 4705 51965 4761 52021
rect 4847 51965 4903 52021
rect 4989 51965 5045 52021
rect 5131 51965 5187 52021
rect 5273 51965 5329 52021
rect 5415 51965 5471 52021
rect 5557 51965 5613 52021
rect 5699 51965 5755 52021
rect 5841 51965 5897 52021
rect 5983 51965 6039 52021
rect 6125 51965 6181 52021
rect 6267 51965 6323 52021
rect 6409 51965 6465 52021
rect 6551 51965 6607 52021
rect 6693 51965 6749 52021
rect 6835 51965 6891 52021
rect 6977 51965 7033 52021
rect 7119 51965 7175 52021
rect 7261 51965 7317 52021
rect 7403 51965 7459 52021
rect 7545 51965 7601 52021
rect 7687 51965 7743 52021
rect 7829 51965 7885 52021
rect 7971 51965 8027 52021
rect 8113 51965 8169 52021
rect 8255 51965 8311 52021
rect 8397 51965 8453 52021
rect 8539 51965 8595 52021
rect 8681 51965 8737 52021
rect 8823 51965 8879 52021
rect 8965 51965 9021 52021
rect 9107 51965 9163 52021
rect 9249 51965 9305 52021
rect 9391 51965 9447 52021
rect 9533 51965 9589 52021
rect 9675 51965 9731 52021
rect 9817 51965 9873 52021
rect 9959 51965 10015 52021
rect 10101 51965 10157 52021
rect 10243 51965 10299 52021
rect 10385 51965 10441 52021
rect 10527 51965 10583 52021
rect 10669 51965 10725 52021
rect 10811 51965 10867 52021
rect 10953 51965 11009 52021
rect 11095 51965 11151 52021
rect 11237 51965 11293 52021
rect 11379 51965 11435 52021
rect 11521 51965 11577 52021
rect 11663 51965 11719 52021
rect 11805 51965 11861 52021
rect 11947 51965 12003 52021
rect 12089 51965 12145 52021
rect 12231 51965 12287 52021
rect 12373 51965 12429 52021
rect 12515 51965 12571 52021
rect 12657 51965 12713 52021
rect 12799 51965 12855 52021
rect 12941 51965 12997 52021
rect 13083 51965 13139 52021
rect 13225 51965 13281 52021
rect 13367 51965 13423 52021
rect 13509 51965 13565 52021
rect 13651 51965 13707 52021
rect 13793 51965 13849 52021
rect 13935 51965 13991 52021
rect 14077 51965 14133 52021
rect 14219 51965 14275 52021
rect 14361 51965 14417 52021
rect 14503 51965 14559 52021
rect 14645 51965 14701 52021
rect 14787 51965 14843 52021
rect 161 51823 217 51879
rect 303 51823 359 51879
rect 445 51823 501 51879
rect 587 51823 643 51879
rect 729 51823 785 51879
rect 871 51823 927 51879
rect 1013 51823 1069 51879
rect 1155 51823 1211 51879
rect 1297 51823 1353 51879
rect 1439 51823 1495 51879
rect 1581 51823 1637 51879
rect 1723 51823 1779 51879
rect 1865 51823 1921 51879
rect 2007 51823 2063 51879
rect 2149 51823 2205 51879
rect 2291 51823 2347 51879
rect 2433 51823 2489 51879
rect 2575 51823 2631 51879
rect 2717 51823 2773 51879
rect 2859 51823 2915 51879
rect 3001 51823 3057 51879
rect 3143 51823 3199 51879
rect 3285 51823 3341 51879
rect 3427 51823 3483 51879
rect 3569 51823 3625 51879
rect 3711 51823 3767 51879
rect 3853 51823 3909 51879
rect 3995 51823 4051 51879
rect 4137 51823 4193 51879
rect 4279 51823 4335 51879
rect 4421 51823 4477 51879
rect 4563 51823 4619 51879
rect 4705 51823 4761 51879
rect 4847 51823 4903 51879
rect 4989 51823 5045 51879
rect 5131 51823 5187 51879
rect 5273 51823 5329 51879
rect 5415 51823 5471 51879
rect 5557 51823 5613 51879
rect 5699 51823 5755 51879
rect 5841 51823 5897 51879
rect 5983 51823 6039 51879
rect 6125 51823 6181 51879
rect 6267 51823 6323 51879
rect 6409 51823 6465 51879
rect 6551 51823 6607 51879
rect 6693 51823 6749 51879
rect 6835 51823 6891 51879
rect 6977 51823 7033 51879
rect 7119 51823 7175 51879
rect 7261 51823 7317 51879
rect 7403 51823 7459 51879
rect 7545 51823 7601 51879
rect 7687 51823 7743 51879
rect 7829 51823 7885 51879
rect 7971 51823 8027 51879
rect 8113 51823 8169 51879
rect 8255 51823 8311 51879
rect 8397 51823 8453 51879
rect 8539 51823 8595 51879
rect 8681 51823 8737 51879
rect 8823 51823 8879 51879
rect 8965 51823 9021 51879
rect 9107 51823 9163 51879
rect 9249 51823 9305 51879
rect 9391 51823 9447 51879
rect 9533 51823 9589 51879
rect 9675 51823 9731 51879
rect 9817 51823 9873 51879
rect 9959 51823 10015 51879
rect 10101 51823 10157 51879
rect 10243 51823 10299 51879
rect 10385 51823 10441 51879
rect 10527 51823 10583 51879
rect 10669 51823 10725 51879
rect 10811 51823 10867 51879
rect 10953 51823 11009 51879
rect 11095 51823 11151 51879
rect 11237 51823 11293 51879
rect 11379 51823 11435 51879
rect 11521 51823 11577 51879
rect 11663 51823 11719 51879
rect 11805 51823 11861 51879
rect 11947 51823 12003 51879
rect 12089 51823 12145 51879
rect 12231 51823 12287 51879
rect 12373 51823 12429 51879
rect 12515 51823 12571 51879
rect 12657 51823 12713 51879
rect 12799 51823 12855 51879
rect 12941 51823 12997 51879
rect 13083 51823 13139 51879
rect 13225 51823 13281 51879
rect 13367 51823 13423 51879
rect 13509 51823 13565 51879
rect 13651 51823 13707 51879
rect 13793 51823 13849 51879
rect 13935 51823 13991 51879
rect 14077 51823 14133 51879
rect 14219 51823 14275 51879
rect 14361 51823 14417 51879
rect 14503 51823 14559 51879
rect 14645 51823 14701 51879
rect 14787 51823 14843 51879
rect 161 51681 217 51737
rect 303 51681 359 51737
rect 445 51681 501 51737
rect 587 51681 643 51737
rect 729 51681 785 51737
rect 871 51681 927 51737
rect 1013 51681 1069 51737
rect 1155 51681 1211 51737
rect 1297 51681 1353 51737
rect 1439 51681 1495 51737
rect 1581 51681 1637 51737
rect 1723 51681 1779 51737
rect 1865 51681 1921 51737
rect 2007 51681 2063 51737
rect 2149 51681 2205 51737
rect 2291 51681 2347 51737
rect 2433 51681 2489 51737
rect 2575 51681 2631 51737
rect 2717 51681 2773 51737
rect 2859 51681 2915 51737
rect 3001 51681 3057 51737
rect 3143 51681 3199 51737
rect 3285 51681 3341 51737
rect 3427 51681 3483 51737
rect 3569 51681 3625 51737
rect 3711 51681 3767 51737
rect 3853 51681 3909 51737
rect 3995 51681 4051 51737
rect 4137 51681 4193 51737
rect 4279 51681 4335 51737
rect 4421 51681 4477 51737
rect 4563 51681 4619 51737
rect 4705 51681 4761 51737
rect 4847 51681 4903 51737
rect 4989 51681 5045 51737
rect 5131 51681 5187 51737
rect 5273 51681 5329 51737
rect 5415 51681 5471 51737
rect 5557 51681 5613 51737
rect 5699 51681 5755 51737
rect 5841 51681 5897 51737
rect 5983 51681 6039 51737
rect 6125 51681 6181 51737
rect 6267 51681 6323 51737
rect 6409 51681 6465 51737
rect 6551 51681 6607 51737
rect 6693 51681 6749 51737
rect 6835 51681 6891 51737
rect 6977 51681 7033 51737
rect 7119 51681 7175 51737
rect 7261 51681 7317 51737
rect 7403 51681 7459 51737
rect 7545 51681 7601 51737
rect 7687 51681 7743 51737
rect 7829 51681 7885 51737
rect 7971 51681 8027 51737
rect 8113 51681 8169 51737
rect 8255 51681 8311 51737
rect 8397 51681 8453 51737
rect 8539 51681 8595 51737
rect 8681 51681 8737 51737
rect 8823 51681 8879 51737
rect 8965 51681 9021 51737
rect 9107 51681 9163 51737
rect 9249 51681 9305 51737
rect 9391 51681 9447 51737
rect 9533 51681 9589 51737
rect 9675 51681 9731 51737
rect 9817 51681 9873 51737
rect 9959 51681 10015 51737
rect 10101 51681 10157 51737
rect 10243 51681 10299 51737
rect 10385 51681 10441 51737
rect 10527 51681 10583 51737
rect 10669 51681 10725 51737
rect 10811 51681 10867 51737
rect 10953 51681 11009 51737
rect 11095 51681 11151 51737
rect 11237 51681 11293 51737
rect 11379 51681 11435 51737
rect 11521 51681 11577 51737
rect 11663 51681 11719 51737
rect 11805 51681 11861 51737
rect 11947 51681 12003 51737
rect 12089 51681 12145 51737
rect 12231 51681 12287 51737
rect 12373 51681 12429 51737
rect 12515 51681 12571 51737
rect 12657 51681 12713 51737
rect 12799 51681 12855 51737
rect 12941 51681 12997 51737
rect 13083 51681 13139 51737
rect 13225 51681 13281 51737
rect 13367 51681 13423 51737
rect 13509 51681 13565 51737
rect 13651 51681 13707 51737
rect 13793 51681 13849 51737
rect 13935 51681 13991 51737
rect 14077 51681 14133 51737
rect 14219 51681 14275 51737
rect 14361 51681 14417 51737
rect 14503 51681 14559 51737
rect 14645 51681 14701 51737
rect 14787 51681 14843 51737
rect 161 51539 217 51595
rect 303 51539 359 51595
rect 445 51539 501 51595
rect 587 51539 643 51595
rect 729 51539 785 51595
rect 871 51539 927 51595
rect 1013 51539 1069 51595
rect 1155 51539 1211 51595
rect 1297 51539 1353 51595
rect 1439 51539 1495 51595
rect 1581 51539 1637 51595
rect 1723 51539 1779 51595
rect 1865 51539 1921 51595
rect 2007 51539 2063 51595
rect 2149 51539 2205 51595
rect 2291 51539 2347 51595
rect 2433 51539 2489 51595
rect 2575 51539 2631 51595
rect 2717 51539 2773 51595
rect 2859 51539 2915 51595
rect 3001 51539 3057 51595
rect 3143 51539 3199 51595
rect 3285 51539 3341 51595
rect 3427 51539 3483 51595
rect 3569 51539 3625 51595
rect 3711 51539 3767 51595
rect 3853 51539 3909 51595
rect 3995 51539 4051 51595
rect 4137 51539 4193 51595
rect 4279 51539 4335 51595
rect 4421 51539 4477 51595
rect 4563 51539 4619 51595
rect 4705 51539 4761 51595
rect 4847 51539 4903 51595
rect 4989 51539 5045 51595
rect 5131 51539 5187 51595
rect 5273 51539 5329 51595
rect 5415 51539 5471 51595
rect 5557 51539 5613 51595
rect 5699 51539 5755 51595
rect 5841 51539 5897 51595
rect 5983 51539 6039 51595
rect 6125 51539 6181 51595
rect 6267 51539 6323 51595
rect 6409 51539 6465 51595
rect 6551 51539 6607 51595
rect 6693 51539 6749 51595
rect 6835 51539 6891 51595
rect 6977 51539 7033 51595
rect 7119 51539 7175 51595
rect 7261 51539 7317 51595
rect 7403 51539 7459 51595
rect 7545 51539 7601 51595
rect 7687 51539 7743 51595
rect 7829 51539 7885 51595
rect 7971 51539 8027 51595
rect 8113 51539 8169 51595
rect 8255 51539 8311 51595
rect 8397 51539 8453 51595
rect 8539 51539 8595 51595
rect 8681 51539 8737 51595
rect 8823 51539 8879 51595
rect 8965 51539 9021 51595
rect 9107 51539 9163 51595
rect 9249 51539 9305 51595
rect 9391 51539 9447 51595
rect 9533 51539 9589 51595
rect 9675 51539 9731 51595
rect 9817 51539 9873 51595
rect 9959 51539 10015 51595
rect 10101 51539 10157 51595
rect 10243 51539 10299 51595
rect 10385 51539 10441 51595
rect 10527 51539 10583 51595
rect 10669 51539 10725 51595
rect 10811 51539 10867 51595
rect 10953 51539 11009 51595
rect 11095 51539 11151 51595
rect 11237 51539 11293 51595
rect 11379 51539 11435 51595
rect 11521 51539 11577 51595
rect 11663 51539 11719 51595
rect 11805 51539 11861 51595
rect 11947 51539 12003 51595
rect 12089 51539 12145 51595
rect 12231 51539 12287 51595
rect 12373 51539 12429 51595
rect 12515 51539 12571 51595
rect 12657 51539 12713 51595
rect 12799 51539 12855 51595
rect 12941 51539 12997 51595
rect 13083 51539 13139 51595
rect 13225 51539 13281 51595
rect 13367 51539 13423 51595
rect 13509 51539 13565 51595
rect 13651 51539 13707 51595
rect 13793 51539 13849 51595
rect 13935 51539 13991 51595
rect 14077 51539 14133 51595
rect 14219 51539 14275 51595
rect 14361 51539 14417 51595
rect 14503 51539 14559 51595
rect 14645 51539 14701 51595
rect 14787 51539 14843 51595
rect 161 51397 217 51453
rect 303 51397 359 51453
rect 445 51397 501 51453
rect 587 51397 643 51453
rect 729 51397 785 51453
rect 871 51397 927 51453
rect 1013 51397 1069 51453
rect 1155 51397 1211 51453
rect 1297 51397 1353 51453
rect 1439 51397 1495 51453
rect 1581 51397 1637 51453
rect 1723 51397 1779 51453
rect 1865 51397 1921 51453
rect 2007 51397 2063 51453
rect 2149 51397 2205 51453
rect 2291 51397 2347 51453
rect 2433 51397 2489 51453
rect 2575 51397 2631 51453
rect 2717 51397 2773 51453
rect 2859 51397 2915 51453
rect 3001 51397 3057 51453
rect 3143 51397 3199 51453
rect 3285 51397 3341 51453
rect 3427 51397 3483 51453
rect 3569 51397 3625 51453
rect 3711 51397 3767 51453
rect 3853 51397 3909 51453
rect 3995 51397 4051 51453
rect 4137 51397 4193 51453
rect 4279 51397 4335 51453
rect 4421 51397 4477 51453
rect 4563 51397 4619 51453
rect 4705 51397 4761 51453
rect 4847 51397 4903 51453
rect 4989 51397 5045 51453
rect 5131 51397 5187 51453
rect 5273 51397 5329 51453
rect 5415 51397 5471 51453
rect 5557 51397 5613 51453
rect 5699 51397 5755 51453
rect 5841 51397 5897 51453
rect 5983 51397 6039 51453
rect 6125 51397 6181 51453
rect 6267 51397 6323 51453
rect 6409 51397 6465 51453
rect 6551 51397 6607 51453
rect 6693 51397 6749 51453
rect 6835 51397 6891 51453
rect 6977 51397 7033 51453
rect 7119 51397 7175 51453
rect 7261 51397 7317 51453
rect 7403 51397 7459 51453
rect 7545 51397 7601 51453
rect 7687 51397 7743 51453
rect 7829 51397 7885 51453
rect 7971 51397 8027 51453
rect 8113 51397 8169 51453
rect 8255 51397 8311 51453
rect 8397 51397 8453 51453
rect 8539 51397 8595 51453
rect 8681 51397 8737 51453
rect 8823 51397 8879 51453
rect 8965 51397 9021 51453
rect 9107 51397 9163 51453
rect 9249 51397 9305 51453
rect 9391 51397 9447 51453
rect 9533 51397 9589 51453
rect 9675 51397 9731 51453
rect 9817 51397 9873 51453
rect 9959 51397 10015 51453
rect 10101 51397 10157 51453
rect 10243 51397 10299 51453
rect 10385 51397 10441 51453
rect 10527 51397 10583 51453
rect 10669 51397 10725 51453
rect 10811 51397 10867 51453
rect 10953 51397 11009 51453
rect 11095 51397 11151 51453
rect 11237 51397 11293 51453
rect 11379 51397 11435 51453
rect 11521 51397 11577 51453
rect 11663 51397 11719 51453
rect 11805 51397 11861 51453
rect 11947 51397 12003 51453
rect 12089 51397 12145 51453
rect 12231 51397 12287 51453
rect 12373 51397 12429 51453
rect 12515 51397 12571 51453
rect 12657 51397 12713 51453
rect 12799 51397 12855 51453
rect 12941 51397 12997 51453
rect 13083 51397 13139 51453
rect 13225 51397 13281 51453
rect 13367 51397 13423 51453
rect 13509 51397 13565 51453
rect 13651 51397 13707 51453
rect 13793 51397 13849 51453
rect 13935 51397 13991 51453
rect 14077 51397 14133 51453
rect 14219 51397 14275 51453
rect 14361 51397 14417 51453
rect 14503 51397 14559 51453
rect 14645 51397 14701 51453
rect 14787 51397 14843 51453
rect 161 51255 217 51311
rect 303 51255 359 51311
rect 445 51255 501 51311
rect 587 51255 643 51311
rect 729 51255 785 51311
rect 871 51255 927 51311
rect 1013 51255 1069 51311
rect 1155 51255 1211 51311
rect 1297 51255 1353 51311
rect 1439 51255 1495 51311
rect 1581 51255 1637 51311
rect 1723 51255 1779 51311
rect 1865 51255 1921 51311
rect 2007 51255 2063 51311
rect 2149 51255 2205 51311
rect 2291 51255 2347 51311
rect 2433 51255 2489 51311
rect 2575 51255 2631 51311
rect 2717 51255 2773 51311
rect 2859 51255 2915 51311
rect 3001 51255 3057 51311
rect 3143 51255 3199 51311
rect 3285 51255 3341 51311
rect 3427 51255 3483 51311
rect 3569 51255 3625 51311
rect 3711 51255 3767 51311
rect 3853 51255 3909 51311
rect 3995 51255 4051 51311
rect 4137 51255 4193 51311
rect 4279 51255 4335 51311
rect 4421 51255 4477 51311
rect 4563 51255 4619 51311
rect 4705 51255 4761 51311
rect 4847 51255 4903 51311
rect 4989 51255 5045 51311
rect 5131 51255 5187 51311
rect 5273 51255 5329 51311
rect 5415 51255 5471 51311
rect 5557 51255 5613 51311
rect 5699 51255 5755 51311
rect 5841 51255 5897 51311
rect 5983 51255 6039 51311
rect 6125 51255 6181 51311
rect 6267 51255 6323 51311
rect 6409 51255 6465 51311
rect 6551 51255 6607 51311
rect 6693 51255 6749 51311
rect 6835 51255 6891 51311
rect 6977 51255 7033 51311
rect 7119 51255 7175 51311
rect 7261 51255 7317 51311
rect 7403 51255 7459 51311
rect 7545 51255 7601 51311
rect 7687 51255 7743 51311
rect 7829 51255 7885 51311
rect 7971 51255 8027 51311
rect 8113 51255 8169 51311
rect 8255 51255 8311 51311
rect 8397 51255 8453 51311
rect 8539 51255 8595 51311
rect 8681 51255 8737 51311
rect 8823 51255 8879 51311
rect 8965 51255 9021 51311
rect 9107 51255 9163 51311
rect 9249 51255 9305 51311
rect 9391 51255 9447 51311
rect 9533 51255 9589 51311
rect 9675 51255 9731 51311
rect 9817 51255 9873 51311
rect 9959 51255 10015 51311
rect 10101 51255 10157 51311
rect 10243 51255 10299 51311
rect 10385 51255 10441 51311
rect 10527 51255 10583 51311
rect 10669 51255 10725 51311
rect 10811 51255 10867 51311
rect 10953 51255 11009 51311
rect 11095 51255 11151 51311
rect 11237 51255 11293 51311
rect 11379 51255 11435 51311
rect 11521 51255 11577 51311
rect 11663 51255 11719 51311
rect 11805 51255 11861 51311
rect 11947 51255 12003 51311
rect 12089 51255 12145 51311
rect 12231 51255 12287 51311
rect 12373 51255 12429 51311
rect 12515 51255 12571 51311
rect 12657 51255 12713 51311
rect 12799 51255 12855 51311
rect 12941 51255 12997 51311
rect 13083 51255 13139 51311
rect 13225 51255 13281 51311
rect 13367 51255 13423 51311
rect 13509 51255 13565 51311
rect 13651 51255 13707 51311
rect 13793 51255 13849 51311
rect 13935 51255 13991 51311
rect 14077 51255 14133 51311
rect 14219 51255 14275 51311
rect 14361 51255 14417 51311
rect 14503 51255 14559 51311
rect 14645 51255 14701 51311
rect 14787 51255 14843 51311
rect 161 51113 217 51169
rect 303 51113 359 51169
rect 445 51113 501 51169
rect 587 51113 643 51169
rect 729 51113 785 51169
rect 871 51113 927 51169
rect 1013 51113 1069 51169
rect 1155 51113 1211 51169
rect 1297 51113 1353 51169
rect 1439 51113 1495 51169
rect 1581 51113 1637 51169
rect 1723 51113 1779 51169
rect 1865 51113 1921 51169
rect 2007 51113 2063 51169
rect 2149 51113 2205 51169
rect 2291 51113 2347 51169
rect 2433 51113 2489 51169
rect 2575 51113 2631 51169
rect 2717 51113 2773 51169
rect 2859 51113 2915 51169
rect 3001 51113 3057 51169
rect 3143 51113 3199 51169
rect 3285 51113 3341 51169
rect 3427 51113 3483 51169
rect 3569 51113 3625 51169
rect 3711 51113 3767 51169
rect 3853 51113 3909 51169
rect 3995 51113 4051 51169
rect 4137 51113 4193 51169
rect 4279 51113 4335 51169
rect 4421 51113 4477 51169
rect 4563 51113 4619 51169
rect 4705 51113 4761 51169
rect 4847 51113 4903 51169
rect 4989 51113 5045 51169
rect 5131 51113 5187 51169
rect 5273 51113 5329 51169
rect 5415 51113 5471 51169
rect 5557 51113 5613 51169
rect 5699 51113 5755 51169
rect 5841 51113 5897 51169
rect 5983 51113 6039 51169
rect 6125 51113 6181 51169
rect 6267 51113 6323 51169
rect 6409 51113 6465 51169
rect 6551 51113 6607 51169
rect 6693 51113 6749 51169
rect 6835 51113 6891 51169
rect 6977 51113 7033 51169
rect 7119 51113 7175 51169
rect 7261 51113 7317 51169
rect 7403 51113 7459 51169
rect 7545 51113 7601 51169
rect 7687 51113 7743 51169
rect 7829 51113 7885 51169
rect 7971 51113 8027 51169
rect 8113 51113 8169 51169
rect 8255 51113 8311 51169
rect 8397 51113 8453 51169
rect 8539 51113 8595 51169
rect 8681 51113 8737 51169
rect 8823 51113 8879 51169
rect 8965 51113 9021 51169
rect 9107 51113 9163 51169
rect 9249 51113 9305 51169
rect 9391 51113 9447 51169
rect 9533 51113 9589 51169
rect 9675 51113 9731 51169
rect 9817 51113 9873 51169
rect 9959 51113 10015 51169
rect 10101 51113 10157 51169
rect 10243 51113 10299 51169
rect 10385 51113 10441 51169
rect 10527 51113 10583 51169
rect 10669 51113 10725 51169
rect 10811 51113 10867 51169
rect 10953 51113 11009 51169
rect 11095 51113 11151 51169
rect 11237 51113 11293 51169
rect 11379 51113 11435 51169
rect 11521 51113 11577 51169
rect 11663 51113 11719 51169
rect 11805 51113 11861 51169
rect 11947 51113 12003 51169
rect 12089 51113 12145 51169
rect 12231 51113 12287 51169
rect 12373 51113 12429 51169
rect 12515 51113 12571 51169
rect 12657 51113 12713 51169
rect 12799 51113 12855 51169
rect 12941 51113 12997 51169
rect 13083 51113 13139 51169
rect 13225 51113 13281 51169
rect 13367 51113 13423 51169
rect 13509 51113 13565 51169
rect 13651 51113 13707 51169
rect 13793 51113 13849 51169
rect 13935 51113 13991 51169
rect 14077 51113 14133 51169
rect 14219 51113 14275 51169
rect 14361 51113 14417 51169
rect 14503 51113 14559 51169
rect 14645 51113 14701 51169
rect 14787 51113 14843 51169
rect 161 50971 217 51027
rect 303 50971 359 51027
rect 445 50971 501 51027
rect 587 50971 643 51027
rect 729 50971 785 51027
rect 871 50971 927 51027
rect 1013 50971 1069 51027
rect 1155 50971 1211 51027
rect 1297 50971 1353 51027
rect 1439 50971 1495 51027
rect 1581 50971 1637 51027
rect 1723 50971 1779 51027
rect 1865 50971 1921 51027
rect 2007 50971 2063 51027
rect 2149 50971 2205 51027
rect 2291 50971 2347 51027
rect 2433 50971 2489 51027
rect 2575 50971 2631 51027
rect 2717 50971 2773 51027
rect 2859 50971 2915 51027
rect 3001 50971 3057 51027
rect 3143 50971 3199 51027
rect 3285 50971 3341 51027
rect 3427 50971 3483 51027
rect 3569 50971 3625 51027
rect 3711 50971 3767 51027
rect 3853 50971 3909 51027
rect 3995 50971 4051 51027
rect 4137 50971 4193 51027
rect 4279 50971 4335 51027
rect 4421 50971 4477 51027
rect 4563 50971 4619 51027
rect 4705 50971 4761 51027
rect 4847 50971 4903 51027
rect 4989 50971 5045 51027
rect 5131 50971 5187 51027
rect 5273 50971 5329 51027
rect 5415 50971 5471 51027
rect 5557 50971 5613 51027
rect 5699 50971 5755 51027
rect 5841 50971 5897 51027
rect 5983 50971 6039 51027
rect 6125 50971 6181 51027
rect 6267 50971 6323 51027
rect 6409 50971 6465 51027
rect 6551 50971 6607 51027
rect 6693 50971 6749 51027
rect 6835 50971 6891 51027
rect 6977 50971 7033 51027
rect 7119 50971 7175 51027
rect 7261 50971 7317 51027
rect 7403 50971 7459 51027
rect 7545 50971 7601 51027
rect 7687 50971 7743 51027
rect 7829 50971 7885 51027
rect 7971 50971 8027 51027
rect 8113 50971 8169 51027
rect 8255 50971 8311 51027
rect 8397 50971 8453 51027
rect 8539 50971 8595 51027
rect 8681 50971 8737 51027
rect 8823 50971 8879 51027
rect 8965 50971 9021 51027
rect 9107 50971 9163 51027
rect 9249 50971 9305 51027
rect 9391 50971 9447 51027
rect 9533 50971 9589 51027
rect 9675 50971 9731 51027
rect 9817 50971 9873 51027
rect 9959 50971 10015 51027
rect 10101 50971 10157 51027
rect 10243 50971 10299 51027
rect 10385 50971 10441 51027
rect 10527 50971 10583 51027
rect 10669 50971 10725 51027
rect 10811 50971 10867 51027
rect 10953 50971 11009 51027
rect 11095 50971 11151 51027
rect 11237 50971 11293 51027
rect 11379 50971 11435 51027
rect 11521 50971 11577 51027
rect 11663 50971 11719 51027
rect 11805 50971 11861 51027
rect 11947 50971 12003 51027
rect 12089 50971 12145 51027
rect 12231 50971 12287 51027
rect 12373 50971 12429 51027
rect 12515 50971 12571 51027
rect 12657 50971 12713 51027
rect 12799 50971 12855 51027
rect 12941 50971 12997 51027
rect 13083 50971 13139 51027
rect 13225 50971 13281 51027
rect 13367 50971 13423 51027
rect 13509 50971 13565 51027
rect 13651 50971 13707 51027
rect 13793 50971 13849 51027
rect 13935 50971 13991 51027
rect 14077 50971 14133 51027
rect 14219 50971 14275 51027
rect 14361 50971 14417 51027
rect 14503 50971 14559 51027
rect 14645 50971 14701 51027
rect 14787 50971 14843 51027
rect 161 50829 217 50885
rect 303 50829 359 50885
rect 445 50829 501 50885
rect 587 50829 643 50885
rect 729 50829 785 50885
rect 871 50829 927 50885
rect 1013 50829 1069 50885
rect 1155 50829 1211 50885
rect 1297 50829 1353 50885
rect 1439 50829 1495 50885
rect 1581 50829 1637 50885
rect 1723 50829 1779 50885
rect 1865 50829 1921 50885
rect 2007 50829 2063 50885
rect 2149 50829 2205 50885
rect 2291 50829 2347 50885
rect 2433 50829 2489 50885
rect 2575 50829 2631 50885
rect 2717 50829 2773 50885
rect 2859 50829 2915 50885
rect 3001 50829 3057 50885
rect 3143 50829 3199 50885
rect 3285 50829 3341 50885
rect 3427 50829 3483 50885
rect 3569 50829 3625 50885
rect 3711 50829 3767 50885
rect 3853 50829 3909 50885
rect 3995 50829 4051 50885
rect 4137 50829 4193 50885
rect 4279 50829 4335 50885
rect 4421 50829 4477 50885
rect 4563 50829 4619 50885
rect 4705 50829 4761 50885
rect 4847 50829 4903 50885
rect 4989 50829 5045 50885
rect 5131 50829 5187 50885
rect 5273 50829 5329 50885
rect 5415 50829 5471 50885
rect 5557 50829 5613 50885
rect 5699 50829 5755 50885
rect 5841 50829 5897 50885
rect 5983 50829 6039 50885
rect 6125 50829 6181 50885
rect 6267 50829 6323 50885
rect 6409 50829 6465 50885
rect 6551 50829 6607 50885
rect 6693 50829 6749 50885
rect 6835 50829 6891 50885
rect 6977 50829 7033 50885
rect 7119 50829 7175 50885
rect 7261 50829 7317 50885
rect 7403 50829 7459 50885
rect 7545 50829 7601 50885
rect 7687 50829 7743 50885
rect 7829 50829 7885 50885
rect 7971 50829 8027 50885
rect 8113 50829 8169 50885
rect 8255 50829 8311 50885
rect 8397 50829 8453 50885
rect 8539 50829 8595 50885
rect 8681 50829 8737 50885
rect 8823 50829 8879 50885
rect 8965 50829 9021 50885
rect 9107 50829 9163 50885
rect 9249 50829 9305 50885
rect 9391 50829 9447 50885
rect 9533 50829 9589 50885
rect 9675 50829 9731 50885
rect 9817 50829 9873 50885
rect 9959 50829 10015 50885
rect 10101 50829 10157 50885
rect 10243 50829 10299 50885
rect 10385 50829 10441 50885
rect 10527 50829 10583 50885
rect 10669 50829 10725 50885
rect 10811 50829 10867 50885
rect 10953 50829 11009 50885
rect 11095 50829 11151 50885
rect 11237 50829 11293 50885
rect 11379 50829 11435 50885
rect 11521 50829 11577 50885
rect 11663 50829 11719 50885
rect 11805 50829 11861 50885
rect 11947 50829 12003 50885
rect 12089 50829 12145 50885
rect 12231 50829 12287 50885
rect 12373 50829 12429 50885
rect 12515 50829 12571 50885
rect 12657 50829 12713 50885
rect 12799 50829 12855 50885
rect 12941 50829 12997 50885
rect 13083 50829 13139 50885
rect 13225 50829 13281 50885
rect 13367 50829 13423 50885
rect 13509 50829 13565 50885
rect 13651 50829 13707 50885
rect 13793 50829 13849 50885
rect 13935 50829 13991 50885
rect 14077 50829 14133 50885
rect 14219 50829 14275 50885
rect 14361 50829 14417 50885
rect 14503 50829 14559 50885
rect 14645 50829 14701 50885
rect 14787 50829 14843 50885
rect 161 50507 217 50563
rect 303 50507 359 50563
rect 445 50507 501 50563
rect 587 50507 643 50563
rect 729 50507 785 50563
rect 871 50507 927 50563
rect 1013 50507 1069 50563
rect 1155 50507 1211 50563
rect 1297 50507 1353 50563
rect 1439 50507 1495 50563
rect 1581 50507 1637 50563
rect 1723 50507 1779 50563
rect 1865 50507 1921 50563
rect 2007 50507 2063 50563
rect 2149 50507 2205 50563
rect 2291 50507 2347 50563
rect 2433 50507 2489 50563
rect 2575 50507 2631 50563
rect 2717 50507 2773 50563
rect 2859 50507 2915 50563
rect 3001 50507 3057 50563
rect 3143 50507 3199 50563
rect 3285 50507 3341 50563
rect 3427 50507 3483 50563
rect 3569 50507 3625 50563
rect 3711 50507 3767 50563
rect 3853 50507 3909 50563
rect 3995 50507 4051 50563
rect 4137 50507 4193 50563
rect 4279 50507 4335 50563
rect 4421 50507 4477 50563
rect 4563 50507 4619 50563
rect 4705 50507 4761 50563
rect 4847 50507 4903 50563
rect 4989 50507 5045 50563
rect 5131 50507 5187 50563
rect 5273 50507 5329 50563
rect 5415 50507 5471 50563
rect 5557 50507 5613 50563
rect 5699 50507 5755 50563
rect 5841 50507 5897 50563
rect 5983 50507 6039 50563
rect 6125 50507 6181 50563
rect 6267 50507 6323 50563
rect 6409 50507 6465 50563
rect 6551 50507 6607 50563
rect 6693 50507 6749 50563
rect 6835 50507 6891 50563
rect 6977 50507 7033 50563
rect 7119 50507 7175 50563
rect 7261 50507 7317 50563
rect 7403 50507 7459 50563
rect 7545 50507 7601 50563
rect 7687 50507 7743 50563
rect 7829 50507 7885 50563
rect 7971 50507 8027 50563
rect 8113 50507 8169 50563
rect 8255 50507 8311 50563
rect 8397 50507 8453 50563
rect 8539 50507 8595 50563
rect 8681 50507 8737 50563
rect 8823 50507 8879 50563
rect 8965 50507 9021 50563
rect 9107 50507 9163 50563
rect 9249 50507 9305 50563
rect 9391 50507 9447 50563
rect 9533 50507 9589 50563
rect 9675 50507 9731 50563
rect 9817 50507 9873 50563
rect 9959 50507 10015 50563
rect 10101 50507 10157 50563
rect 10243 50507 10299 50563
rect 10385 50507 10441 50563
rect 10527 50507 10583 50563
rect 10669 50507 10725 50563
rect 10811 50507 10867 50563
rect 10953 50507 11009 50563
rect 11095 50507 11151 50563
rect 11237 50507 11293 50563
rect 11379 50507 11435 50563
rect 11521 50507 11577 50563
rect 11663 50507 11719 50563
rect 11805 50507 11861 50563
rect 11947 50507 12003 50563
rect 12089 50507 12145 50563
rect 12231 50507 12287 50563
rect 12373 50507 12429 50563
rect 12515 50507 12571 50563
rect 12657 50507 12713 50563
rect 12799 50507 12855 50563
rect 12941 50507 12997 50563
rect 13083 50507 13139 50563
rect 13225 50507 13281 50563
rect 13367 50507 13423 50563
rect 13509 50507 13565 50563
rect 13651 50507 13707 50563
rect 13793 50507 13849 50563
rect 13935 50507 13991 50563
rect 14077 50507 14133 50563
rect 14219 50507 14275 50563
rect 14361 50507 14417 50563
rect 14503 50507 14559 50563
rect 14645 50507 14701 50563
rect 14787 50507 14843 50563
rect 161 50365 217 50421
rect 303 50365 359 50421
rect 445 50365 501 50421
rect 587 50365 643 50421
rect 729 50365 785 50421
rect 871 50365 927 50421
rect 1013 50365 1069 50421
rect 1155 50365 1211 50421
rect 1297 50365 1353 50421
rect 1439 50365 1495 50421
rect 1581 50365 1637 50421
rect 1723 50365 1779 50421
rect 1865 50365 1921 50421
rect 2007 50365 2063 50421
rect 2149 50365 2205 50421
rect 2291 50365 2347 50421
rect 2433 50365 2489 50421
rect 2575 50365 2631 50421
rect 2717 50365 2773 50421
rect 2859 50365 2915 50421
rect 3001 50365 3057 50421
rect 3143 50365 3199 50421
rect 3285 50365 3341 50421
rect 3427 50365 3483 50421
rect 3569 50365 3625 50421
rect 3711 50365 3767 50421
rect 3853 50365 3909 50421
rect 3995 50365 4051 50421
rect 4137 50365 4193 50421
rect 4279 50365 4335 50421
rect 4421 50365 4477 50421
rect 4563 50365 4619 50421
rect 4705 50365 4761 50421
rect 4847 50365 4903 50421
rect 4989 50365 5045 50421
rect 5131 50365 5187 50421
rect 5273 50365 5329 50421
rect 5415 50365 5471 50421
rect 5557 50365 5613 50421
rect 5699 50365 5755 50421
rect 5841 50365 5897 50421
rect 5983 50365 6039 50421
rect 6125 50365 6181 50421
rect 6267 50365 6323 50421
rect 6409 50365 6465 50421
rect 6551 50365 6607 50421
rect 6693 50365 6749 50421
rect 6835 50365 6891 50421
rect 6977 50365 7033 50421
rect 7119 50365 7175 50421
rect 7261 50365 7317 50421
rect 7403 50365 7459 50421
rect 7545 50365 7601 50421
rect 7687 50365 7743 50421
rect 7829 50365 7885 50421
rect 7971 50365 8027 50421
rect 8113 50365 8169 50421
rect 8255 50365 8311 50421
rect 8397 50365 8453 50421
rect 8539 50365 8595 50421
rect 8681 50365 8737 50421
rect 8823 50365 8879 50421
rect 8965 50365 9021 50421
rect 9107 50365 9163 50421
rect 9249 50365 9305 50421
rect 9391 50365 9447 50421
rect 9533 50365 9589 50421
rect 9675 50365 9731 50421
rect 9817 50365 9873 50421
rect 9959 50365 10015 50421
rect 10101 50365 10157 50421
rect 10243 50365 10299 50421
rect 10385 50365 10441 50421
rect 10527 50365 10583 50421
rect 10669 50365 10725 50421
rect 10811 50365 10867 50421
rect 10953 50365 11009 50421
rect 11095 50365 11151 50421
rect 11237 50365 11293 50421
rect 11379 50365 11435 50421
rect 11521 50365 11577 50421
rect 11663 50365 11719 50421
rect 11805 50365 11861 50421
rect 11947 50365 12003 50421
rect 12089 50365 12145 50421
rect 12231 50365 12287 50421
rect 12373 50365 12429 50421
rect 12515 50365 12571 50421
rect 12657 50365 12713 50421
rect 12799 50365 12855 50421
rect 12941 50365 12997 50421
rect 13083 50365 13139 50421
rect 13225 50365 13281 50421
rect 13367 50365 13423 50421
rect 13509 50365 13565 50421
rect 13651 50365 13707 50421
rect 13793 50365 13849 50421
rect 13935 50365 13991 50421
rect 14077 50365 14133 50421
rect 14219 50365 14275 50421
rect 14361 50365 14417 50421
rect 14503 50365 14559 50421
rect 14645 50365 14701 50421
rect 14787 50365 14843 50421
rect 161 50223 217 50279
rect 303 50223 359 50279
rect 445 50223 501 50279
rect 587 50223 643 50279
rect 729 50223 785 50279
rect 871 50223 927 50279
rect 1013 50223 1069 50279
rect 1155 50223 1211 50279
rect 1297 50223 1353 50279
rect 1439 50223 1495 50279
rect 1581 50223 1637 50279
rect 1723 50223 1779 50279
rect 1865 50223 1921 50279
rect 2007 50223 2063 50279
rect 2149 50223 2205 50279
rect 2291 50223 2347 50279
rect 2433 50223 2489 50279
rect 2575 50223 2631 50279
rect 2717 50223 2773 50279
rect 2859 50223 2915 50279
rect 3001 50223 3057 50279
rect 3143 50223 3199 50279
rect 3285 50223 3341 50279
rect 3427 50223 3483 50279
rect 3569 50223 3625 50279
rect 3711 50223 3767 50279
rect 3853 50223 3909 50279
rect 3995 50223 4051 50279
rect 4137 50223 4193 50279
rect 4279 50223 4335 50279
rect 4421 50223 4477 50279
rect 4563 50223 4619 50279
rect 4705 50223 4761 50279
rect 4847 50223 4903 50279
rect 4989 50223 5045 50279
rect 5131 50223 5187 50279
rect 5273 50223 5329 50279
rect 5415 50223 5471 50279
rect 5557 50223 5613 50279
rect 5699 50223 5755 50279
rect 5841 50223 5897 50279
rect 5983 50223 6039 50279
rect 6125 50223 6181 50279
rect 6267 50223 6323 50279
rect 6409 50223 6465 50279
rect 6551 50223 6607 50279
rect 6693 50223 6749 50279
rect 6835 50223 6891 50279
rect 6977 50223 7033 50279
rect 7119 50223 7175 50279
rect 7261 50223 7317 50279
rect 7403 50223 7459 50279
rect 7545 50223 7601 50279
rect 7687 50223 7743 50279
rect 7829 50223 7885 50279
rect 7971 50223 8027 50279
rect 8113 50223 8169 50279
rect 8255 50223 8311 50279
rect 8397 50223 8453 50279
rect 8539 50223 8595 50279
rect 8681 50223 8737 50279
rect 8823 50223 8879 50279
rect 8965 50223 9021 50279
rect 9107 50223 9163 50279
rect 9249 50223 9305 50279
rect 9391 50223 9447 50279
rect 9533 50223 9589 50279
rect 9675 50223 9731 50279
rect 9817 50223 9873 50279
rect 9959 50223 10015 50279
rect 10101 50223 10157 50279
rect 10243 50223 10299 50279
rect 10385 50223 10441 50279
rect 10527 50223 10583 50279
rect 10669 50223 10725 50279
rect 10811 50223 10867 50279
rect 10953 50223 11009 50279
rect 11095 50223 11151 50279
rect 11237 50223 11293 50279
rect 11379 50223 11435 50279
rect 11521 50223 11577 50279
rect 11663 50223 11719 50279
rect 11805 50223 11861 50279
rect 11947 50223 12003 50279
rect 12089 50223 12145 50279
rect 12231 50223 12287 50279
rect 12373 50223 12429 50279
rect 12515 50223 12571 50279
rect 12657 50223 12713 50279
rect 12799 50223 12855 50279
rect 12941 50223 12997 50279
rect 13083 50223 13139 50279
rect 13225 50223 13281 50279
rect 13367 50223 13423 50279
rect 13509 50223 13565 50279
rect 13651 50223 13707 50279
rect 13793 50223 13849 50279
rect 13935 50223 13991 50279
rect 14077 50223 14133 50279
rect 14219 50223 14275 50279
rect 14361 50223 14417 50279
rect 14503 50223 14559 50279
rect 14645 50223 14701 50279
rect 14787 50223 14843 50279
rect 161 50081 217 50137
rect 303 50081 359 50137
rect 445 50081 501 50137
rect 587 50081 643 50137
rect 729 50081 785 50137
rect 871 50081 927 50137
rect 1013 50081 1069 50137
rect 1155 50081 1211 50137
rect 1297 50081 1353 50137
rect 1439 50081 1495 50137
rect 1581 50081 1637 50137
rect 1723 50081 1779 50137
rect 1865 50081 1921 50137
rect 2007 50081 2063 50137
rect 2149 50081 2205 50137
rect 2291 50081 2347 50137
rect 2433 50081 2489 50137
rect 2575 50081 2631 50137
rect 2717 50081 2773 50137
rect 2859 50081 2915 50137
rect 3001 50081 3057 50137
rect 3143 50081 3199 50137
rect 3285 50081 3341 50137
rect 3427 50081 3483 50137
rect 3569 50081 3625 50137
rect 3711 50081 3767 50137
rect 3853 50081 3909 50137
rect 3995 50081 4051 50137
rect 4137 50081 4193 50137
rect 4279 50081 4335 50137
rect 4421 50081 4477 50137
rect 4563 50081 4619 50137
rect 4705 50081 4761 50137
rect 4847 50081 4903 50137
rect 4989 50081 5045 50137
rect 5131 50081 5187 50137
rect 5273 50081 5329 50137
rect 5415 50081 5471 50137
rect 5557 50081 5613 50137
rect 5699 50081 5755 50137
rect 5841 50081 5897 50137
rect 5983 50081 6039 50137
rect 6125 50081 6181 50137
rect 6267 50081 6323 50137
rect 6409 50081 6465 50137
rect 6551 50081 6607 50137
rect 6693 50081 6749 50137
rect 6835 50081 6891 50137
rect 6977 50081 7033 50137
rect 7119 50081 7175 50137
rect 7261 50081 7317 50137
rect 7403 50081 7459 50137
rect 7545 50081 7601 50137
rect 7687 50081 7743 50137
rect 7829 50081 7885 50137
rect 7971 50081 8027 50137
rect 8113 50081 8169 50137
rect 8255 50081 8311 50137
rect 8397 50081 8453 50137
rect 8539 50081 8595 50137
rect 8681 50081 8737 50137
rect 8823 50081 8879 50137
rect 8965 50081 9021 50137
rect 9107 50081 9163 50137
rect 9249 50081 9305 50137
rect 9391 50081 9447 50137
rect 9533 50081 9589 50137
rect 9675 50081 9731 50137
rect 9817 50081 9873 50137
rect 9959 50081 10015 50137
rect 10101 50081 10157 50137
rect 10243 50081 10299 50137
rect 10385 50081 10441 50137
rect 10527 50081 10583 50137
rect 10669 50081 10725 50137
rect 10811 50081 10867 50137
rect 10953 50081 11009 50137
rect 11095 50081 11151 50137
rect 11237 50081 11293 50137
rect 11379 50081 11435 50137
rect 11521 50081 11577 50137
rect 11663 50081 11719 50137
rect 11805 50081 11861 50137
rect 11947 50081 12003 50137
rect 12089 50081 12145 50137
rect 12231 50081 12287 50137
rect 12373 50081 12429 50137
rect 12515 50081 12571 50137
rect 12657 50081 12713 50137
rect 12799 50081 12855 50137
rect 12941 50081 12997 50137
rect 13083 50081 13139 50137
rect 13225 50081 13281 50137
rect 13367 50081 13423 50137
rect 13509 50081 13565 50137
rect 13651 50081 13707 50137
rect 13793 50081 13849 50137
rect 13935 50081 13991 50137
rect 14077 50081 14133 50137
rect 14219 50081 14275 50137
rect 14361 50081 14417 50137
rect 14503 50081 14559 50137
rect 14645 50081 14701 50137
rect 14787 50081 14843 50137
rect 161 49939 217 49995
rect 303 49939 359 49995
rect 445 49939 501 49995
rect 587 49939 643 49995
rect 729 49939 785 49995
rect 871 49939 927 49995
rect 1013 49939 1069 49995
rect 1155 49939 1211 49995
rect 1297 49939 1353 49995
rect 1439 49939 1495 49995
rect 1581 49939 1637 49995
rect 1723 49939 1779 49995
rect 1865 49939 1921 49995
rect 2007 49939 2063 49995
rect 2149 49939 2205 49995
rect 2291 49939 2347 49995
rect 2433 49939 2489 49995
rect 2575 49939 2631 49995
rect 2717 49939 2773 49995
rect 2859 49939 2915 49995
rect 3001 49939 3057 49995
rect 3143 49939 3199 49995
rect 3285 49939 3341 49995
rect 3427 49939 3483 49995
rect 3569 49939 3625 49995
rect 3711 49939 3767 49995
rect 3853 49939 3909 49995
rect 3995 49939 4051 49995
rect 4137 49939 4193 49995
rect 4279 49939 4335 49995
rect 4421 49939 4477 49995
rect 4563 49939 4619 49995
rect 4705 49939 4761 49995
rect 4847 49939 4903 49995
rect 4989 49939 5045 49995
rect 5131 49939 5187 49995
rect 5273 49939 5329 49995
rect 5415 49939 5471 49995
rect 5557 49939 5613 49995
rect 5699 49939 5755 49995
rect 5841 49939 5897 49995
rect 5983 49939 6039 49995
rect 6125 49939 6181 49995
rect 6267 49939 6323 49995
rect 6409 49939 6465 49995
rect 6551 49939 6607 49995
rect 6693 49939 6749 49995
rect 6835 49939 6891 49995
rect 6977 49939 7033 49995
rect 7119 49939 7175 49995
rect 7261 49939 7317 49995
rect 7403 49939 7459 49995
rect 7545 49939 7601 49995
rect 7687 49939 7743 49995
rect 7829 49939 7885 49995
rect 7971 49939 8027 49995
rect 8113 49939 8169 49995
rect 8255 49939 8311 49995
rect 8397 49939 8453 49995
rect 8539 49939 8595 49995
rect 8681 49939 8737 49995
rect 8823 49939 8879 49995
rect 8965 49939 9021 49995
rect 9107 49939 9163 49995
rect 9249 49939 9305 49995
rect 9391 49939 9447 49995
rect 9533 49939 9589 49995
rect 9675 49939 9731 49995
rect 9817 49939 9873 49995
rect 9959 49939 10015 49995
rect 10101 49939 10157 49995
rect 10243 49939 10299 49995
rect 10385 49939 10441 49995
rect 10527 49939 10583 49995
rect 10669 49939 10725 49995
rect 10811 49939 10867 49995
rect 10953 49939 11009 49995
rect 11095 49939 11151 49995
rect 11237 49939 11293 49995
rect 11379 49939 11435 49995
rect 11521 49939 11577 49995
rect 11663 49939 11719 49995
rect 11805 49939 11861 49995
rect 11947 49939 12003 49995
rect 12089 49939 12145 49995
rect 12231 49939 12287 49995
rect 12373 49939 12429 49995
rect 12515 49939 12571 49995
rect 12657 49939 12713 49995
rect 12799 49939 12855 49995
rect 12941 49939 12997 49995
rect 13083 49939 13139 49995
rect 13225 49939 13281 49995
rect 13367 49939 13423 49995
rect 13509 49939 13565 49995
rect 13651 49939 13707 49995
rect 13793 49939 13849 49995
rect 13935 49939 13991 49995
rect 14077 49939 14133 49995
rect 14219 49939 14275 49995
rect 14361 49939 14417 49995
rect 14503 49939 14559 49995
rect 14645 49939 14701 49995
rect 14787 49939 14843 49995
rect 161 49797 217 49853
rect 303 49797 359 49853
rect 445 49797 501 49853
rect 587 49797 643 49853
rect 729 49797 785 49853
rect 871 49797 927 49853
rect 1013 49797 1069 49853
rect 1155 49797 1211 49853
rect 1297 49797 1353 49853
rect 1439 49797 1495 49853
rect 1581 49797 1637 49853
rect 1723 49797 1779 49853
rect 1865 49797 1921 49853
rect 2007 49797 2063 49853
rect 2149 49797 2205 49853
rect 2291 49797 2347 49853
rect 2433 49797 2489 49853
rect 2575 49797 2631 49853
rect 2717 49797 2773 49853
rect 2859 49797 2915 49853
rect 3001 49797 3057 49853
rect 3143 49797 3199 49853
rect 3285 49797 3341 49853
rect 3427 49797 3483 49853
rect 3569 49797 3625 49853
rect 3711 49797 3767 49853
rect 3853 49797 3909 49853
rect 3995 49797 4051 49853
rect 4137 49797 4193 49853
rect 4279 49797 4335 49853
rect 4421 49797 4477 49853
rect 4563 49797 4619 49853
rect 4705 49797 4761 49853
rect 4847 49797 4903 49853
rect 4989 49797 5045 49853
rect 5131 49797 5187 49853
rect 5273 49797 5329 49853
rect 5415 49797 5471 49853
rect 5557 49797 5613 49853
rect 5699 49797 5755 49853
rect 5841 49797 5897 49853
rect 5983 49797 6039 49853
rect 6125 49797 6181 49853
rect 6267 49797 6323 49853
rect 6409 49797 6465 49853
rect 6551 49797 6607 49853
rect 6693 49797 6749 49853
rect 6835 49797 6891 49853
rect 6977 49797 7033 49853
rect 7119 49797 7175 49853
rect 7261 49797 7317 49853
rect 7403 49797 7459 49853
rect 7545 49797 7601 49853
rect 7687 49797 7743 49853
rect 7829 49797 7885 49853
rect 7971 49797 8027 49853
rect 8113 49797 8169 49853
rect 8255 49797 8311 49853
rect 8397 49797 8453 49853
rect 8539 49797 8595 49853
rect 8681 49797 8737 49853
rect 8823 49797 8879 49853
rect 8965 49797 9021 49853
rect 9107 49797 9163 49853
rect 9249 49797 9305 49853
rect 9391 49797 9447 49853
rect 9533 49797 9589 49853
rect 9675 49797 9731 49853
rect 9817 49797 9873 49853
rect 9959 49797 10015 49853
rect 10101 49797 10157 49853
rect 10243 49797 10299 49853
rect 10385 49797 10441 49853
rect 10527 49797 10583 49853
rect 10669 49797 10725 49853
rect 10811 49797 10867 49853
rect 10953 49797 11009 49853
rect 11095 49797 11151 49853
rect 11237 49797 11293 49853
rect 11379 49797 11435 49853
rect 11521 49797 11577 49853
rect 11663 49797 11719 49853
rect 11805 49797 11861 49853
rect 11947 49797 12003 49853
rect 12089 49797 12145 49853
rect 12231 49797 12287 49853
rect 12373 49797 12429 49853
rect 12515 49797 12571 49853
rect 12657 49797 12713 49853
rect 12799 49797 12855 49853
rect 12941 49797 12997 49853
rect 13083 49797 13139 49853
rect 13225 49797 13281 49853
rect 13367 49797 13423 49853
rect 13509 49797 13565 49853
rect 13651 49797 13707 49853
rect 13793 49797 13849 49853
rect 13935 49797 13991 49853
rect 14077 49797 14133 49853
rect 14219 49797 14275 49853
rect 14361 49797 14417 49853
rect 14503 49797 14559 49853
rect 14645 49797 14701 49853
rect 14787 49797 14843 49853
rect 161 49655 217 49711
rect 303 49655 359 49711
rect 445 49655 501 49711
rect 587 49655 643 49711
rect 729 49655 785 49711
rect 871 49655 927 49711
rect 1013 49655 1069 49711
rect 1155 49655 1211 49711
rect 1297 49655 1353 49711
rect 1439 49655 1495 49711
rect 1581 49655 1637 49711
rect 1723 49655 1779 49711
rect 1865 49655 1921 49711
rect 2007 49655 2063 49711
rect 2149 49655 2205 49711
rect 2291 49655 2347 49711
rect 2433 49655 2489 49711
rect 2575 49655 2631 49711
rect 2717 49655 2773 49711
rect 2859 49655 2915 49711
rect 3001 49655 3057 49711
rect 3143 49655 3199 49711
rect 3285 49655 3341 49711
rect 3427 49655 3483 49711
rect 3569 49655 3625 49711
rect 3711 49655 3767 49711
rect 3853 49655 3909 49711
rect 3995 49655 4051 49711
rect 4137 49655 4193 49711
rect 4279 49655 4335 49711
rect 4421 49655 4477 49711
rect 4563 49655 4619 49711
rect 4705 49655 4761 49711
rect 4847 49655 4903 49711
rect 4989 49655 5045 49711
rect 5131 49655 5187 49711
rect 5273 49655 5329 49711
rect 5415 49655 5471 49711
rect 5557 49655 5613 49711
rect 5699 49655 5755 49711
rect 5841 49655 5897 49711
rect 5983 49655 6039 49711
rect 6125 49655 6181 49711
rect 6267 49655 6323 49711
rect 6409 49655 6465 49711
rect 6551 49655 6607 49711
rect 6693 49655 6749 49711
rect 6835 49655 6891 49711
rect 6977 49655 7033 49711
rect 7119 49655 7175 49711
rect 7261 49655 7317 49711
rect 7403 49655 7459 49711
rect 7545 49655 7601 49711
rect 7687 49655 7743 49711
rect 7829 49655 7885 49711
rect 7971 49655 8027 49711
rect 8113 49655 8169 49711
rect 8255 49655 8311 49711
rect 8397 49655 8453 49711
rect 8539 49655 8595 49711
rect 8681 49655 8737 49711
rect 8823 49655 8879 49711
rect 8965 49655 9021 49711
rect 9107 49655 9163 49711
rect 9249 49655 9305 49711
rect 9391 49655 9447 49711
rect 9533 49655 9589 49711
rect 9675 49655 9731 49711
rect 9817 49655 9873 49711
rect 9959 49655 10015 49711
rect 10101 49655 10157 49711
rect 10243 49655 10299 49711
rect 10385 49655 10441 49711
rect 10527 49655 10583 49711
rect 10669 49655 10725 49711
rect 10811 49655 10867 49711
rect 10953 49655 11009 49711
rect 11095 49655 11151 49711
rect 11237 49655 11293 49711
rect 11379 49655 11435 49711
rect 11521 49655 11577 49711
rect 11663 49655 11719 49711
rect 11805 49655 11861 49711
rect 11947 49655 12003 49711
rect 12089 49655 12145 49711
rect 12231 49655 12287 49711
rect 12373 49655 12429 49711
rect 12515 49655 12571 49711
rect 12657 49655 12713 49711
rect 12799 49655 12855 49711
rect 12941 49655 12997 49711
rect 13083 49655 13139 49711
rect 13225 49655 13281 49711
rect 13367 49655 13423 49711
rect 13509 49655 13565 49711
rect 13651 49655 13707 49711
rect 13793 49655 13849 49711
rect 13935 49655 13991 49711
rect 14077 49655 14133 49711
rect 14219 49655 14275 49711
rect 14361 49655 14417 49711
rect 14503 49655 14559 49711
rect 14645 49655 14701 49711
rect 14787 49655 14843 49711
rect 161 49513 217 49569
rect 303 49513 359 49569
rect 445 49513 501 49569
rect 587 49513 643 49569
rect 729 49513 785 49569
rect 871 49513 927 49569
rect 1013 49513 1069 49569
rect 1155 49513 1211 49569
rect 1297 49513 1353 49569
rect 1439 49513 1495 49569
rect 1581 49513 1637 49569
rect 1723 49513 1779 49569
rect 1865 49513 1921 49569
rect 2007 49513 2063 49569
rect 2149 49513 2205 49569
rect 2291 49513 2347 49569
rect 2433 49513 2489 49569
rect 2575 49513 2631 49569
rect 2717 49513 2773 49569
rect 2859 49513 2915 49569
rect 3001 49513 3057 49569
rect 3143 49513 3199 49569
rect 3285 49513 3341 49569
rect 3427 49513 3483 49569
rect 3569 49513 3625 49569
rect 3711 49513 3767 49569
rect 3853 49513 3909 49569
rect 3995 49513 4051 49569
rect 4137 49513 4193 49569
rect 4279 49513 4335 49569
rect 4421 49513 4477 49569
rect 4563 49513 4619 49569
rect 4705 49513 4761 49569
rect 4847 49513 4903 49569
rect 4989 49513 5045 49569
rect 5131 49513 5187 49569
rect 5273 49513 5329 49569
rect 5415 49513 5471 49569
rect 5557 49513 5613 49569
rect 5699 49513 5755 49569
rect 5841 49513 5897 49569
rect 5983 49513 6039 49569
rect 6125 49513 6181 49569
rect 6267 49513 6323 49569
rect 6409 49513 6465 49569
rect 6551 49513 6607 49569
rect 6693 49513 6749 49569
rect 6835 49513 6891 49569
rect 6977 49513 7033 49569
rect 7119 49513 7175 49569
rect 7261 49513 7317 49569
rect 7403 49513 7459 49569
rect 7545 49513 7601 49569
rect 7687 49513 7743 49569
rect 7829 49513 7885 49569
rect 7971 49513 8027 49569
rect 8113 49513 8169 49569
rect 8255 49513 8311 49569
rect 8397 49513 8453 49569
rect 8539 49513 8595 49569
rect 8681 49513 8737 49569
rect 8823 49513 8879 49569
rect 8965 49513 9021 49569
rect 9107 49513 9163 49569
rect 9249 49513 9305 49569
rect 9391 49513 9447 49569
rect 9533 49513 9589 49569
rect 9675 49513 9731 49569
rect 9817 49513 9873 49569
rect 9959 49513 10015 49569
rect 10101 49513 10157 49569
rect 10243 49513 10299 49569
rect 10385 49513 10441 49569
rect 10527 49513 10583 49569
rect 10669 49513 10725 49569
rect 10811 49513 10867 49569
rect 10953 49513 11009 49569
rect 11095 49513 11151 49569
rect 11237 49513 11293 49569
rect 11379 49513 11435 49569
rect 11521 49513 11577 49569
rect 11663 49513 11719 49569
rect 11805 49513 11861 49569
rect 11947 49513 12003 49569
rect 12089 49513 12145 49569
rect 12231 49513 12287 49569
rect 12373 49513 12429 49569
rect 12515 49513 12571 49569
rect 12657 49513 12713 49569
rect 12799 49513 12855 49569
rect 12941 49513 12997 49569
rect 13083 49513 13139 49569
rect 13225 49513 13281 49569
rect 13367 49513 13423 49569
rect 13509 49513 13565 49569
rect 13651 49513 13707 49569
rect 13793 49513 13849 49569
rect 13935 49513 13991 49569
rect 14077 49513 14133 49569
rect 14219 49513 14275 49569
rect 14361 49513 14417 49569
rect 14503 49513 14559 49569
rect 14645 49513 14701 49569
rect 14787 49513 14843 49569
rect 161 49371 217 49427
rect 303 49371 359 49427
rect 445 49371 501 49427
rect 587 49371 643 49427
rect 729 49371 785 49427
rect 871 49371 927 49427
rect 1013 49371 1069 49427
rect 1155 49371 1211 49427
rect 1297 49371 1353 49427
rect 1439 49371 1495 49427
rect 1581 49371 1637 49427
rect 1723 49371 1779 49427
rect 1865 49371 1921 49427
rect 2007 49371 2063 49427
rect 2149 49371 2205 49427
rect 2291 49371 2347 49427
rect 2433 49371 2489 49427
rect 2575 49371 2631 49427
rect 2717 49371 2773 49427
rect 2859 49371 2915 49427
rect 3001 49371 3057 49427
rect 3143 49371 3199 49427
rect 3285 49371 3341 49427
rect 3427 49371 3483 49427
rect 3569 49371 3625 49427
rect 3711 49371 3767 49427
rect 3853 49371 3909 49427
rect 3995 49371 4051 49427
rect 4137 49371 4193 49427
rect 4279 49371 4335 49427
rect 4421 49371 4477 49427
rect 4563 49371 4619 49427
rect 4705 49371 4761 49427
rect 4847 49371 4903 49427
rect 4989 49371 5045 49427
rect 5131 49371 5187 49427
rect 5273 49371 5329 49427
rect 5415 49371 5471 49427
rect 5557 49371 5613 49427
rect 5699 49371 5755 49427
rect 5841 49371 5897 49427
rect 5983 49371 6039 49427
rect 6125 49371 6181 49427
rect 6267 49371 6323 49427
rect 6409 49371 6465 49427
rect 6551 49371 6607 49427
rect 6693 49371 6749 49427
rect 6835 49371 6891 49427
rect 6977 49371 7033 49427
rect 7119 49371 7175 49427
rect 7261 49371 7317 49427
rect 7403 49371 7459 49427
rect 7545 49371 7601 49427
rect 7687 49371 7743 49427
rect 7829 49371 7885 49427
rect 7971 49371 8027 49427
rect 8113 49371 8169 49427
rect 8255 49371 8311 49427
rect 8397 49371 8453 49427
rect 8539 49371 8595 49427
rect 8681 49371 8737 49427
rect 8823 49371 8879 49427
rect 8965 49371 9021 49427
rect 9107 49371 9163 49427
rect 9249 49371 9305 49427
rect 9391 49371 9447 49427
rect 9533 49371 9589 49427
rect 9675 49371 9731 49427
rect 9817 49371 9873 49427
rect 9959 49371 10015 49427
rect 10101 49371 10157 49427
rect 10243 49371 10299 49427
rect 10385 49371 10441 49427
rect 10527 49371 10583 49427
rect 10669 49371 10725 49427
rect 10811 49371 10867 49427
rect 10953 49371 11009 49427
rect 11095 49371 11151 49427
rect 11237 49371 11293 49427
rect 11379 49371 11435 49427
rect 11521 49371 11577 49427
rect 11663 49371 11719 49427
rect 11805 49371 11861 49427
rect 11947 49371 12003 49427
rect 12089 49371 12145 49427
rect 12231 49371 12287 49427
rect 12373 49371 12429 49427
rect 12515 49371 12571 49427
rect 12657 49371 12713 49427
rect 12799 49371 12855 49427
rect 12941 49371 12997 49427
rect 13083 49371 13139 49427
rect 13225 49371 13281 49427
rect 13367 49371 13423 49427
rect 13509 49371 13565 49427
rect 13651 49371 13707 49427
rect 13793 49371 13849 49427
rect 13935 49371 13991 49427
rect 14077 49371 14133 49427
rect 14219 49371 14275 49427
rect 14361 49371 14417 49427
rect 14503 49371 14559 49427
rect 14645 49371 14701 49427
rect 14787 49371 14843 49427
rect 161 49229 217 49285
rect 303 49229 359 49285
rect 445 49229 501 49285
rect 587 49229 643 49285
rect 729 49229 785 49285
rect 871 49229 927 49285
rect 1013 49229 1069 49285
rect 1155 49229 1211 49285
rect 1297 49229 1353 49285
rect 1439 49229 1495 49285
rect 1581 49229 1637 49285
rect 1723 49229 1779 49285
rect 1865 49229 1921 49285
rect 2007 49229 2063 49285
rect 2149 49229 2205 49285
rect 2291 49229 2347 49285
rect 2433 49229 2489 49285
rect 2575 49229 2631 49285
rect 2717 49229 2773 49285
rect 2859 49229 2915 49285
rect 3001 49229 3057 49285
rect 3143 49229 3199 49285
rect 3285 49229 3341 49285
rect 3427 49229 3483 49285
rect 3569 49229 3625 49285
rect 3711 49229 3767 49285
rect 3853 49229 3909 49285
rect 3995 49229 4051 49285
rect 4137 49229 4193 49285
rect 4279 49229 4335 49285
rect 4421 49229 4477 49285
rect 4563 49229 4619 49285
rect 4705 49229 4761 49285
rect 4847 49229 4903 49285
rect 4989 49229 5045 49285
rect 5131 49229 5187 49285
rect 5273 49229 5329 49285
rect 5415 49229 5471 49285
rect 5557 49229 5613 49285
rect 5699 49229 5755 49285
rect 5841 49229 5897 49285
rect 5983 49229 6039 49285
rect 6125 49229 6181 49285
rect 6267 49229 6323 49285
rect 6409 49229 6465 49285
rect 6551 49229 6607 49285
rect 6693 49229 6749 49285
rect 6835 49229 6891 49285
rect 6977 49229 7033 49285
rect 7119 49229 7175 49285
rect 7261 49229 7317 49285
rect 7403 49229 7459 49285
rect 7545 49229 7601 49285
rect 7687 49229 7743 49285
rect 7829 49229 7885 49285
rect 7971 49229 8027 49285
rect 8113 49229 8169 49285
rect 8255 49229 8311 49285
rect 8397 49229 8453 49285
rect 8539 49229 8595 49285
rect 8681 49229 8737 49285
rect 8823 49229 8879 49285
rect 8965 49229 9021 49285
rect 9107 49229 9163 49285
rect 9249 49229 9305 49285
rect 9391 49229 9447 49285
rect 9533 49229 9589 49285
rect 9675 49229 9731 49285
rect 9817 49229 9873 49285
rect 9959 49229 10015 49285
rect 10101 49229 10157 49285
rect 10243 49229 10299 49285
rect 10385 49229 10441 49285
rect 10527 49229 10583 49285
rect 10669 49229 10725 49285
rect 10811 49229 10867 49285
rect 10953 49229 11009 49285
rect 11095 49229 11151 49285
rect 11237 49229 11293 49285
rect 11379 49229 11435 49285
rect 11521 49229 11577 49285
rect 11663 49229 11719 49285
rect 11805 49229 11861 49285
rect 11947 49229 12003 49285
rect 12089 49229 12145 49285
rect 12231 49229 12287 49285
rect 12373 49229 12429 49285
rect 12515 49229 12571 49285
rect 12657 49229 12713 49285
rect 12799 49229 12855 49285
rect 12941 49229 12997 49285
rect 13083 49229 13139 49285
rect 13225 49229 13281 49285
rect 13367 49229 13423 49285
rect 13509 49229 13565 49285
rect 13651 49229 13707 49285
rect 13793 49229 13849 49285
rect 13935 49229 13991 49285
rect 14077 49229 14133 49285
rect 14219 49229 14275 49285
rect 14361 49229 14417 49285
rect 14503 49229 14559 49285
rect 14645 49229 14701 49285
rect 14787 49229 14843 49285
rect 161 48885 217 48941
rect 303 48885 359 48941
rect 445 48885 501 48941
rect 587 48885 643 48941
rect 729 48885 785 48941
rect 871 48885 927 48941
rect 1013 48885 1069 48941
rect 1155 48885 1211 48941
rect 1297 48885 1353 48941
rect 1439 48885 1495 48941
rect 1581 48885 1637 48941
rect 1723 48885 1779 48941
rect 1865 48885 1921 48941
rect 2007 48885 2063 48941
rect 2149 48885 2205 48941
rect 2291 48885 2347 48941
rect 2433 48885 2489 48941
rect 2575 48885 2631 48941
rect 2717 48885 2773 48941
rect 2859 48885 2915 48941
rect 3001 48885 3057 48941
rect 3143 48885 3199 48941
rect 3285 48885 3341 48941
rect 3427 48885 3483 48941
rect 3569 48885 3625 48941
rect 3711 48885 3767 48941
rect 3853 48885 3909 48941
rect 3995 48885 4051 48941
rect 4137 48885 4193 48941
rect 4279 48885 4335 48941
rect 4421 48885 4477 48941
rect 4563 48885 4619 48941
rect 4705 48885 4761 48941
rect 4847 48885 4903 48941
rect 4989 48885 5045 48941
rect 5131 48885 5187 48941
rect 5273 48885 5329 48941
rect 5415 48885 5471 48941
rect 5557 48885 5613 48941
rect 5699 48885 5755 48941
rect 5841 48885 5897 48941
rect 5983 48885 6039 48941
rect 6125 48885 6181 48941
rect 6267 48885 6323 48941
rect 6409 48885 6465 48941
rect 6551 48885 6607 48941
rect 6693 48885 6749 48941
rect 6835 48885 6891 48941
rect 6977 48885 7033 48941
rect 7119 48885 7175 48941
rect 7261 48885 7317 48941
rect 7403 48885 7459 48941
rect 7545 48885 7601 48941
rect 7687 48885 7743 48941
rect 7829 48885 7885 48941
rect 7971 48885 8027 48941
rect 8113 48885 8169 48941
rect 8255 48885 8311 48941
rect 8397 48885 8453 48941
rect 8539 48885 8595 48941
rect 8681 48885 8737 48941
rect 8823 48885 8879 48941
rect 8965 48885 9021 48941
rect 9107 48885 9163 48941
rect 9249 48885 9305 48941
rect 9391 48885 9447 48941
rect 9533 48885 9589 48941
rect 9675 48885 9731 48941
rect 9817 48885 9873 48941
rect 9959 48885 10015 48941
rect 10101 48885 10157 48941
rect 10243 48885 10299 48941
rect 10385 48885 10441 48941
rect 10527 48885 10583 48941
rect 10669 48885 10725 48941
rect 10811 48885 10867 48941
rect 10953 48885 11009 48941
rect 11095 48885 11151 48941
rect 11237 48885 11293 48941
rect 11379 48885 11435 48941
rect 11521 48885 11577 48941
rect 11663 48885 11719 48941
rect 11805 48885 11861 48941
rect 11947 48885 12003 48941
rect 12089 48885 12145 48941
rect 12231 48885 12287 48941
rect 12373 48885 12429 48941
rect 12515 48885 12571 48941
rect 12657 48885 12713 48941
rect 12799 48885 12855 48941
rect 12941 48885 12997 48941
rect 13083 48885 13139 48941
rect 13225 48885 13281 48941
rect 13367 48885 13423 48941
rect 13509 48885 13565 48941
rect 13651 48885 13707 48941
rect 13793 48885 13849 48941
rect 13935 48885 13991 48941
rect 14077 48885 14133 48941
rect 14219 48885 14275 48941
rect 14361 48885 14417 48941
rect 14503 48885 14559 48941
rect 14645 48885 14701 48941
rect 14787 48885 14843 48941
rect 161 48743 217 48799
rect 303 48743 359 48799
rect 445 48743 501 48799
rect 587 48743 643 48799
rect 729 48743 785 48799
rect 871 48743 927 48799
rect 1013 48743 1069 48799
rect 1155 48743 1211 48799
rect 1297 48743 1353 48799
rect 1439 48743 1495 48799
rect 1581 48743 1637 48799
rect 1723 48743 1779 48799
rect 1865 48743 1921 48799
rect 2007 48743 2063 48799
rect 2149 48743 2205 48799
rect 2291 48743 2347 48799
rect 2433 48743 2489 48799
rect 2575 48743 2631 48799
rect 2717 48743 2773 48799
rect 2859 48743 2915 48799
rect 3001 48743 3057 48799
rect 3143 48743 3199 48799
rect 3285 48743 3341 48799
rect 3427 48743 3483 48799
rect 3569 48743 3625 48799
rect 3711 48743 3767 48799
rect 3853 48743 3909 48799
rect 3995 48743 4051 48799
rect 4137 48743 4193 48799
rect 4279 48743 4335 48799
rect 4421 48743 4477 48799
rect 4563 48743 4619 48799
rect 4705 48743 4761 48799
rect 4847 48743 4903 48799
rect 4989 48743 5045 48799
rect 5131 48743 5187 48799
rect 5273 48743 5329 48799
rect 5415 48743 5471 48799
rect 5557 48743 5613 48799
rect 5699 48743 5755 48799
rect 5841 48743 5897 48799
rect 5983 48743 6039 48799
rect 6125 48743 6181 48799
rect 6267 48743 6323 48799
rect 6409 48743 6465 48799
rect 6551 48743 6607 48799
rect 6693 48743 6749 48799
rect 6835 48743 6891 48799
rect 6977 48743 7033 48799
rect 7119 48743 7175 48799
rect 7261 48743 7317 48799
rect 7403 48743 7459 48799
rect 7545 48743 7601 48799
rect 7687 48743 7743 48799
rect 7829 48743 7885 48799
rect 7971 48743 8027 48799
rect 8113 48743 8169 48799
rect 8255 48743 8311 48799
rect 8397 48743 8453 48799
rect 8539 48743 8595 48799
rect 8681 48743 8737 48799
rect 8823 48743 8879 48799
rect 8965 48743 9021 48799
rect 9107 48743 9163 48799
rect 9249 48743 9305 48799
rect 9391 48743 9447 48799
rect 9533 48743 9589 48799
rect 9675 48743 9731 48799
rect 9817 48743 9873 48799
rect 9959 48743 10015 48799
rect 10101 48743 10157 48799
rect 10243 48743 10299 48799
rect 10385 48743 10441 48799
rect 10527 48743 10583 48799
rect 10669 48743 10725 48799
rect 10811 48743 10867 48799
rect 10953 48743 11009 48799
rect 11095 48743 11151 48799
rect 11237 48743 11293 48799
rect 11379 48743 11435 48799
rect 11521 48743 11577 48799
rect 11663 48743 11719 48799
rect 11805 48743 11861 48799
rect 11947 48743 12003 48799
rect 12089 48743 12145 48799
rect 12231 48743 12287 48799
rect 12373 48743 12429 48799
rect 12515 48743 12571 48799
rect 12657 48743 12713 48799
rect 12799 48743 12855 48799
rect 12941 48743 12997 48799
rect 13083 48743 13139 48799
rect 13225 48743 13281 48799
rect 13367 48743 13423 48799
rect 13509 48743 13565 48799
rect 13651 48743 13707 48799
rect 13793 48743 13849 48799
rect 13935 48743 13991 48799
rect 14077 48743 14133 48799
rect 14219 48743 14275 48799
rect 14361 48743 14417 48799
rect 14503 48743 14559 48799
rect 14645 48743 14701 48799
rect 14787 48743 14843 48799
rect 161 48601 217 48657
rect 303 48601 359 48657
rect 445 48601 501 48657
rect 587 48601 643 48657
rect 729 48601 785 48657
rect 871 48601 927 48657
rect 1013 48601 1069 48657
rect 1155 48601 1211 48657
rect 1297 48601 1353 48657
rect 1439 48601 1495 48657
rect 1581 48601 1637 48657
rect 1723 48601 1779 48657
rect 1865 48601 1921 48657
rect 2007 48601 2063 48657
rect 2149 48601 2205 48657
rect 2291 48601 2347 48657
rect 2433 48601 2489 48657
rect 2575 48601 2631 48657
rect 2717 48601 2773 48657
rect 2859 48601 2915 48657
rect 3001 48601 3057 48657
rect 3143 48601 3199 48657
rect 3285 48601 3341 48657
rect 3427 48601 3483 48657
rect 3569 48601 3625 48657
rect 3711 48601 3767 48657
rect 3853 48601 3909 48657
rect 3995 48601 4051 48657
rect 4137 48601 4193 48657
rect 4279 48601 4335 48657
rect 4421 48601 4477 48657
rect 4563 48601 4619 48657
rect 4705 48601 4761 48657
rect 4847 48601 4903 48657
rect 4989 48601 5045 48657
rect 5131 48601 5187 48657
rect 5273 48601 5329 48657
rect 5415 48601 5471 48657
rect 5557 48601 5613 48657
rect 5699 48601 5755 48657
rect 5841 48601 5897 48657
rect 5983 48601 6039 48657
rect 6125 48601 6181 48657
rect 6267 48601 6323 48657
rect 6409 48601 6465 48657
rect 6551 48601 6607 48657
rect 6693 48601 6749 48657
rect 6835 48601 6891 48657
rect 6977 48601 7033 48657
rect 7119 48601 7175 48657
rect 7261 48601 7317 48657
rect 7403 48601 7459 48657
rect 7545 48601 7601 48657
rect 7687 48601 7743 48657
rect 7829 48601 7885 48657
rect 7971 48601 8027 48657
rect 8113 48601 8169 48657
rect 8255 48601 8311 48657
rect 8397 48601 8453 48657
rect 8539 48601 8595 48657
rect 8681 48601 8737 48657
rect 8823 48601 8879 48657
rect 8965 48601 9021 48657
rect 9107 48601 9163 48657
rect 9249 48601 9305 48657
rect 9391 48601 9447 48657
rect 9533 48601 9589 48657
rect 9675 48601 9731 48657
rect 9817 48601 9873 48657
rect 9959 48601 10015 48657
rect 10101 48601 10157 48657
rect 10243 48601 10299 48657
rect 10385 48601 10441 48657
rect 10527 48601 10583 48657
rect 10669 48601 10725 48657
rect 10811 48601 10867 48657
rect 10953 48601 11009 48657
rect 11095 48601 11151 48657
rect 11237 48601 11293 48657
rect 11379 48601 11435 48657
rect 11521 48601 11577 48657
rect 11663 48601 11719 48657
rect 11805 48601 11861 48657
rect 11947 48601 12003 48657
rect 12089 48601 12145 48657
rect 12231 48601 12287 48657
rect 12373 48601 12429 48657
rect 12515 48601 12571 48657
rect 12657 48601 12713 48657
rect 12799 48601 12855 48657
rect 12941 48601 12997 48657
rect 13083 48601 13139 48657
rect 13225 48601 13281 48657
rect 13367 48601 13423 48657
rect 13509 48601 13565 48657
rect 13651 48601 13707 48657
rect 13793 48601 13849 48657
rect 13935 48601 13991 48657
rect 14077 48601 14133 48657
rect 14219 48601 14275 48657
rect 14361 48601 14417 48657
rect 14503 48601 14559 48657
rect 14645 48601 14701 48657
rect 14787 48601 14843 48657
rect 161 48459 217 48515
rect 303 48459 359 48515
rect 445 48459 501 48515
rect 587 48459 643 48515
rect 729 48459 785 48515
rect 871 48459 927 48515
rect 1013 48459 1069 48515
rect 1155 48459 1211 48515
rect 1297 48459 1353 48515
rect 1439 48459 1495 48515
rect 1581 48459 1637 48515
rect 1723 48459 1779 48515
rect 1865 48459 1921 48515
rect 2007 48459 2063 48515
rect 2149 48459 2205 48515
rect 2291 48459 2347 48515
rect 2433 48459 2489 48515
rect 2575 48459 2631 48515
rect 2717 48459 2773 48515
rect 2859 48459 2915 48515
rect 3001 48459 3057 48515
rect 3143 48459 3199 48515
rect 3285 48459 3341 48515
rect 3427 48459 3483 48515
rect 3569 48459 3625 48515
rect 3711 48459 3767 48515
rect 3853 48459 3909 48515
rect 3995 48459 4051 48515
rect 4137 48459 4193 48515
rect 4279 48459 4335 48515
rect 4421 48459 4477 48515
rect 4563 48459 4619 48515
rect 4705 48459 4761 48515
rect 4847 48459 4903 48515
rect 4989 48459 5045 48515
rect 5131 48459 5187 48515
rect 5273 48459 5329 48515
rect 5415 48459 5471 48515
rect 5557 48459 5613 48515
rect 5699 48459 5755 48515
rect 5841 48459 5897 48515
rect 5983 48459 6039 48515
rect 6125 48459 6181 48515
rect 6267 48459 6323 48515
rect 6409 48459 6465 48515
rect 6551 48459 6607 48515
rect 6693 48459 6749 48515
rect 6835 48459 6891 48515
rect 6977 48459 7033 48515
rect 7119 48459 7175 48515
rect 7261 48459 7317 48515
rect 7403 48459 7459 48515
rect 7545 48459 7601 48515
rect 7687 48459 7743 48515
rect 7829 48459 7885 48515
rect 7971 48459 8027 48515
rect 8113 48459 8169 48515
rect 8255 48459 8311 48515
rect 8397 48459 8453 48515
rect 8539 48459 8595 48515
rect 8681 48459 8737 48515
rect 8823 48459 8879 48515
rect 8965 48459 9021 48515
rect 9107 48459 9163 48515
rect 9249 48459 9305 48515
rect 9391 48459 9447 48515
rect 9533 48459 9589 48515
rect 9675 48459 9731 48515
rect 9817 48459 9873 48515
rect 9959 48459 10015 48515
rect 10101 48459 10157 48515
rect 10243 48459 10299 48515
rect 10385 48459 10441 48515
rect 10527 48459 10583 48515
rect 10669 48459 10725 48515
rect 10811 48459 10867 48515
rect 10953 48459 11009 48515
rect 11095 48459 11151 48515
rect 11237 48459 11293 48515
rect 11379 48459 11435 48515
rect 11521 48459 11577 48515
rect 11663 48459 11719 48515
rect 11805 48459 11861 48515
rect 11947 48459 12003 48515
rect 12089 48459 12145 48515
rect 12231 48459 12287 48515
rect 12373 48459 12429 48515
rect 12515 48459 12571 48515
rect 12657 48459 12713 48515
rect 12799 48459 12855 48515
rect 12941 48459 12997 48515
rect 13083 48459 13139 48515
rect 13225 48459 13281 48515
rect 13367 48459 13423 48515
rect 13509 48459 13565 48515
rect 13651 48459 13707 48515
rect 13793 48459 13849 48515
rect 13935 48459 13991 48515
rect 14077 48459 14133 48515
rect 14219 48459 14275 48515
rect 14361 48459 14417 48515
rect 14503 48459 14559 48515
rect 14645 48459 14701 48515
rect 14787 48459 14843 48515
rect 161 48317 217 48373
rect 303 48317 359 48373
rect 445 48317 501 48373
rect 587 48317 643 48373
rect 729 48317 785 48373
rect 871 48317 927 48373
rect 1013 48317 1069 48373
rect 1155 48317 1211 48373
rect 1297 48317 1353 48373
rect 1439 48317 1495 48373
rect 1581 48317 1637 48373
rect 1723 48317 1779 48373
rect 1865 48317 1921 48373
rect 2007 48317 2063 48373
rect 2149 48317 2205 48373
rect 2291 48317 2347 48373
rect 2433 48317 2489 48373
rect 2575 48317 2631 48373
rect 2717 48317 2773 48373
rect 2859 48317 2915 48373
rect 3001 48317 3057 48373
rect 3143 48317 3199 48373
rect 3285 48317 3341 48373
rect 3427 48317 3483 48373
rect 3569 48317 3625 48373
rect 3711 48317 3767 48373
rect 3853 48317 3909 48373
rect 3995 48317 4051 48373
rect 4137 48317 4193 48373
rect 4279 48317 4335 48373
rect 4421 48317 4477 48373
rect 4563 48317 4619 48373
rect 4705 48317 4761 48373
rect 4847 48317 4903 48373
rect 4989 48317 5045 48373
rect 5131 48317 5187 48373
rect 5273 48317 5329 48373
rect 5415 48317 5471 48373
rect 5557 48317 5613 48373
rect 5699 48317 5755 48373
rect 5841 48317 5897 48373
rect 5983 48317 6039 48373
rect 6125 48317 6181 48373
rect 6267 48317 6323 48373
rect 6409 48317 6465 48373
rect 6551 48317 6607 48373
rect 6693 48317 6749 48373
rect 6835 48317 6891 48373
rect 6977 48317 7033 48373
rect 7119 48317 7175 48373
rect 7261 48317 7317 48373
rect 7403 48317 7459 48373
rect 7545 48317 7601 48373
rect 7687 48317 7743 48373
rect 7829 48317 7885 48373
rect 7971 48317 8027 48373
rect 8113 48317 8169 48373
rect 8255 48317 8311 48373
rect 8397 48317 8453 48373
rect 8539 48317 8595 48373
rect 8681 48317 8737 48373
rect 8823 48317 8879 48373
rect 8965 48317 9021 48373
rect 9107 48317 9163 48373
rect 9249 48317 9305 48373
rect 9391 48317 9447 48373
rect 9533 48317 9589 48373
rect 9675 48317 9731 48373
rect 9817 48317 9873 48373
rect 9959 48317 10015 48373
rect 10101 48317 10157 48373
rect 10243 48317 10299 48373
rect 10385 48317 10441 48373
rect 10527 48317 10583 48373
rect 10669 48317 10725 48373
rect 10811 48317 10867 48373
rect 10953 48317 11009 48373
rect 11095 48317 11151 48373
rect 11237 48317 11293 48373
rect 11379 48317 11435 48373
rect 11521 48317 11577 48373
rect 11663 48317 11719 48373
rect 11805 48317 11861 48373
rect 11947 48317 12003 48373
rect 12089 48317 12145 48373
rect 12231 48317 12287 48373
rect 12373 48317 12429 48373
rect 12515 48317 12571 48373
rect 12657 48317 12713 48373
rect 12799 48317 12855 48373
rect 12941 48317 12997 48373
rect 13083 48317 13139 48373
rect 13225 48317 13281 48373
rect 13367 48317 13423 48373
rect 13509 48317 13565 48373
rect 13651 48317 13707 48373
rect 13793 48317 13849 48373
rect 13935 48317 13991 48373
rect 14077 48317 14133 48373
rect 14219 48317 14275 48373
rect 14361 48317 14417 48373
rect 14503 48317 14559 48373
rect 14645 48317 14701 48373
rect 14787 48317 14843 48373
rect 161 48175 217 48231
rect 303 48175 359 48231
rect 445 48175 501 48231
rect 587 48175 643 48231
rect 729 48175 785 48231
rect 871 48175 927 48231
rect 1013 48175 1069 48231
rect 1155 48175 1211 48231
rect 1297 48175 1353 48231
rect 1439 48175 1495 48231
rect 1581 48175 1637 48231
rect 1723 48175 1779 48231
rect 1865 48175 1921 48231
rect 2007 48175 2063 48231
rect 2149 48175 2205 48231
rect 2291 48175 2347 48231
rect 2433 48175 2489 48231
rect 2575 48175 2631 48231
rect 2717 48175 2773 48231
rect 2859 48175 2915 48231
rect 3001 48175 3057 48231
rect 3143 48175 3199 48231
rect 3285 48175 3341 48231
rect 3427 48175 3483 48231
rect 3569 48175 3625 48231
rect 3711 48175 3767 48231
rect 3853 48175 3909 48231
rect 3995 48175 4051 48231
rect 4137 48175 4193 48231
rect 4279 48175 4335 48231
rect 4421 48175 4477 48231
rect 4563 48175 4619 48231
rect 4705 48175 4761 48231
rect 4847 48175 4903 48231
rect 4989 48175 5045 48231
rect 5131 48175 5187 48231
rect 5273 48175 5329 48231
rect 5415 48175 5471 48231
rect 5557 48175 5613 48231
rect 5699 48175 5755 48231
rect 5841 48175 5897 48231
rect 5983 48175 6039 48231
rect 6125 48175 6181 48231
rect 6267 48175 6323 48231
rect 6409 48175 6465 48231
rect 6551 48175 6607 48231
rect 6693 48175 6749 48231
rect 6835 48175 6891 48231
rect 6977 48175 7033 48231
rect 7119 48175 7175 48231
rect 7261 48175 7317 48231
rect 7403 48175 7459 48231
rect 7545 48175 7601 48231
rect 7687 48175 7743 48231
rect 7829 48175 7885 48231
rect 7971 48175 8027 48231
rect 8113 48175 8169 48231
rect 8255 48175 8311 48231
rect 8397 48175 8453 48231
rect 8539 48175 8595 48231
rect 8681 48175 8737 48231
rect 8823 48175 8879 48231
rect 8965 48175 9021 48231
rect 9107 48175 9163 48231
rect 9249 48175 9305 48231
rect 9391 48175 9447 48231
rect 9533 48175 9589 48231
rect 9675 48175 9731 48231
rect 9817 48175 9873 48231
rect 9959 48175 10015 48231
rect 10101 48175 10157 48231
rect 10243 48175 10299 48231
rect 10385 48175 10441 48231
rect 10527 48175 10583 48231
rect 10669 48175 10725 48231
rect 10811 48175 10867 48231
rect 10953 48175 11009 48231
rect 11095 48175 11151 48231
rect 11237 48175 11293 48231
rect 11379 48175 11435 48231
rect 11521 48175 11577 48231
rect 11663 48175 11719 48231
rect 11805 48175 11861 48231
rect 11947 48175 12003 48231
rect 12089 48175 12145 48231
rect 12231 48175 12287 48231
rect 12373 48175 12429 48231
rect 12515 48175 12571 48231
rect 12657 48175 12713 48231
rect 12799 48175 12855 48231
rect 12941 48175 12997 48231
rect 13083 48175 13139 48231
rect 13225 48175 13281 48231
rect 13367 48175 13423 48231
rect 13509 48175 13565 48231
rect 13651 48175 13707 48231
rect 13793 48175 13849 48231
rect 13935 48175 13991 48231
rect 14077 48175 14133 48231
rect 14219 48175 14275 48231
rect 14361 48175 14417 48231
rect 14503 48175 14559 48231
rect 14645 48175 14701 48231
rect 14787 48175 14843 48231
rect 161 48033 217 48089
rect 303 48033 359 48089
rect 445 48033 501 48089
rect 587 48033 643 48089
rect 729 48033 785 48089
rect 871 48033 927 48089
rect 1013 48033 1069 48089
rect 1155 48033 1211 48089
rect 1297 48033 1353 48089
rect 1439 48033 1495 48089
rect 1581 48033 1637 48089
rect 1723 48033 1779 48089
rect 1865 48033 1921 48089
rect 2007 48033 2063 48089
rect 2149 48033 2205 48089
rect 2291 48033 2347 48089
rect 2433 48033 2489 48089
rect 2575 48033 2631 48089
rect 2717 48033 2773 48089
rect 2859 48033 2915 48089
rect 3001 48033 3057 48089
rect 3143 48033 3199 48089
rect 3285 48033 3341 48089
rect 3427 48033 3483 48089
rect 3569 48033 3625 48089
rect 3711 48033 3767 48089
rect 3853 48033 3909 48089
rect 3995 48033 4051 48089
rect 4137 48033 4193 48089
rect 4279 48033 4335 48089
rect 4421 48033 4477 48089
rect 4563 48033 4619 48089
rect 4705 48033 4761 48089
rect 4847 48033 4903 48089
rect 4989 48033 5045 48089
rect 5131 48033 5187 48089
rect 5273 48033 5329 48089
rect 5415 48033 5471 48089
rect 5557 48033 5613 48089
rect 5699 48033 5755 48089
rect 5841 48033 5897 48089
rect 5983 48033 6039 48089
rect 6125 48033 6181 48089
rect 6267 48033 6323 48089
rect 6409 48033 6465 48089
rect 6551 48033 6607 48089
rect 6693 48033 6749 48089
rect 6835 48033 6891 48089
rect 6977 48033 7033 48089
rect 7119 48033 7175 48089
rect 7261 48033 7317 48089
rect 7403 48033 7459 48089
rect 7545 48033 7601 48089
rect 7687 48033 7743 48089
rect 7829 48033 7885 48089
rect 7971 48033 8027 48089
rect 8113 48033 8169 48089
rect 8255 48033 8311 48089
rect 8397 48033 8453 48089
rect 8539 48033 8595 48089
rect 8681 48033 8737 48089
rect 8823 48033 8879 48089
rect 8965 48033 9021 48089
rect 9107 48033 9163 48089
rect 9249 48033 9305 48089
rect 9391 48033 9447 48089
rect 9533 48033 9589 48089
rect 9675 48033 9731 48089
rect 9817 48033 9873 48089
rect 9959 48033 10015 48089
rect 10101 48033 10157 48089
rect 10243 48033 10299 48089
rect 10385 48033 10441 48089
rect 10527 48033 10583 48089
rect 10669 48033 10725 48089
rect 10811 48033 10867 48089
rect 10953 48033 11009 48089
rect 11095 48033 11151 48089
rect 11237 48033 11293 48089
rect 11379 48033 11435 48089
rect 11521 48033 11577 48089
rect 11663 48033 11719 48089
rect 11805 48033 11861 48089
rect 11947 48033 12003 48089
rect 12089 48033 12145 48089
rect 12231 48033 12287 48089
rect 12373 48033 12429 48089
rect 12515 48033 12571 48089
rect 12657 48033 12713 48089
rect 12799 48033 12855 48089
rect 12941 48033 12997 48089
rect 13083 48033 13139 48089
rect 13225 48033 13281 48089
rect 13367 48033 13423 48089
rect 13509 48033 13565 48089
rect 13651 48033 13707 48089
rect 13793 48033 13849 48089
rect 13935 48033 13991 48089
rect 14077 48033 14133 48089
rect 14219 48033 14275 48089
rect 14361 48033 14417 48089
rect 14503 48033 14559 48089
rect 14645 48033 14701 48089
rect 14787 48033 14843 48089
rect 161 47891 217 47947
rect 303 47891 359 47947
rect 445 47891 501 47947
rect 587 47891 643 47947
rect 729 47891 785 47947
rect 871 47891 927 47947
rect 1013 47891 1069 47947
rect 1155 47891 1211 47947
rect 1297 47891 1353 47947
rect 1439 47891 1495 47947
rect 1581 47891 1637 47947
rect 1723 47891 1779 47947
rect 1865 47891 1921 47947
rect 2007 47891 2063 47947
rect 2149 47891 2205 47947
rect 2291 47891 2347 47947
rect 2433 47891 2489 47947
rect 2575 47891 2631 47947
rect 2717 47891 2773 47947
rect 2859 47891 2915 47947
rect 3001 47891 3057 47947
rect 3143 47891 3199 47947
rect 3285 47891 3341 47947
rect 3427 47891 3483 47947
rect 3569 47891 3625 47947
rect 3711 47891 3767 47947
rect 3853 47891 3909 47947
rect 3995 47891 4051 47947
rect 4137 47891 4193 47947
rect 4279 47891 4335 47947
rect 4421 47891 4477 47947
rect 4563 47891 4619 47947
rect 4705 47891 4761 47947
rect 4847 47891 4903 47947
rect 4989 47891 5045 47947
rect 5131 47891 5187 47947
rect 5273 47891 5329 47947
rect 5415 47891 5471 47947
rect 5557 47891 5613 47947
rect 5699 47891 5755 47947
rect 5841 47891 5897 47947
rect 5983 47891 6039 47947
rect 6125 47891 6181 47947
rect 6267 47891 6323 47947
rect 6409 47891 6465 47947
rect 6551 47891 6607 47947
rect 6693 47891 6749 47947
rect 6835 47891 6891 47947
rect 6977 47891 7033 47947
rect 7119 47891 7175 47947
rect 7261 47891 7317 47947
rect 7403 47891 7459 47947
rect 7545 47891 7601 47947
rect 7687 47891 7743 47947
rect 7829 47891 7885 47947
rect 7971 47891 8027 47947
rect 8113 47891 8169 47947
rect 8255 47891 8311 47947
rect 8397 47891 8453 47947
rect 8539 47891 8595 47947
rect 8681 47891 8737 47947
rect 8823 47891 8879 47947
rect 8965 47891 9021 47947
rect 9107 47891 9163 47947
rect 9249 47891 9305 47947
rect 9391 47891 9447 47947
rect 9533 47891 9589 47947
rect 9675 47891 9731 47947
rect 9817 47891 9873 47947
rect 9959 47891 10015 47947
rect 10101 47891 10157 47947
rect 10243 47891 10299 47947
rect 10385 47891 10441 47947
rect 10527 47891 10583 47947
rect 10669 47891 10725 47947
rect 10811 47891 10867 47947
rect 10953 47891 11009 47947
rect 11095 47891 11151 47947
rect 11237 47891 11293 47947
rect 11379 47891 11435 47947
rect 11521 47891 11577 47947
rect 11663 47891 11719 47947
rect 11805 47891 11861 47947
rect 11947 47891 12003 47947
rect 12089 47891 12145 47947
rect 12231 47891 12287 47947
rect 12373 47891 12429 47947
rect 12515 47891 12571 47947
rect 12657 47891 12713 47947
rect 12799 47891 12855 47947
rect 12941 47891 12997 47947
rect 13083 47891 13139 47947
rect 13225 47891 13281 47947
rect 13367 47891 13423 47947
rect 13509 47891 13565 47947
rect 13651 47891 13707 47947
rect 13793 47891 13849 47947
rect 13935 47891 13991 47947
rect 14077 47891 14133 47947
rect 14219 47891 14275 47947
rect 14361 47891 14417 47947
rect 14503 47891 14559 47947
rect 14645 47891 14701 47947
rect 14787 47891 14843 47947
rect 161 47749 217 47805
rect 303 47749 359 47805
rect 445 47749 501 47805
rect 587 47749 643 47805
rect 729 47749 785 47805
rect 871 47749 927 47805
rect 1013 47749 1069 47805
rect 1155 47749 1211 47805
rect 1297 47749 1353 47805
rect 1439 47749 1495 47805
rect 1581 47749 1637 47805
rect 1723 47749 1779 47805
rect 1865 47749 1921 47805
rect 2007 47749 2063 47805
rect 2149 47749 2205 47805
rect 2291 47749 2347 47805
rect 2433 47749 2489 47805
rect 2575 47749 2631 47805
rect 2717 47749 2773 47805
rect 2859 47749 2915 47805
rect 3001 47749 3057 47805
rect 3143 47749 3199 47805
rect 3285 47749 3341 47805
rect 3427 47749 3483 47805
rect 3569 47749 3625 47805
rect 3711 47749 3767 47805
rect 3853 47749 3909 47805
rect 3995 47749 4051 47805
rect 4137 47749 4193 47805
rect 4279 47749 4335 47805
rect 4421 47749 4477 47805
rect 4563 47749 4619 47805
rect 4705 47749 4761 47805
rect 4847 47749 4903 47805
rect 4989 47749 5045 47805
rect 5131 47749 5187 47805
rect 5273 47749 5329 47805
rect 5415 47749 5471 47805
rect 5557 47749 5613 47805
rect 5699 47749 5755 47805
rect 5841 47749 5897 47805
rect 5983 47749 6039 47805
rect 6125 47749 6181 47805
rect 6267 47749 6323 47805
rect 6409 47749 6465 47805
rect 6551 47749 6607 47805
rect 6693 47749 6749 47805
rect 6835 47749 6891 47805
rect 6977 47749 7033 47805
rect 7119 47749 7175 47805
rect 7261 47749 7317 47805
rect 7403 47749 7459 47805
rect 7545 47749 7601 47805
rect 7687 47749 7743 47805
rect 7829 47749 7885 47805
rect 7971 47749 8027 47805
rect 8113 47749 8169 47805
rect 8255 47749 8311 47805
rect 8397 47749 8453 47805
rect 8539 47749 8595 47805
rect 8681 47749 8737 47805
rect 8823 47749 8879 47805
rect 8965 47749 9021 47805
rect 9107 47749 9163 47805
rect 9249 47749 9305 47805
rect 9391 47749 9447 47805
rect 9533 47749 9589 47805
rect 9675 47749 9731 47805
rect 9817 47749 9873 47805
rect 9959 47749 10015 47805
rect 10101 47749 10157 47805
rect 10243 47749 10299 47805
rect 10385 47749 10441 47805
rect 10527 47749 10583 47805
rect 10669 47749 10725 47805
rect 10811 47749 10867 47805
rect 10953 47749 11009 47805
rect 11095 47749 11151 47805
rect 11237 47749 11293 47805
rect 11379 47749 11435 47805
rect 11521 47749 11577 47805
rect 11663 47749 11719 47805
rect 11805 47749 11861 47805
rect 11947 47749 12003 47805
rect 12089 47749 12145 47805
rect 12231 47749 12287 47805
rect 12373 47749 12429 47805
rect 12515 47749 12571 47805
rect 12657 47749 12713 47805
rect 12799 47749 12855 47805
rect 12941 47749 12997 47805
rect 13083 47749 13139 47805
rect 13225 47749 13281 47805
rect 13367 47749 13423 47805
rect 13509 47749 13565 47805
rect 13651 47749 13707 47805
rect 13793 47749 13849 47805
rect 13935 47749 13991 47805
rect 14077 47749 14133 47805
rect 14219 47749 14275 47805
rect 14361 47749 14417 47805
rect 14503 47749 14559 47805
rect 14645 47749 14701 47805
rect 14787 47749 14843 47805
rect 161 47607 217 47663
rect 303 47607 359 47663
rect 445 47607 501 47663
rect 587 47607 643 47663
rect 729 47607 785 47663
rect 871 47607 927 47663
rect 1013 47607 1069 47663
rect 1155 47607 1211 47663
rect 1297 47607 1353 47663
rect 1439 47607 1495 47663
rect 1581 47607 1637 47663
rect 1723 47607 1779 47663
rect 1865 47607 1921 47663
rect 2007 47607 2063 47663
rect 2149 47607 2205 47663
rect 2291 47607 2347 47663
rect 2433 47607 2489 47663
rect 2575 47607 2631 47663
rect 2717 47607 2773 47663
rect 2859 47607 2915 47663
rect 3001 47607 3057 47663
rect 3143 47607 3199 47663
rect 3285 47607 3341 47663
rect 3427 47607 3483 47663
rect 3569 47607 3625 47663
rect 3711 47607 3767 47663
rect 3853 47607 3909 47663
rect 3995 47607 4051 47663
rect 4137 47607 4193 47663
rect 4279 47607 4335 47663
rect 4421 47607 4477 47663
rect 4563 47607 4619 47663
rect 4705 47607 4761 47663
rect 4847 47607 4903 47663
rect 4989 47607 5045 47663
rect 5131 47607 5187 47663
rect 5273 47607 5329 47663
rect 5415 47607 5471 47663
rect 5557 47607 5613 47663
rect 5699 47607 5755 47663
rect 5841 47607 5897 47663
rect 5983 47607 6039 47663
rect 6125 47607 6181 47663
rect 6267 47607 6323 47663
rect 6409 47607 6465 47663
rect 6551 47607 6607 47663
rect 6693 47607 6749 47663
rect 6835 47607 6891 47663
rect 6977 47607 7033 47663
rect 7119 47607 7175 47663
rect 7261 47607 7317 47663
rect 7403 47607 7459 47663
rect 7545 47607 7601 47663
rect 7687 47607 7743 47663
rect 7829 47607 7885 47663
rect 7971 47607 8027 47663
rect 8113 47607 8169 47663
rect 8255 47607 8311 47663
rect 8397 47607 8453 47663
rect 8539 47607 8595 47663
rect 8681 47607 8737 47663
rect 8823 47607 8879 47663
rect 8965 47607 9021 47663
rect 9107 47607 9163 47663
rect 9249 47607 9305 47663
rect 9391 47607 9447 47663
rect 9533 47607 9589 47663
rect 9675 47607 9731 47663
rect 9817 47607 9873 47663
rect 9959 47607 10015 47663
rect 10101 47607 10157 47663
rect 10243 47607 10299 47663
rect 10385 47607 10441 47663
rect 10527 47607 10583 47663
rect 10669 47607 10725 47663
rect 10811 47607 10867 47663
rect 10953 47607 11009 47663
rect 11095 47607 11151 47663
rect 11237 47607 11293 47663
rect 11379 47607 11435 47663
rect 11521 47607 11577 47663
rect 11663 47607 11719 47663
rect 11805 47607 11861 47663
rect 11947 47607 12003 47663
rect 12089 47607 12145 47663
rect 12231 47607 12287 47663
rect 12373 47607 12429 47663
rect 12515 47607 12571 47663
rect 12657 47607 12713 47663
rect 12799 47607 12855 47663
rect 12941 47607 12997 47663
rect 13083 47607 13139 47663
rect 13225 47607 13281 47663
rect 13367 47607 13423 47663
rect 13509 47607 13565 47663
rect 13651 47607 13707 47663
rect 13793 47607 13849 47663
rect 13935 47607 13991 47663
rect 14077 47607 14133 47663
rect 14219 47607 14275 47663
rect 14361 47607 14417 47663
rect 14503 47607 14559 47663
rect 14645 47607 14701 47663
rect 14787 47607 14843 47663
rect 161 47465 217 47521
rect 303 47465 359 47521
rect 445 47465 501 47521
rect 587 47465 643 47521
rect 729 47465 785 47521
rect 871 47465 927 47521
rect 1013 47465 1069 47521
rect 1155 47465 1211 47521
rect 1297 47465 1353 47521
rect 1439 47465 1495 47521
rect 1581 47465 1637 47521
rect 1723 47465 1779 47521
rect 1865 47465 1921 47521
rect 2007 47465 2063 47521
rect 2149 47465 2205 47521
rect 2291 47465 2347 47521
rect 2433 47465 2489 47521
rect 2575 47465 2631 47521
rect 2717 47465 2773 47521
rect 2859 47465 2915 47521
rect 3001 47465 3057 47521
rect 3143 47465 3199 47521
rect 3285 47465 3341 47521
rect 3427 47465 3483 47521
rect 3569 47465 3625 47521
rect 3711 47465 3767 47521
rect 3853 47465 3909 47521
rect 3995 47465 4051 47521
rect 4137 47465 4193 47521
rect 4279 47465 4335 47521
rect 4421 47465 4477 47521
rect 4563 47465 4619 47521
rect 4705 47465 4761 47521
rect 4847 47465 4903 47521
rect 4989 47465 5045 47521
rect 5131 47465 5187 47521
rect 5273 47465 5329 47521
rect 5415 47465 5471 47521
rect 5557 47465 5613 47521
rect 5699 47465 5755 47521
rect 5841 47465 5897 47521
rect 5983 47465 6039 47521
rect 6125 47465 6181 47521
rect 6267 47465 6323 47521
rect 6409 47465 6465 47521
rect 6551 47465 6607 47521
rect 6693 47465 6749 47521
rect 6835 47465 6891 47521
rect 6977 47465 7033 47521
rect 7119 47465 7175 47521
rect 7261 47465 7317 47521
rect 7403 47465 7459 47521
rect 7545 47465 7601 47521
rect 7687 47465 7743 47521
rect 7829 47465 7885 47521
rect 7971 47465 8027 47521
rect 8113 47465 8169 47521
rect 8255 47465 8311 47521
rect 8397 47465 8453 47521
rect 8539 47465 8595 47521
rect 8681 47465 8737 47521
rect 8823 47465 8879 47521
rect 8965 47465 9021 47521
rect 9107 47465 9163 47521
rect 9249 47465 9305 47521
rect 9391 47465 9447 47521
rect 9533 47465 9589 47521
rect 9675 47465 9731 47521
rect 9817 47465 9873 47521
rect 9959 47465 10015 47521
rect 10101 47465 10157 47521
rect 10243 47465 10299 47521
rect 10385 47465 10441 47521
rect 10527 47465 10583 47521
rect 10669 47465 10725 47521
rect 10811 47465 10867 47521
rect 10953 47465 11009 47521
rect 11095 47465 11151 47521
rect 11237 47465 11293 47521
rect 11379 47465 11435 47521
rect 11521 47465 11577 47521
rect 11663 47465 11719 47521
rect 11805 47465 11861 47521
rect 11947 47465 12003 47521
rect 12089 47465 12145 47521
rect 12231 47465 12287 47521
rect 12373 47465 12429 47521
rect 12515 47465 12571 47521
rect 12657 47465 12713 47521
rect 12799 47465 12855 47521
rect 12941 47465 12997 47521
rect 13083 47465 13139 47521
rect 13225 47465 13281 47521
rect 13367 47465 13423 47521
rect 13509 47465 13565 47521
rect 13651 47465 13707 47521
rect 13793 47465 13849 47521
rect 13935 47465 13991 47521
rect 14077 47465 14133 47521
rect 14219 47465 14275 47521
rect 14361 47465 14417 47521
rect 14503 47465 14559 47521
rect 14645 47465 14701 47521
rect 14787 47465 14843 47521
rect 161 47323 217 47379
rect 303 47323 359 47379
rect 445 47323 501 47379
rect 587 47323 643 47379
rect 729 47323 785 47379
rect 871 47323 927 47379
rect 1013 47323 1069 47379
rect 1155 47323 1211 47379
rect 1297 47323 1353 47379
rect 1439 47323 1495 47379
rect 1581 47323 1637 47379
rect 1723 47323 1779 47379
rect 1865 47323 1921 47379
rect 2007 47323 2063 47379
rect 2149 47323 2205 47379
rect 2291 47323 2347 47379
rect 2433 47323 2489 47379
rect 2575 47323 2631 47379
rect 2717 47323 2773 47379
rect 2859 47323 2915 47379
rect 3001 47323 3057 47379
rect 3143 47323 3199 47379
rect 3285 47323 3341 47379
rect 3427 47323 3483 47379
rect 3569 47323 3625 47379
rect 3711 47323 3767 47379
rect 3853 47323 3909 47379
rect 3995 47323 4051 47379
rect 4137 47323 4193 47379
rect 4279 47323 4335 47379
rect 4421 47323 4477 47379
rect 4563 47323 4619 47379
rect 4705 47323 4761 47379
rect 4847 47323 4903 47379
rect 4989 47323 5045 47379
rect 5131 47323 5187 47379
rect 5273 47323 5329 47379
rect 5415 47323 5471 47379
rect 5557 47323 5613 47379
rect 5699 47323 5755 47379
rect 5841 47323 5897 47379
rect 5983 47323 6039 47379
rect 6125 47323 6181 47379
rect 6267 47323 6323 47379
rect 6409 47323 6465 47379
rect 6551 47323 6607 47379
rect 6693 47323 6749 47379
rect 6835 47323 6891 47379
rect 6977 47323 7033 47379
rect 7119 47323 7175 47379
rect 7261 47323 7317 47379
rect 7403 47323 7459 47379
rect 7545 47323 7601 47379
rect 7687 47323 7743 47379
rect 7829 47323 7885 47379
rect 7971 47323 8027 47379
rect 8113 47323 8169 47379
rect 8255 47323 8311 47379
rect 8397 47323 8453 47379
rect 8539 47323 8595 47379
rect 8681 47323 8737 47379
rect 8823 47323 8879 47379
rect 8965 47323 9021 47379
rect 9107 47323 9163 47379
rect 9249 47323 9305 47379
rect 9391 47323 9447 47379
rect 9533 47323 9589 47379
rect 9675 47323 9731 47379
rect 9817 47323 9873 47379
rect 9959 47323 10015 47379
rect 10101 47323 10157 47379
rect 10243 47323 10299 47379
rect 10385 47323 10441 47379
rect 10527 47323 10583 47379
rect 10669 47323 10725 47379
rect 10811 47323 10867 47379
rect 10953 47323 11009 47379
rect 11095 47323 11151 47379
rect 11237 47323 11293 47379
rect 11379 47323 11435 47379
rect 11521 47323 11577 47379
rect 11663 47323 11719 47379
rect 11805 47323 11861 47379
rect 11947 47323 12003 47379
rect 12089 47323 12145 47379
rect 12231 47323 12287 47379
rect 12373 47323 12429 47379
rect 12515 47323 12571 47379
rect 12657 47323 12713 47379
rect 12799 47323 12855 47379
rect 12941 47323 12997 47379
rect 13083 47323 13139 47379
rect 13225 47323 13281 47379
rect 13367 47323 13423 47379
rect 13509 47323 13565 47379
rect 13651 47323 13707 47379
rect 13793 47323 13849 47379
rect 13935 47323 13991 47379
rect 14077 47323 14133 47379
rect 14219 47323 14275 47379
rect 14361 47323 14417 47379
rect 14503 47323 14559 47379
rect 14645 47323 14701 47379
rect 14787 47323 14843 47379
rect 161 47181 217 47237
rect 303 47181 359 47237
rect 445 47181 501 47237
rect 587 47181 643 47237
rect 729 47181 785 47237
rect 871 47181 927 47237
rect 1013 47181 1069 47237
rect 1155 47181 1211 47237
rect 1297 47181 1353 47237
rect 1439 47181 1495 47237
rect 1581 47181 1637 47237
rect 1723 47181 1779 47237
rect 1865 47181 1921 47237
rect 2007 47181 2063 47237
rect 2149 47181 2205 47237
rect 2291 47181 2347 47237
rect 2433 47181 2489 47237
rect 2575 47181 2631 47237
rect 2717 47181 2773 47237
rect 2859 47181 2915 47237
rect 3001 47181 3057 47237
rect 3143 47181 3199 47237
rect 3285 47181 3341 47237
rect 3427 47181 3483 47237
rect 3569 47181 3625 47237
rect 3711 47181 3767 47237
rect 3853 47181 3909 47237
rect 3995 47181 4051 47237
rect 4137 47181 4193 47237
rect 4279 47181 4335 47237
rect 4421 47181 4477 47237
rect 4563 47181 4619 47237
rect 4705 47181 4761 47237
rect 4847 47181 4903 47237
rect 4989 47181 5045 47237
rect 5131 47181 5187 47237
rect 5273 47181 5329 47237
rect 5415 47181 5471 47237
rect 5557 47181 5613 47237
rect 5699 47181 5755 47237
rect 5841 47181 5897 47237
rect 5983 47181 6039 47237
rect 6125 47181 6181 47237
rect 6267 47181 6323 47237
rect 6409 47181 6465 47237
rect 6551 47181 6607 47237
rect 6693 47181 6749 47237
rect 6835 47181 6891 47237
rect 6977 47181 7033 47237
rect 7119 47181 7175 47237
rect 7261 47181 7317 47237
rect 7403 47181 7459 47237
rect 7545 47181 7601 47237
rect 7687 47181 7743 47237
rect 7829 47181 7885 47237
rect 7971 47181 8027 47237
rect 8113 47181 8169 47237
rect 8255 47181 8311 47237
rect 8397 47181 8453 47237
rect 8539 47181 8595 47237
rect 8681 47181 8737 47237
rect 8823 47181 8879 47237
rect 8965 47181 9021 47237
rect 9107 47181 9163 47237
rect 9249 47181 9305 47237
rect 9391 47181 9447 47237
rect 9533 47181 9589 47237
rect 9675 47181 9731 47237
rect 9817 47181 9873 47237
rect 9959 47181 10015 47237
rect 10101 47181 10157 47237
rect 10243 47181 10299 47237
rect 10385 47181 10441 47237
rect 10527 47181 10583 47237
rect 10669 47181 10725 47237
rect 10811 47181 10867 47237
rect 10953 47181 11009 47237
rect 11095 47181 11151 47237
rect 11237 47181 11293 47237
rect 11379 47181 11435 47237
rect 11521 47181 11577 47237
rect 11663 47181 11719 47237
rect 11805 47181 11861 47237
rect 11947 47181 12003 47237
rect 12089 47181 12145 47237
rect 12231 47181 12287 47237
rect 12373 47181 12429 47237
rect 12515 47181 12571 47237
rect 12657 47181 12713 47237
rect 12799 47181 12855 47237
rect 12941 47181 12997 47237
rect 13083 47181 13139 47237
rect 13225 47181 13281 47237
rect 13367 47181 13423 47237
rect 13509 47181 13565 47237
rect 13651 47181 13707 47237
rect 13793 47181 13849 47237
rect 13935 47181 13991 47237
rect 14077 47181 14133 47237
rect 14219 47181 14275 47237
rect 14361 47181 14417 47237
rect 14503 47181 14559 47237
rect 14645 47181 14701 47237
rect 14787 47181 14843 47237
rect 161 47039 217 47095
rect 303 47039 359 47095
rect 445 47039 501 47095
rect 587 47039 643 47095
rect 729 47039 785 47095
rect 871 47039 927 47095
rect 1013 47039 1069 47095
rect 1155 47039 1211 47095
rect 1297 47039 1353 47095
rect 1439 47039 1495 47095
rect 1581 47039 1637 47095
rect 1723 47039 1779 47095
rect 1865 47039 1921 47095
rect 2007 47039 2063 47095
rect 2149 47039 2205 47095
rect 2291 47039 2347 47095
rect 2433 47039 2489 47095
rect 2575 47039 2631 47095
rect 2717 47039 2773 47095
rect 2859 47039 2915 47095
rect 3001 47039 3057 47095
rect 3143 47039 3199 47095
rect 3285 47039 3341 47095
rect 3427 47039 3483 47095
rect 3569 47039 3625 47095
rect 3711 47039 3767 47095
rect 3853 47039 3909 47095
rect 3995 47039 4051 47095
rect 4137 47039 4193 47095
rect 4279 47039 4335 47095
rect 4421 47039 4477 47095
rect 4563 47039 4619 47095
rect 4705 47039 4761 47095
rect 4847 47039 4903 47095
rect 4989 47039 5045 47095
rect 5131 47039 5187 47095
rect 5273 47039 5329 47095
rect 5415 47039 5471 47095
rect 5557 47039 5613 47095
rect 5699 47039 5755 47095
rect 5841 47039 5897 47095
rect 5983 47039 6039 47095
rect 6125 47039 6181 47095
rect 6267 47039 6323 47095
rect 6409 47039 6465 47095
rect 6551 47039 6607 47095
rect 6693 47039 6749 47095
rect 6835 47039 6891 47095
rect 6977 47039 7033 47095
rect 7119 47039 7175 47095
rect 7261 47039 7317 47095
rect 7403 47039 7459 47095
rect 7545 47039 7601 47095
rect 7687 47039 7743 47095
rect 7829 47039 7885 47095
rect 7971 47039 8027 47095
rect 8113 47039 8169 47095
rect 8255 47039 8311 47095
rect 8397 47039 8453 47095
rect 8539 47039 8595 47095
rect 8681 47039 8737 47095
rect 8823 47039 8879 47095
rect 8965 47039 9021 47095
rect 9107 47039 9163 47095
rect 9249 47039 9305 47095
rect 9391 47039 9447 47095
rect 9533 47039 9589 47095
rect 9675 47039 9731 47095
rect 9817 47039 9873 47095
rect 9959 47039 10015 47095
rect 10101 47039 10157 47095
rect 10243 47039 10299 47095
rect 10385 47039 10441 47095
rect 10527 47039 10583 47095
rect 10669 47039 10725 47095
rect 10811 47039 10867 47095
rect 10953 47039 11009 47095
rect 11095 47039 11151 47095
rect 11237 47039 11293 47095
rect 11379 47039 11435 47095
rect 11521 47039 11577 47095
rect 11663 47039 11719 47095
rect 11805 47039 11861 47095
rect 11947 47039 12003 47095
rect 12089 47039 12145 47095
rect 12231 47039 12287 47095
rect 12373 47039 12429 47095
rect 12515 47039 12571 47095
rect 12657 47039 12713 47095
rect 12799 47039 12855 47095
rect 12941 47039 12997 47095
rect 13083 47039 13139 47095
rect 13225 47039 13281 47095
rect 13367 47039 13423 47095
rect 13509 47039 13565 47095
rect 13651 47039 13707 47095
rect 13793 47039 13849 47095
rect 13935 47039 13991 47095
rect 14077 47039 14133 47095
rect 14219 47039 14275 47095
rect 14361 47039 14417 47095
rect 14503 47039 14559 47095
rect 14645 47039 14701 47095
rect 14787 47039 14843 47095
rect 161 46897 217 46953
rect 303 46897 359 46953
rect 445 46897 501 46953
rect 587 46897 643 46953
rect 729 46897 785 46953
rect 871 46897 927 46953
rect 1013 46897 1069 46953
rect 1155 46897 1211 46953
rect 1297 46897 1353 46953
rect 1439 46897 1495 46953
rect 1581 46897 1637 46953
rect 1723 46897 1779 46953
rect 1865 46897 1921 46953
rect 2007 46897 2063 46953
rect 2149 46897 2205 46953
rect 2291 46897 2347 46953
rect 2433 46897 2489 46953
rect 2575 46897 2631 46953
rect 2717 46897 2773 46953
rect 2859 46897 2915 46953
rect 3001 46897 3057 46953
rect 3143 46897 3199 46953
rect 3285 46897 3341 46953
rect 3427 46897 3483 46953
rect 3569 46897 3625 46953
rect 3711 46897 3767 46953
rect 3853 46897 3909 46953
rect 3995 46897 4051 46953
rect 4137 46897 4193 46953
rect 4279 46897 4335 46953
rect 4421 46897 4477 46953
rect 4563 46897 4619 46953
rect 4705 46897 4761 46953
rect 4847 46897 4903 46953
rect 4989 46897 5045 46953
rect 5131 46897 5187 46953
rect 5273 46897 5329 46953
rect 5415 46897 5471 46953
rect 5557 46897 5613 46953
rect 5699 46897 5755 46953
rect 5841 46897 5897 46953
rect 5983 46897 6039 46953
rect 6125 46897 6181 46953
rect 6267 46897 6323 46953
rect 6409 46897 6465 46953
rect 6551 46897 6607 46953
rect 6693 46897 6749 46953
rect 6835 46897 6891 46953
rect 6977 46897 7033 46953
rect 7119 46897 7175 46953
rect 7261 46897 7317 46953
rect 7403 46897 7459 46953
rect 7545 46897 7601 46953
rect 7687 46897 7743 46953
rect 7829 46897 7885 46953
rect 7971 46897 8027 46953
rect 8113 46897 8169 46953
rect 8255 46897 8311 46953
rect 8397 46897 8453 46953
rect 8539 46897 8595 46953
rect 8681 46897 8737 46953
rect 8823 46897 8879 46953
rect 8965 46897 9021 46953
rect 9107 46897 9163 46953
rect 9249 46897 9305 46953
rect 9391 46897 9447 46953
rect 9533 46897 9589 46953
rect 9675 46897 9731 46953
rect 9817 46897 9873 46953
rect 9959 46897 10015 46953
rect 10101 46897 10157 46953
rect 10243 46897 10299 46953
rect 10385 46897 10441 46953
rect 10527 46897 10583 46953
rect 10669 46897 10725 46953
rect 10811 46897 10867 46953
rect 10953 46897 11009 46953
rect 11095 46897 11151 46953
rect 11237 46897 11293 46953
rect 11379 46897 11435 46953
rect 11521 46897 11577 46953
rect 11663 46897 11719 46953
rect 11805 46897 11861 46953
rect 11947 46897 12003 46953
rect 12089 46897 12145 46953
rect 12231 46897 12287 46953
rect 12373 46897 12429 46953
rect 12515 46897 12571 46953
rect 12657 46897 12713 46953
rect 12799 46897 12855 46953
rect 12941 46897 12997 46953
rect 13083 46897 13139 46953
rect 13225 46897 13281 46953
rect 13367 46897 13423 46953
rect 13509 46897 13565 46953
rect 13651 46897 13707 46953
rect 13793 46897 13849 46953
rect 13935 46897 13991 46953
rect 14077 46897 14133 46953
rect 14219 46897 14275 46953
rect 14361 46897 14417 46953
rect 14503 46897 14559 46953
rect 14645 46897 14701 46953
rect 14787 46897 14843 46953
rect 161 46755 217 46811
rect 303 46755 359 46811
rect 445 46755 501 46811
rect 587 46755 643 46811
rect 729 46755 785 46811
rect 871 46755 927 46811
rect 1013 46755 1069 46811
rect 1155 46755 1211 46811
rect 1297 46755 1353 46811
rect 1439 46755 1495 46811
rect 1581 46755 1637 46811
rect 1723 46755 1779 46811
rect 1865 46755 1921 46811
rect 2007 46755 2063 46811
rect 2149 46755 2205 46811
rect 2291 46755 2347 46811
rect 2433 46755 2489 46811
rect 2575 46755 2631 46811
rect 2717 46755 2773 46811
rect 2859 46755 2915 46811
rect 3001 46755 3057 46811
rect 3143 46755 3199 46811
rect 3285 46755 3341 46811
rect 3427 46755 3483 46811
rect 3569 46755 3625 46811
rect 3711 46755 3767 46811
rect 3853 46755 3909 46811
rect 3995 46755 4051 46811
rect 4137 46755 4193 46811
rect 4279 46755 4335 46811
rect 4421 46755 4477 46811
rect 4563 46755 4619 46811
rect 4705 46755 4761 46811
rect 4847 46755 4903 46811
rect 4989 46755 5045 46811
rect 5131 46755 5187 46811
rect 5273 46755 5329 46811
rect 5415 46755 5471 46811
rect 5557 46755 5613 46811
rect 5699 46755 5755 46811
rect 5841 46755 5897 46811
rect 5983 46755 6039 46811
rect 6125 46755 6181 46811
rect 6267 46755 6323 46811
rect 6409 46755 6465 46811
rect 6551 46755 6607 46811
rect 6693 46755 6749 46811
rect 6835 46755 6891 46811
rect 6977 46755 7033 46811
rect 7119 46755 7175 46811
rect 7261 46755 7317 46811
rect 7403 46755 7459 46811
rect 7545 46755 7601 46811
rect 7687 46755 7743 46811
rect 7829 46755 7885 46811
rect 7971 46755 8027 46811
rect 8113 46755 8169 46811
rect 8255 46755 8311 46811
rect 8397 46755 8453 46811
rect 8539 46755 8595 46811
rect 8681 46755 8737 46811
rect 8823 46755 8879 46811
rect 8965 46755 9021 46811
rect 9107 46755 9163 46811
rect 9249 46755 9305 46811
rect 9391 46755 9447 46811
rect 9533 46755 9589 46811
rect 9675 46755 9731 46811
rect 9817 46755 9873 46811
rect 9959 46755 10015 46811
rect 10101 46755 10157 46811
rect 10243 46755 10299 46811
rect 10385 46755 10441 46811
rect 10527 46755 10583 46811
rect 10669 46755 10725 46811
rect 10811 46755 10867 46811
rect 10953 46755 11009 46811
rect 11095 46755 11151 46811
rect 11237 46755 11293 46811
rect 11379 46755 11435 46811
rect 11521 46755 11577 46811
rect 11663 46755 11719 46811
rect 11805 46755 11861 46811
rect 11947 46755 12003 46811
rect 12089 46755 12145 46811
rect 12231 46755 12287 46811
rect 12373 46755 12429 46811
rect 12515 46755 12571 46811
rect 12657 46755 12713 46811
rect 12799 46755 12855 46811
rect 12941 46755 12997 46811
rect 13083 46755 13139 46811
rect 13225 46755 13281 46811
rect 13367 46755 13423 46811
rect 13509 46755 13565 46811
rect 13651 46755 13707 46811
rect 13793 46755 13849 46811
rect 13935 46755 13991 46811
rect 14077 46755 14133 46811
rect 14219 46755 14275 46811
rect 14361 46755 14417 46811
rect 14503 46755 14559 46811
rect 14645 46755 14701 46811
rect 14787 46755 14843 46811
rect 161 46613 217 46669
rect 303 46613 359 46669
rect 445 46613 501 46669
rect 587 46613 643 46669
rect 729 46613 785 46669
rect 871 46613 927 46669
rect 1013 46613 1069 46669
rect 1155 46613 1211 46669
rect 1297 46613 1353 46669
rect 1439 46613 1495 46669
rect 1581 46613 1637 46669
rect 1723 46613 1779 46669
rect 1865 46613 1921 46669
rect 2007 46613 2063 46669
rect 2149 46613 2205 46669
rect 2291 46613 2347 46669
rect 2433 46613 2489 46669
rect 2575 46613 2631 46669
rect 2717 46613 2773 46669
rect 2859 46613 2915 46669
rect 3001 46613 3057 46669
rect 3143 46613 3199 46669
rect 3285 46613 3341 46669
rect 3427 46613 3483 46669
rect 3569 46613 3625 46669
rect 3711 46613 3767 46669
rect 3853 46613 3909 46669
rect 3995 46613 4051 46669
rect 4137 46613 4193 46669
rect 4279 46613 4335 46669
rect 4421 46613 4477 46669
rect 4563 46613 4619 46669
rect 4705 46613 4761 46669
rect 4847 46613 4903 46669
rect 4989 46613 5045 46669
rect 5131 46613 5187 46669
rect 5273 46613 5329 46669
rect 5415 46613 5471 46669
rect 5557 46613 5613 46669
rect 5699 46613 5755 46669
rect 5841 46613 5897 46669
rect 5983 46613 6039 46669
rect 6125 46613 6181 46669
rect 6267 46613 6323 46669
rect 6409 46613 6465 46669
rect 6551 46613 6607 46669
rect 6693 46613 6749 46669
rect 6835 46613 6891 46669
rect 6977 46613 7033 46669
rect 7119 46613 7175 46669
rect 7261 46613 7317 46669
rect 7403 46613 7459 46669
rect 7545 46613 7601 46669
rect 7687 46613 7743 46669
rect 7829 46613 7885 46669
rect 7971 46613 8027 46669
rect 8113 46613 8169 46669
rect 8255 46613 8311 46669
rect 8397 46613 8453 46669
rect 8539 46613 8595 46669
rect 8681 46613 8737 46669
rect 8823 46613 8879 46669
rect 8965 46613 9021 46669
rect 9107 46613 9163 46669
rect 9249 46613 9305 46669
rect 9391 46613 9447 46669
rect 9533 46613 9589 46669
rect 9675 46613 9731 46669
rect 9817 46613 9873 46669
rect 9959 46613 10015 46669
rect 10101 46613 10157 46669
rect 10243 46613 10299 46669
rect 10385 46613 10441 46669
rect 10527 46613 10583 46669
rect 10669 46613 10725 46669
rect 10811 46613 10867 46669
rect 10953 46613 11009 46669
rect 11095 46613 11151 46669
rect 11237 46613 11293 46669
rect 11379 46613 11435 46669
rect 11521 46613 11577 46669
rect 11663 46613 11719 46669
rect 11805 46613 11861 46669
rect 11947 46613 12003 46669
rect 12089 46613 12145 46669
rect 12231 46613 12287 46669
rect 12373 46613 12429 46669
rect 12515 46613 12571 46669
rect 12657 46613 12713 46669
rect 12799 46613 12855 46669
rect 12941 46613 12997 46669
rect 13083 46613 13139 46669
rect 13225 46613 13281 46669
rect 13367 46613 13423 46669
rect 13509 46613 13565 46669
rect 13651 46613 13707 46669
rect 13793 46613 13849 46669
rect 13935 46613 13991 46669
rect 14077 46613 14133 46669
rect 14219 46613 14275 46669
rect 14361 46613 14417 46669
rect 14503 46613 14559 46669
rect 14645 46613 14701 46669
rect 14787 46613 14843 46669
rect 161 46471 217 46527
rect 303 46471 359 46527
rect 445 46471 501 46527
rect 587 46471 643 46527
rect 729 46471 785 46527
rect 871 46471 927 46527
rect 1013 46471 1069 46527
rect 1155 46471 1211 46527
rect 1297 46471 1353 46527
rect 1439 46471 1495 46527
rect 1581 46471 1637 46527
rect 1723 46471 1779 46527
rect 1865 46471 1921 46527
rect 2007 46471 2063 46527
rect 2149 46471 2205 46527
rect 2291 46471 2347 46527
rect 2433 46471 2489 46527
rect 2575 46471 2631 46527
rect 2717 46471 2773 46527
rect 2859 46471 2915 46527
rect 3001 46471 3057 46527
rect 3143 46471 3199 46527
rect 3285 46471 3341 46527
rect 3427 46471 3483 46527
rect 3569 46471 3625 46527
rect 3711 46471 3767 46527
rect 3853 46471 3909 46527
rect 3995 46471 4051 46527
rect 4137 46471 4193 46527
rect 4279 46471 4335 46527
rect 4421 46471 4477 46527
rect 4563 46471 4619 46527
rect 4705 46471 4761 46527
rect 4847 46471 4903 46527
rect 4989 46471 5045 46527
rect 5131 46471 5187 46527
rect 5273 46471 5329 46527
rect 5415 46471 5471 46527
rect 5557 46471 5613 46527
rect 5699 46471 5755 46527
rect 5841 46471 5897 46527
rect 5983 46471 6039 46527
rect 6125 46471 6181 46527
rect 6267 46471 6323 46527
rect 6409 46471 6465 46527
rect 6551 46471 6607 46527
rect 6693 46471 6749 46527
rect 6835 46471 6891 46527
rect 6977 46471 7033 46527
rect 7119 46471 7175 46527
rect 7261 46471 7317 46527
rect 7403 46471 7459 46527
rect 7545 46471 7601 46527
rect 7687 46471 7743 46527
rect 7829 46471 7885 46527
rect 7971 46471 8027 46527
rect 8113 46471 8169 46527
rect 8255 46471 8311 46527
rect 8397 46471 8453 46527
rect 8539 46471 8595 46527
rect 8681 46471 8737 46527
rect 8823 46471 8879 46527
rect 8965 46471 9021 46527
rect 9107 46471 9163 46527
rect 9249 46471 9305 46527
rect 9391 46471 9447 46527
rect 9533 46471 9589 46527
rect 9675 46471 9731 46527
rect 9817 46471 9873 46527
rect 9959 46471 10015 46527
rect 10101 46471 10157 46527
rect 10243 46471 10299 46527
rect 10385 46471 10441 46527
rect 10527 46471 10583 46527
rect 10669 46471 10725 46527
rect 10811 46471 10867 46527
rect 10953 46471 11009 46527
rect 11095 46471 11151 46527
rect 11237 46471 11293 46527
rect 11379 46471 11435 46527
rect 11521 46471 11577 46527
rect 11663 46471 11719 46527
rect 11805 46471 11861 46527
rect 11947 46471 12003 46527
rect 12089 46471 12145 46527
rect 12231 46471 12287 46527
rect 12373 46471 12429 46527
rect 12515 46471 12571 46527
rect 12657 46471 12713 46527
rect 12799 46471 12855 46527
rect 12941 46471 12997 46527
rect 13083 46471 13139 46527
rect 13225 46471 13281 46527
rect 13367 46471 13423 46527
rect 13509 46471 13565 46527
rect 13651 46471 13707 46527
rect 13793 46471 13849 46527
rect 13935 46471 13991 46527
rect 14077 46471 14133 46527
rect 14219 46471 14275 46527
rect 14361 46471 14417 46527
rect 14503 46471 14559 46527
rect 14645 46471 14701 46527
rect 14787 46471 14843 46527
rect 161 46329 217 46385
rect 303 46329 359 46385
rect 445 46329 501 46385
rect 587 46329 643 46385
rect 729 46329 785 46385
rect 871 46329 927 46385
rect 1013 46329 1069 46385
rect 1155 46329 1211 46385
rect 1297 46329 1353 46385
rect 1439 46329 1495 46385
rect 1581 46329 1637 46385
rect 1723 46329 1779 46385
rect 1865 46329 1921 46385
rect 2007 46329 2063 46385
rect 2149 46329 2205 46385
rect 2291 46329 2347 46385
rect 2433 46329 2489 46385
rect 2575 46329 2631 46385
rect 2717 46329 2773 46385
rect 2859 46329 2915 46385
rect 3001 46329 3057 46385
rect 3143 46329 3199 46385
rect 3285 46329 3341 46385
rect 3427 46329 3483 46385
rect 3569 46329 3625 46385
rect 3711 46329 3767 46385
rect 3853 46329 3909 46385
rect 3995 46329 4051 46385
rect 4137 46329 4193 46385
rect 4279 46329 4335 46385
rect 4421 46329 4477 46385
rect 4563 46329 4619 46385
rect 4705 46329 4761 46385
rect 4847 46329 4903 46385
rect 4989 46329 5045 46385
rect 5131 46329 5187 46385
rect 5273 46329 5329 46385
rect 5415 46329 5471 46385
rect 5557 46329 5613 46385
rect 5699 46329 5755 46385
rect 5841 46329 5897 46385
rect 5983 46329 6039 46385
rect 6125 46329 6181 46385
rect 6267 46329 6323 46385
rect 6409 46329 6465 46385
rect 6551 46329 6607 46385
rect 6693 46329 6749 46385
rect 6835 46329 6891 46385
rect 6977 46329 7033 46385
rect 7119 46329 7175 46385
rect 7261 46329 7317 46385
rect 7403 46329 7459 46385
rect 7545 46329 7601 46385
rect 7687 46329 7743 46385
rect 7829 46329 7885 46385
rect 7971 46329 8027 46385
rect 8113 46329 8169 46385
rect 8255 46329 8311 46385
rect 8397 46329 8453 46385
rect 8539 46329 8595 46385
rect 8681 46329 8737 46385
rect 8823 46329 8879 46385
rect 8965 46329 9021 46385
rect 9107 46329 9163 46385
rect 9249 46329 9305 46385
rect 9391 46329 9447 46385
rect 9533 46329 9589 46385
rect 9675 46329 9731 46385
rect 9817 46329 9873 46385
rect 9959 46329 10015 46385
rect 10101 46329 10157 46385
rect 10243 46329 10299 46385
rect 10385 46329 10441 46385
rect 10527 46329 10583 46385
rect 10669 46329 10725 46385
rect 10811 46329 10867 46385
rect 10953 46329 11009 46385
rect 11095 46329 11151 46385
rect 11237 46329 11293 46385
rect 11379 46329 11435 46385
rect 11521 46329 11577 46385
rect 11663 46329 11719 46385
rect 11805 46329 11861 46385
rect 11947 46329 12003 46385
rect 12089 46329 12145 46385
rect 12231 46329 12287 46385
rect 12373 46329 12429 46385
rect 12515 46329 12571 46385
rect 12657 46329 12713 46385
rect 12799 46329 12855 46385
rect 12941 46329 12997 46385
rect 13083 46329 13139 46385
rect 13225 46329 13281 46385
rect 13367 46329 13423 46385
rect 13509 46329 13565 46385
rect 13651 46329 13707 46385
rect 13793 46329 13849 46385
rect 13935 46329 13991 46385
rect 14077 46329 14133 46385
rect 14219 46329 14275 46385
rect 14361 46329 14417 46385
rect 14503 46329 14559 46385
rect 14645 46329 14701 46385
rect 14787 46329 14843 46385
rect 161 46187 217 46243
rect 303 46187 359 46243
rect 445 46187 501 46243
rect 587 46187 643 46243
rect 729 46187 785 46243
rect 871 46187 927 46243
rect 1013 46187 1069 46243
rect 1155 46187 1211 46243
rect 1297 46187 1353 46243
rect 1439 46187 1495 46243
rect 1581 46187 1637 46243
rect 1723 46187 1779 46243
rect 1865 46187 1921 46243
rect 2007 46187 2063 46243
rect 2149 46187 2205 46243
rect 2291 46187 2347 46243
rect 2433 46187 2489 46243
rect 2575 46187 2631 46243
rect 2717 46187 2773 46243
rect 2859 46187 2915 46243
rect 3001 46187 3057 46243
rect 3143 46187 3199 46243
rect 3285 46187 3341 46243
rect 3427 46187 3483 46243
rect 3569 46187 3625 46243
rect 3711 46187 3767 46243
rect 3853 46187 3909 46243
rect 3995 46187 4051 46243
rect 4137 46187 4193 46243
rect 4279 46187 4335 46243
rect 4421 46187 4477 46243
rect 4563 46187 4619 46243
rect 4705 46187 4761 46243
rect 4847 46187 4903 46243
rect 4989 46187 5045 46243
rect 5131 46187 5187 46243
rect 5273 46187 5329 46243
rect 5415 46187 5471 46243
rect 5557 46187 5613 46243
rect 5699 46187 5755 46243
rect 5841 46187 5897 46243
rect 5983 46187 6039 46243
rect 6125 46187 6181 46243
rect 6267 46187 6323 46243
rect 6409 46187 6465 46243
rect 6551 46187 6607 46243
rect 6693 46187 6749 46243
rect 6835 46187 6891 46243
rect 6977 46187 7033 46243
rect 7119 46187 7175 46243
rect 7261 46187 7317 46243
rect 7403 46187 7459 46243
rect 7545 46187 7601 46243
rect 7687 46187 7743 46243
rect 7829 46187 7885 46243
rect 7971 46187 8027 46243
rect 8113 46187 8169 46243
rect 8255 46187 8311 46243
rect 8397 46187 8453 46243
rect 8539 46187 8595 46243
rect 8681 46187 8737 46243
rect 8823 46187 8879 46243
rect 8965 46187 9021 46243
rect 9107 46187 9163 46243
rect 9249 46187 9305 46243
rect 9391 46187 9447 46243
rect 9533 46187 9589 46243
rect 9675 46187 9731 46243
rect 9817 46187 9873 46243
rect 9959 46187 10015 46243
rect 10101 46187 10157 46243
rect 10243 46187 10299 46243
rect 10385 46187 10441 46243
rect 10527 46187 10583 46243
rect 10669 46187 10725 46243
rect 10811 46187 10867 46243
rect 10953 46187 11009 46243
rect 11095 46187 11151 46243
rect 11237 46187 11293 46243
rect 11379 46187 11435 46243
rect 11521 46187 11577 46243
rect 11663 46187 11719 46243
rect 11805 46187 11861 46243
rect 11947 46187 12003 46243
rect 12089 46187 12145 46243
rect 12231 46187 12287 46243
rect 12373 46187 12429 46243
rect 12515 46187 12571 46243
rect 12657 46187 12713 46243
rect 12799 46187 12855 46243
rect 12941 46187 12997 46243
rect 13083 46187 13139 46243
rect 13225 46187 13281 46243
rect 13367 46187 13423 46243
rect 13509 46187 13565 46243
rect 13651 46187 13707 46243
rect 13793 46187 13849 46243
rect 13935 46187 13991 46243
rect 14077 46187 14133 46243
rect 14219 46187 14275 46243
rect 14361 46187 14417 46243
rect 14503 46187 14559 46243
rect 14645 46187 14701 46243
rect 14787 46187 14843 46243
rect 161 46045 217 46101
rect 303 46045 359 46101
rect 445 46045 501 46101
rect 587 46045 643 46101
rect 729 46045 785 46101
rect 871 46045 927 46101
rect 1013 46045 1069 46101
rect 1155 46045 1211 46101
rect 1297 46045 1353 46101
rect 1439 46045 1495 46101
rect 1581 46045 1637 46101
rect 1723 46045 1779 46101
rect 1865 46045 1921 46101
rect 2007 46045 2063 46101
rect 2149 46045 2205 46101
rect 2291 46045 2347 46101
rect 2433 46045 2489 46101
rect 2575 46045 2631 46101
rect 2717 46045 2773 46101
rect 2859 46045 2915 46101
rect 3001 46045 3057 46101
rect 3143 46045 3199 46101
rect 3285 46045 3341 46101
rect 3427 46045 3483 46101
rect 3569 46045 3625 46101
rect 3711 46045 3767 46101
rect 3853 46045 3909 46101
rect 3995 46045 4051 46101
rect 4137 46045 4193 46101
rect 4279 46045 4335 46101
rect 4421 46045 4477 46101
rect 4563 46045 4619 46101
rect 4705 46045 4761 46101
rect 4847 46045 4903 46101
rect 4989 46045 5045 46101
rect 5131 46045 5187 46101
rect 5273 46045 5329 46101
rect 5415 46045 5471 46101
rect 5557 46045 5613 46101
rect 5699 46045 5755 46101
rect 5841 46045 5897 46101
rect 5983 46045 6039 46101
rect 6125 46045 6181 46101
rect 6267 46045 6323 46101
rect 6409 46045 6465 46101
rect 6551 46045 6607 46101
rect 6693 46045 6749 46101
rect 6835 46045 6891 46101
rect 6977 46045 7033 46101
rect 7119 46045 7175 46101
rect 7261 46045 7317 46101
rect 7403 46045 7459 46101
rect 7545 46045 7601 46101
rect 7687 46045 7743 46101
rect 7829 46045 7885 46101
rect 7971 46045 8027 46101
rect 8113 46045 8169 46101
rect 8255 46045 8311 46101
rect 8397 46045 8453 46101
rect 8539 46045 8595 46101
rect 8681 46045 8737 46101
rect 8823 46045 8879 46101
rect 8965 46045 9021 46101
rect 9107 46045 9163 46101
rect 9249 46045 9305 46101
rect 9391 46045 9447 46101
rect 9533 46045 9589 46101
rect 9675 46045 9731 46101
rect 9817 46045 9873 46101
rect 9959 46045 10015 46101
rect 10101 46045 10157 46101
rect 10243 46045 10299 46101
rect 10385 46045 10441 46101
rect 10527 46045 10583 46101
rect 10669 46045 10725 46101
rect 10811 46045 10867 46101
rect 10953 46045 11009 46101
rect 11095 46045 11151 46101
rect 11237 46045 11293 46101
rect 11379 46045 11435 46101
rect 11521 46045 11577 46101
rect 11663 46045 11719 46101
rect 11805 46045 11861 46101
rect 11947 46045 12003 46101
rect 12089 46045 12145 46101
rect 12231 46045 12287 46101
rect 12373 46045 12429 46101
rect 12515 46045 12571 46101
rect 12657 46045 12713 46101
rect 12799 46045 12855 46101
rect 12941 46045 12997 46101
rect 13083 46045 13139 46101
rect 13225 46045 13281 46101
rect 13367 46045 13423 46101
rect 13509 46045 13565 46101
rect 13651 46045 13707 46101
rect 13793 46045 13849 46101
rect 13935 46045 13991 46101
rect 14077 46045 14133 46101
rect 14219 46045 14275 46101
rect 14361 46045 14417 46101
rect 14503 46045 14559 46101
rect 14645 46045 14701 46101
rect 14787 46045 14843 46101
rect 161 45685 217 45741
rect 303 45685 359 45741
rect 445 45685 501 45741
rect 587 45685 643 45741
rect 729 45685 785 45741
rect 871 45685 927 45741
rect 1013 45685 1069 45741
rect 1155 45685 1211 45741
rect 1297 45685 1353 45741
rect 1439 45685 1495 45741
rect 1581 45685 1637 45741
rect 1723 45685 1779 45741
rect 1865 45685 1921 45741
rect 2007 45685 2063 45741
rect 2149 45685 2205 45741
rect 2291 45685 2347 45741
rect 2433 45685 2489 45741
rect 2575 45685 2631 45741
rect 2717 45685 2773 45741
rect 2859 45685 2915 45741
rect 3001 45685 3057 45741
rect 3143 45685 3199 45741
rect 3285 45685 3341 45741
rect 3427 45685 3483 45741
rect 3569 45685 3625 45741
rect 3711 45685 3767 45741
rect 3853 45685 3909 45741
rect 3995 45685 4051 45741
rect 4137 45685 4193 45741
rect 4279 45685 4335 45741
rect 4421 45685 4477 45741
rect 4563 45685 4619 45741
rect 4705 45685 4761 45741
rect 4847 45685 4903 45741
rect 4989 45685 5045 45741
rect 5131 45685 5187 45741
rect 5273 45685 5329 45741
rect 5415 45685 5471 45741
rect 5557 45685 5613 45741
rect 5699 45685 5755 45741
rect 5841 45685 5897 45741
rect 5983 45685 6039 45741
rect 6125 45685 6181 45741
rect 6267 45685 6323 45741
rect 6409 45685 6465 45741
rect 6551 45685 6607 45741
rect 6693 45685 6749 45741
rect 6835 45685 6891 45741
rect 6977 45685 7033 45741
rect 7119 45685 7175 45741
rect 7261 45685 7317 45741
rect 7403 45685 7459 45741
rect 7545 45685 7601 45741
rect 7687 45685 7743 45741
rect 7829 45685 7885 45741
rect 7971 45685 8027 45741
rect 8113 45685 8169 45741
rect 8255 45685 8311 45741
rect 8397 45685 8453 45741
rect 8539 45685 8595 45741
rect 8681 45685 8737 45741
rect 8823 45685 8879 45741
rect 8965 45685 9021 45741
rect 9107 45685 9163 45741
rect 9249 45685 9305 45741
rect 9391 45685 9447 45741
rect 9533 45685 9589 45741
rect 9675 45685 9731 45741
rect 9817 45685 9873 45741
rect 9959 45685 10015 45741
rect 10101 45685 10157 45741
rect 10243 45685 10299 45741
rect 10385 45685 10441 45741
rect 10527 45685 10583 45741
rect 10669 45685 10725 45741
rect 10811 45685 10867 45741
rect 10953 45685 11009 45741
rect 11095 45685 11151 45741
rect 11237 45685 11293 45741
rect 11379 45685 11435 45741
rect 11521 45685 11577 45741
rect 11663 45685 11719 45741
rect 11805 45685 11861 45741
rect 11947 45685 12003 45741
rect 12089 45685 12145 45741
rect 12231 45685 12287 45741
rect 12373 45685 12429 45741
rect 12515 45685 12571 45741
rect 12657 45685 12713 45741
rect 12799 45685 12855 45741
rect 12941 45685 12997 45741
rect 13083 45685 13139 45741
rect 13225 45685 13281 45741
rect 13367 45685 13423 45741
rect 13509 45685 13565 45741
rect 13651 45685 13707 45741
rect 13793 45685 13849 45741
rect 13935 45685 13991 45741
rect 14077 45685 14133 45741
rect 14219 45685 14275 45741
rect 14361 45685 14417 45741
rect 14503 45685 14559 45741
rect 14645 45685 14701 45741
rect 14787 45685 14843 45741
rect 161 45543 217 45599
rect 303 45543 359 45599
rect 445 45543 501 45599
rect 587 45543 643 45599
rect 729 45543 785 45599
rect 871 45543 927 45599
rect 1013 45543 1069 45599
rect 1155 45543 1211 45599
rect 1297 45543 1353 45599
rect 1439 45543 1495 45599
rect 1581 45543 1637 45599
rect 1723 45543 1779 45599
rect 1865 45543 1921 45599
rect 2007 45543 2063 45599
rect 2149 45543 2205 45599
rect 2291 45543 2347 45599
rect 2433 45543 2489 45599
rect 2575 45543 2631 45599
rect 2717 45543 2773 45599
rect 2859 45543 2915 45599
rect 3001 45543 3057 45599
rect 3143 45543 3199 45599
rect 3285 45543 3341 45599
rect 3427 45543 3483 45599
rect 3569 45543 3625 45599
rect 3711 45543 3767 45599
rect 3853 45543 3909 45599
rect 3995 45543 4051 45599
rect 4137 45543 4193 45599
rect 4279 45543 4335 45599
rect 4421 45543 4477 45599
rect 4563 45543 4619 45599
rect 4705 45543 4761 45599
rect 4847 45543 4903 45599
rect 4989 45543 5045 45599
rect 5131 45543 5187 45599
rect 5273 45543 5329 45599
rect 5415 45543 5471 45599
rect 5557 45543 5613 45599
rect 5699 45543 5755 45599
rect 5841 45543 5897 45599
rect 5983 45543 6039 45599
rect 6125 45543 6181 45599
rect 6267 45543 6323 45599
rect 6409 45543 6465 45599
rect 6551 45543 6607 45599
rect 6693 45543 6749 45599
rect 6835 45543 6891 45599
rect 6977 45543 7033 45599
rect 7119 45543 7175 45599
rect 7261 45543 7317 45599
rect 7403 45543 7459 45599
rect 7545 45543 7601 45599
rect 7687 45543 7743 45599
rect 7829 45543 7885 45599
rect 7971 45543 8027 45599
rect 8113 45543 8169 45599
rect 8255 45543 8311 45599
rect 8397 45543 8453 45599
rect 8539 45543 8595 45599
rect 8681 45543 8737 45599
rect 8823 45543 8879 45599
rect 8965 45543 9021 45599
rect 9107 45543 9163 45599
rect 9249 45543 9305 45599
rect 9391 45543 9447 45599
rect 9533 45543 9589 45599
rect 9675 45543 9731 45599
rect 9817 45543 9873 45599
rect 9959 45543 10015 45599
rect 10101 45543 10157 45599
rect 10243 45543 10299 45599
rect 10385 45543 10441 45599
rect 10527 45543 10583 45599
rect 10669 45543 10725 45599
rect 10811 45543 10867 45599
rect 10953 45543 11009 45599
rect 11095 45543 11151 45599
rect 11237 45543 11293 45599
rect 11379 45543 11435 45599
rect 11521 45543 11577 45599
rect 11663 45543 11719 45599
rect 11805 45543 11861 45599
rect 11947 45543 12003 45599
rect 12089 45543 12145 45599
rect 12231 45543 12287 45599
rect 12373 45543 12429 45599
rect 12515 45543 12571 45599
rect 12657 45543 12713 45599
rect 12799 45543 12855 45599
rect 12941 45543 12997 45599
rect 13083 45543 13139 45599
rect 13225 45543 13281 45599
rect 13367 45543 13423 45599
rect 13509 45543 13565 45599
rect 13651 45543 13707 45599
rect 13793 45543 13849 45599
rect 13935 45543 13991 45599
rect 14077 45543 14133 45599
rect 14219 45543 14275 45599
rect 14361 45543 14417 45599
rect 14503 45543 14559 45599
rect 14645 45543 14701 45599
rect 14787 45543 14843 45599
rect 161 45401 217 45457
rect 303 45401 359 45457
rect 445 45401 501 45457
rect 587 45401 643 45457
rect 729 45401 785 45457
rect 871 45401 927 45457
rect 1013 45401 1069 45457
rect 1155 45401 1211 45457
rect 1297 45401 1353 45457
rect 1439 45401 1495 45457
rect 1581 45401 1637 45457
rect 1723 45401 1779 45457
rect 1865 45401 1921 45457
rect 2007 45401 2063 45457
rect 2149 45401 2205 45457
rect 2291 45401 2347 45457
rect 2433 45401 2489 45457
rect 2575 45401 2631 45457
rect 2717 45401 2773 45457
rect 2859 45401 2915 45457
rect 3001 45401 3057 45457
rect 3143 45401 3199 45457
rect 3285 45401 3341 45457
rect 3427 45401 3483 45457
rect 3569 45401 3625 45457
rect 3711 45401 3767 45457
rect 3853 45401 3909 45457
rect 3995 45401 4051 45457
rect 4137 45401 4193 45457
rect 4279 45401 4335 45457
rect 4421 45401 4477 45457
rect 4563 45401 4619 45457
rect 4705 45401 4761 45457
rect 4847 45401 4903 45457
rect 4989 45401 5045 45457
rect 5131 45401 5187 45457
rect 5273 45401 5329 45457
rect 5415 45401 5471 45457
rect 5557 45401 5613 45457
rect 5699 45401 5755 45457
rect 5841 45401 5897 45457
rect 5983 45401 6039 45457
rect 6125 45401 6181 45457
rect 6267 45401 6323 45457
rect 6409 45401 6465 45457
rect 6551 45401 6607 45457
rect 6693 45401 6749 45457
rect 6835 45401 6891 45457
rect 6977 45401 7033 45457
rect 7119 45401 7175 45457
rect 7261 45401 7317 45457
rect 7403 45401 7459 45457
rect 7545 45401 7601 45457
rect 7687 45401 7743 45457
rect 7829 45401 7885 45457
rect 7971 45401 8027 45457
rect 8113 45401 8169 45457
rect 8255 45401 8311 45457
rect 8397 45401 8453 45457
rect 8539 45401 8595 45457
rect 8681 45401 8737 45457
rect 8823 45401 8879 45457
rect 8965 45401 9021 45457
rect 9107 45401 9163 45457
rect 9249 45401 9305 45457
rect 9391 45401 9447 45457
rect 9533 45401 9589 45457
rect 9675 45401 9731 45457
rect 9817 45401 9873 45457
rect 9959 45401 10015 45457
rect 10101 45401 10157 45457
rect 10243 45401 10299 45457
rect 10385 45401 10441 45457
rect 10527 45401 10583 45457
rect 10669 45401 10725 45457
rect 10811 45401 10867 45457
rect 10953 45401 11009 45457
rect 11095 45401 11151 45457
rect 11237 45401 11293 45457
rect 11379 45401 11435 45457
rect 11521 45401 11577 45457
rect 11663 45401 11719 45457
rect 11805 45401 11861 45457
rect 11947 45401 12003 45457
rect 12089 45401 12145 45457
rect 12231 45401 12287 45457
rect 12373 45401 12429 45457
rect 12515 45401 12571 45457
rect 12657 45401 12713 45457
rect 12799 45401 12855 45457
rect 12941 45401 12997 45457
rect 13083 45401 13139 45457
rect 13225 45401 13281 45457
rect 13367 45401 13423 45457
rect 13509 45401 13565 45457
rect 13651 45401 13707 45457
rect 13793 45401 13849 45457
rect 13935 45401 13991 45457
rect 14077 45401 14133 45457
rect 14219 45401 14275 45457
rect 14361 45401 14417 45457
rect 14503 45401 14559 45457
rect 14645 45401 14701 45457
rect 14787 45401 14843 45457
rect 161 45259 217 45315
rect 303 45259 359 45315
rect 445 45259 501 45315
rect 587 45259 643 45315
rect 729 45259 785 45315
rect 871 45259 927 45315
rect 1013 45259 1069 45315
rect 1155 45259 1211 45315
rect 1297 45259 1353 45315
rect 1439 45259 1495 45315
rect 1581 45259 1637 45315
rect 1723 45259 1779 45315
rect 1865 45259 1921 45315
rect 2007 45259 2063 45315
rect 2149 45259 2205 45315
rect 2291 45259 2347 45315
rect 2433 45259 2489 45315
rect 2575 45259 2631 45315
rect 2717 45259 2773 45315
rect 2859 45259 2915 45315
rect 3001 45259 3057 45315
rect 3143 45259 3199 45315
rect 3285 45259 3341 45315
rect 3427 45259 3483 45315
rect 3569 45259 3625 45315
rect 3711 45259 3767 45315
rect 3853 45259 3909 45315
rect 3995 45259 4051 45315
rect 4137 45259 4193 45315
rect 4279 45259 4335 45315
rect 4421 45259 4477 45315
rect 4563 45259 4619 45315
rect 4705 45259 4761 45315
rect 4847 45259 4903 45315
rect 4989 45259 5045 45315
rect 5131 45259 5187 45315
rect 5273 45259 5329 45315
rect 5415 45259 5471 45315
rect 5557 45259 5613 45315
rect 5699 45259 5755 45315
rect 5841 45259 5897 45315
rect 5983 45259 6039 45315
rect 6125 45259 6181 45315
rect 6267 45259 6323 45315
rect 6409 45259 6465 45315
rect 6551 45259 6607 45315
rect 6693 45259 6749 45315
rect 6835 45259 6891 45315
rect 6977 45259 7033 45315
rect 7119 45259 7175 45315
rect 7261 45259 7317 45315
rect 7403 45259 7459 45315
rect 7545 45259 7601 45315
rect 7687 45259 7743 45315
rect 7829 45259 7885 45315
rect 7971 45259 8027 45315
rect 8113 45259 8169 45315
rect 8255 45259 8311 45315
rect 8397 45259 8453 45315
rect 8539 45259 8595 45315
rect 8681 45259 8737 45315
rect 8823 45259 8879 45315
rect 8965 45259 9021 45315
rect 9107 45259 9163 45315
rect 9249 45259 9305 45315
rect 9391 45259 9447 45315
rect 9533 45259 9589 45315
rect 9675 45259 9731 45315
rect 9817 45259 9873 45315
rect 9959 45259 10015 45315
rect 10101 45259 10157 45315
rect 10243 45259 10299 45315
rect 10385 45259 10441 45315
rect 10527 45259 10583 45315
rect 10669 45259 10725 45315
rect 10811 45259 10867 45315
rect 10953 45259 11009 45315
rect 11095 45259 11151 45315
rect 11237 45259 11293 45315
rect 11379 45259 11435 45315
rect 11521 45259 11577 45315
rect 11663 45259 11719 45315
rect 11805 45259 11861 45315
rect 11947 45259 12003 45315
rect 12089 45259 12145 45315
rect 12231 45259 12287 45315
rect 12373 45259 12429 45315
rect 12515 45259 12571 45315
rect 12657 45259 12713 45315
rect 12799 45259 12855 45315
rect 12941 45259 12997 45315
rect 13083 45259 13139 45315
rect 13225 45259 13281 45315
rect 13367 45259 13423 45315
rect 13509 45259 13565 45315
rect 13651 45259 13707 45315
rect 13793 45259 13849 45315
rect 13935 45259 13991 45315
rect 14077 45259 14133 45315
rect 14219 45259 14275 45315
rect 14361 45259 14417 45315
rect 14503 45259 14559 45315
rect 14645 45259 14701 45315
rect 14787 45259 14843 45315
rect 161 45117 217 45173
rect 303 45117 359 45173
rect 445 45117 501 45173
rect 587 45117 643 45173
rect 729 45117 785 45173
rect 871 45117 927 45173
rect 1013 45117 1069 45173
rect 1155 45117 1211 45173
rect 1297 45117 1353 45173
rect 1439 45117 1495 45173
rect 1581 45117 1637 45173
rect 1723 45117 1779 45173
rect 1865 45117 1921 45173
rect 2007 45117 2063 45173
rect 2149 45117 2205 45173
rect 2291 45117 2347 45173
rect 2433 45117 2489 45173
rect 2575 45117 2631 45173
rect 2717 45117 2773 45173
rect 2859 45117 2915 45173
rect 3001 45117 3057 45173
rect 3143 45117 3199 45173
rect 3285 45117 3341 45173
rect 3427 45117 3483 45173
rect 3569 45117 3625 45173
rect 3711 45117 3767 45173
rect 3853 45117 3909 45173
rect 3995 45117 4051 45173
rect 4137 45117 4193 45173
rect 4279 45117 4335 45173
rect 4421 45117 4477 45173
rect 4563 45117 4619 45173
rect 4705 45117 4761 45173
rect 4847 45117 4903 45173
rect 4989 45117 5045 45173
rect 5131 45117 5187 45173
rect 5273 45117 5329 45173
rect 5415 45117 5471 45173
rect 5557 45117 5613 45173
rect 5699 45117 5755 45173
rect 5841 45117 5897 45173
rect 5983 45117 6039 45173
rect 6125 45117 6181 45173
rect 6267 45117 6323 45173
rect 6409 45117 6465 45173
rect 6551 45117 6607 45173
rect 6693 45117 6749 45173
rect 6835 45117 6891 45173
rect 6977 45117 7033 45173
rect 7119 45117 7175 45173
rect 7261 45117 7317 45173
rect 7403 45117 7459 45173
rect 7545 45117 7601 45173
rect 7687 45117 7743 45173
rect 7829 45117 7885 45173
rect 7971 45117 8027 45173
rect 8113 45117 8169 45173
rect 8255 45117 8311 45173
rect 8397 45117 8453 45173
rect 8539 45117 8595 45173
rect 8681 45117 8737 45173
rect 8823 45117 8879 45173
rect 8965 45117 9021 45173
rect 9107 45117 9163 45173
rect 9249 45117 9305 45173
rect 9391 45117 9447 45173
rect 9533 45117 9589 45173
rect 9675 45117 9731 45173
rect 9817 45117 9873 45173
rect 9959 45117 10015 45173
rect 10101 45117 10157 45173
rect 10243 45117 10299 45173
rect 10385 45117 10441 45173
rect 10527 45117 10583 45173
rect 10669 45117 10725 45173
rect 10811 45117 10867 45173
rect 10953 45117 11009 45173
rect 11095 45117 11151 45173
rect 11237 45117 11293 45173
rect 11379 45117 11435 45173
rect 11521 45117 11577 45173
rect 11663 45117 11719 45173
rect 11805 45117 11861 45173
rect 11947 45117 12003 45173
rect 12089 45117 12145 45173
rect 12231 45117 12287 45173
rect 12373 45117 12429 45173
rect 12515 45117 12571 45173
rect 12657 45117 12713 45173
rect 12799 45117 12855 45173
rect 12941 45117 12997 45173
rect 13083 45117 13139 45173
rect 13225 45117 13281 45173
rect 13367 45117 13423 45173
rect 13509 45117 13565 45173
rect 13651 45117 13707 45173
rect 13793 45117 13849 45173
rect 13935 45117 13991 45173
rect 14077 45117 14133 45173
rect 14219 45117 14275 45173
rect 14361 45117 14417 45173
rect 14503 45117 14559 45173
rect 14645 45117 14701 45173
rect 14787 45117 14843 45173
rect 161 44975 217 45031
rect 303 44975 359 45031
rect 445 44975 501 45031
rect 587 44975 643 45031
rect 729 44975 785 45031
rect 871 44975 927 45031
rect 1013 44975 1069 45031
rect 1155 44975 1211 45031
rect 1297 44975 1353 45031
rect 1439 44975 1495 45031
rect 1581 44975 1637 45031
rect 1723 44975 1779 45031
rect 1865 44975 1921 45031
rect 2007 44975 2063 45031
rect 2149 44975 2205 45031
rect 2291 44975 2347 45031
rect 2433 44975 2489 45031
rect 2575 44975 2631 45031
rect 2717 44975 2773 45031
rect 2859 44975 2915 45031
rect 3001 44975 3057 45031
rect 3143 44975 3199 45031
rect 3285 44975 3341 45031
rect 3427 44975 3483 45031
rect 3569 44975 3625 45031
rect 3711 44975 3767 45031
rect 3853 44975 3909 45031
rect 3995 44975 4051 45031
rect 4137 44975 4193 45031
rect 4279 44975 4335 45031
rect 4421 44975 4477 45031
rect 4563 44975 4619 45031
rect 4705 44975 4761 45031
rect 4847 44975 4903 45031
rect 4989 44975 5045 45031
rect 5131 44975 5187 45031
rect 5273 44975 5329 45031
rect 5415 44975 5471 45031
rect 5557 44975 5613 45031
rect 5699 44975 5755 45031
rect 5841 44975 5897 45031
rect 5983 44975 6039 45031
rect 6125 44975 6181 45031
rect 6267 44975 6323 45031
rect 6409 44975 6465 45031
rect 6551 44975 6607 45031
rect 6693 44975 6749 45031
rect 6835 44975 6891 45031
rect 6977 44975 7033 45031
rect 7119 44975 7175 45031
rect 7261 44975 7317 45031
rect 7403 44975 7459 45031
rect 7545 44975 7601 45031
rect 7687 44975 7743 45031
rect 7829 44975 7885 45031
rect 7971 44975 8027 45031
rect 8113 44975 8169 45031
rect 8255 44975 8311 45031
rect 8397 44975 8453 45031
rect 8539 44975 8595 45031
rect 8681 44975 8737 45031
rect 8823 44975 8879 45031
rect 8965 44975 9021 45031
rect 9107 44975 9163 45031
rect 9249 44975 9305 45031
rect 9391 44975 9447 45031
rect 9533 44975 9589 45031
rect 9675 44975 9731 45031
rect 9817 44975 9873 45031
rect 9959 44975 10015 45031
rect 10101 44975 10157 45031
rect 10243 44975 10299 45031
rect 10385 44975 10441 45031
rect 10527 44975 10583 45031
rect 10669 44975 10725 45031
rect 10811 44975 10867 45031
rect 10953 44975 11009 45031
rect 11095 44975 11151 45031
rect 11237 44975 11293 45031
rect 11379 44975 11435 45031
rect 11521 44975 11577 45031
rect 11663 44975 11719 45031
rect 11805 44975 11861 45031
rect 11947 44975 12003 45031
rect 12089 44975 12145 45031
rect 12231 44975 12287 45031
rect 12373 44975 12429 45031
rect 12515 44975 12571 45031
rect 12657 44975 12713 45031
rect 12799 44975 12855 45031
rect 12941 44975 12997 45031
rect 13083 44975 13139 45031
rect 13225 44975 13281 45031
rect 13367 44975 13423 45031
rect 13509 44975 13565 45031
rect 13651 44975 13707 45031
rect 13793 44975 13849 45031
rect 13935 44975 13991 45031
rect 14077 44975 14133 45031
rect 14219 44975 14275 45031
rect 14361 44975 14417 45031
rect 14503 44975 14559 45031
rect 14645 44975 14701 45031
rect 14787 44975 14843 45031
rect 161 44833 217 44889
rect 303 44833 359 44889
rect 445 44833 501 44889
rect 587 44833 643 44889
rect 729 44833 785 44889
rect 871 44833 927 44889
rect 1013 44833 1069 44889
rect 1155 44833 1211 44889
rect 1297 44833 1353 44889
rect 1439 44833 1495 44889
rect 1581 44833 1637 44889
rect 1723 44833 1779 44889
rect 1865 44833 1921 44889
rect 2007 44833 2063 44889
rect 2149 44833 2205 44889
rect 2291 44833 2347 44889
rect 2433 44833 2489 44889
rect 2575 44833 2631 44889
rect 2717 44833 2773 44889
rect 2859 44833 2915 44889
rect 3001 44833 3057 44889
rect 3143 44833 3199 44889
rect 3285 44833 3341 44889
rect 3427 44833 3483 44889
rect 3569 44833 3625 44889
rect 3711 44833 3767 44889
rect 3853 44833 3909 44889
rect 3995 44833 4051 44889
rect 4137 44833 4193 44889
rect 4279 44833 4335 44889
rect 4421 44833 4477 44889
rect 4563 44833 4619 44889
rect 4705 44833 4761 44889
rect 4847 44833 4903 44889
rect 4989 44833 5045 44889
rect 5131 44833 5187 44889
rect 5273 44833 5329 44889
rect 5415 44833 5471 44889
rect 5557 44833 5613 44889
rect 5699 44833 5755 44889
rect 5841 44833 5897 44889
rect 5983 44833 6039 44889
rect 6125 44833 6181 44889
rect 6267 44833 6323 44889
rect 6409 44833 6465 44889
rect 6551 44833 6607 44889
rect 6693 44833 6749 44889
rect 6835 44833 6891 44889
rect 6977 44833 7033 44889
rect 7119 44833 7175 44889
rect 7261 44833 7317 44889
rect 7403 44833 7459 44889
rect 7545 44833 7601 44889
rect 7687 44833 7743 44889
rect 7829 44833 7885 44889
rect 7971 44833 8027 44889
rect 8113 44833 8169 44889
rect 8255 44833 8311 44889
rect 8397 44833 8453 44889
rect 8539 44833 8595 44889
rect 8681 44833 8737 44889
rect 8823 44833 8879 44889
rect 8965 44833 9021 44889
rect 9107 44833 9163 44889
rect 9249 44833 9305 44889
rect 9391 44833 9447 44889
rect 9533 44833 9589 44889
rect 9675 44833 9731 44889
rect 9817 44833 9873 44889
rect 9959 44833 10015 44889
rect 10101 44833 10157 44889
rect 10243 44833 10299 44889
rect 10385 44833 10441 44889
rect 10527 44833 10583 44889
rect 10669 44833 10725 44889
rect 10811 44833 10867 44889
rect 10953 44833 11009 44889
rect 11095 44833 11151 44889
rect 11237 44833 11293 44889
rect 11379 44833 11435 44889
rect 11521 44833 11577 44889
rect 11663 44833 11719 44889
rect 11805 44833 11861 44889
rect 11947 44833 12003 44889
rect 12089 44833 12145 44889
rect 12231 44833 12287 44889
rect 12373 44833 12429 44889
rect 12515 44833 12571 44889
rect 12657 44833 12713 44889
rect 12799 44833 12855 44889
rect 12941 44833 12997 44889
rect 13083 44833 13139 44889
rect 13225 44833 13281 44889
rect 13367 44833 13423 44889
rect 13509 44833 13565 44889
rect 13651 44833 13707 44889
rect 13793 44833 13849 44889
rect 13935 44833 13991 44889
rect 14077 44833 14133 44889
rect 14219 44833 14275 44889
rect 14361 44833 14417 44889
rect 14503 44833 14559 44889
rect 14645 44833 14701 44889
rect 14787 44833 14843 44889
rect 161 44691 217 44747
rect 303 44691 359 44747
rect 445 44691 501 44747
rect 587 44691 643 44747
rect 729 44691 785 44747
rect 871 44691 927 44747
rect 1013 44691 1069 44747
rect 1155 44691 1211 44747
rect 1297 44691 1353 44747
rect 1439 44691 1495 44747
rect 1581 44691 1637 44747
rect 1723 44691 1779 44747
rect 1865 44691 1921 44747
rect 2007 44691 2063 44747
rect 2149 44691 2205 44747
rect 2291 44691 2347 44747
rect 2433 44691 2489 44747
rect 2575 44691 2631 44747
rect 2717 44691 2773 44747
rect 2859 44691 2915 44747
rect 3001 44691 3057 44747
rect 3143 44691 3199 44747
rect 3285 44691 3341 44747
rect 3427 44691 3483 44747
rect 3569 44691 3625 44747
rect 3711 44691 3767 44747
rect 3853 44691 3909 44747
rect 3995 44691 4051 44747
rect 4137 44691 4193 44747
rect 4279 44691 4335 44747
rect 4421 44691 4477 44747
rect 4563 44691 4619 44747
rect 4705 44691 4761 44747
rect 4847 44691 4903 44747
rect 4989 44691 5045 44747
rect 5131 44691 5187 44747
rect 5273 44691 5329 44747
rect 5415 44691 5471 44747
rect 5557 44691 5613 44747
rect 5699 44691 5755 44747
rect 5841 44691 5897 44747
rect 5983 44691 6039 44747
rect 6125 44691 6181 44747
rect 6267 44691 6323 44747
rect 6409 44691 6465 44747
rect 6551 44691 6607 44747
rect 6693 44691 6749 44747
rect 6835 44691 6891 44747
rect 6977 44691 7033 44747
rect 7119 44691 7175 44747
rect 7261 44691 7317 44747
rect 7403 44691 7459 44747
rect 7545 44691 7601 44747
rect 7687 44691 7743 44747
rect 7829 44691 7885 44747
rect 7971 44691 8027 44747
rect 8113 44691 8169 44747
rect 8255 44691 8311 44747
rect 8397 44691 8453 44747
rect 8539 44691 8595 44747
rect 8681 44691 8737 44747
rect 8823 44691 8879 44747
rect 8965 44691 9021 44747
rect 9107 44691 9163 44747
rect 9249 44691 9305 44747
rect 9391 44691 9447 44747
rect 9533 44691 9589 44747
rect 9675 44691 9731 44747
rect 9817 44691 9873 44747
rect 9959 44691 10015 44747
rect 10101 44691 10157 44747
rect 10243 44691 10299 44747
rect 10385 44691 10441 44747
rect 10527 44691 10583 44747
rect 10669 44691 10725 44747
rect 10811 44691 10867 44747
rect 10953 44691 11009 44747
rect 11095 44691 11151 44747
rect 11237 44691 11293 44747
rect 11379 44691 11435 44747
rect 11521 44691 11577 44747
rect 11663 44691 11719 44747
rect 11805 44691 11861 44747
rect 11947 44691 12003 44747
rect 12089 44691 12145 44747
rect 12231 44691 12287 44747
rect 12373 44691 12429 44747
rect 12515 44691 12571 44747
rect 12657 44691 12713 44747
rect 12799 44691 12855 44747
rect 12941 44691 12997 44747
rect 13083 44691 13139 44747
rect 13225 44691 13281 44747
rect 13367 44691 13423 44747
rect 13509 44691 13565 44747
rect 13651 44691 13707 44747
rect 13793 44691 13849 44747
rect 13935 44691 13991 44747
rect 14077 44691 14133 44747
rect 14219 44691 14275 44747
rect 14361 44691 14417 44747
rect 14503 44691 14559 44747
rect 14645 44691 14701 44747
rect 14787 44691 14843 44747
rect 161 44549 217 44605
rect 303 44549 359 44605
rect 445 44549 501 44605
rect 587 44549 643 44605
rect 729 44549 785 44605
rect 871 44549 927 44605
rect 1013 44549 1069 44605
rect 1155 44549 1211 44605
rect 1297 44549 1353 44605
rect 1439 44549 1495 44605
rect 1581 44549 1637 44605
rect 1723 44549 1779 44605
rect 1865 44549 1921 44605
rect 2007 44549 2063 44605
rect 2149 44549 2205 44605
rect 2291 44549 2347 44605
rect 2433 44549 2489 44605
rect 2575 44549 2631 44605
rect 2717 44549 2773 44605
rect 2859 44549 2915 44605
rect 3001 44549 3057 44605
rect 3143 44549 3199 44605
rect 3285 44549 3341 44605
rect 3427 44549 3483 44605
rect 3569 44549 3625 44605
rect 3711 44549 3767 44605
rect 3853 44549 3909 44605
rect 3995 44549 4051 44605
rect 4137 44549 4193 44605
rect 4279 44549 4335 44605
rect 4421 44549 4477 44605
rect 4563 44549 4619 44605
rect 4705 44549 4761 44605
rect 4847 44549 4903 44605
rect 4989 44549 5045 44605
rect 5131 44549 5187 44605
rect 5273 44549 5329 44605
rect 5415 44549 5471 44605
rect 5557 44549 5613 44605
rect 5699 44549 5755 44605
rect 5841 44549 5897 44605
rect 5983 44549 6039 44605
rect 6125 44549 6181 44605
rect 6267 44549 6323 44605
rect 6409 44549 6465 44605
rect 6551 44549 6607 44605
rect 6693 44549 6749 44605
rect 6835 44549 6891 44605
rect 6977 44549 7033 44605
rect 7119 44549 7175 44605
rect 7261 44549 7317 44605
rect 7403 44549 7459 44605
rect 7545 44549 7601 44605
rect 7687 44549 7743 44605
rect 7829 44549 7885 44605
rect 7971 44549 8027 44605
rect 8113 44549 8169 44605
rect 8255 44549 8311 44605
rect 8397 44549 8453 44605
rect 8539 44549 8595 44605
rect 8681 44549 8737 44605
rect 8823 44549 8879 44605
rect 8965 44549 9021 44605
rect 9107 44549 9163 44605
rect 9249 44549 9305 44605
rect 9391 44549 9447 44605
rect 9533 44549 9589 44605
rect 9675 44549 9731 44605
rect 9817 44549 9873 44605
rect 9959 44549 10015 44605
rect 10101 44549 10157 44605
rect 10243 44549 10299 44605
rect 10385 44549 10441 44605
rect 10527 44549 10583 44605
rect 10669 44549 10725 44605
rect 10811 44549 10867 44605
rect 10953 44549 11009 44605
rect 11095 44549 11151 44605
rect 11237 44549 11293 44605
rect 11379 44549 11435 44605
rect 11521 44549 11577 44605
rect 11663 44549 11719 44605
rect 11805 44549 11861 44605
rect 11947 44549 12003 44605
rect 12089 44549 12145 44605
rect 12231 44549 12287 44605
rect 12373 44549 12429 44605
rect 12515 44549 12571 44605
rect 12657 44549 12713 44605
rect 12799 44549 12855 44605
rect 12941 44549 12997 44605
rect 13083 44549 13139 44605
rect 13225 44549 13281 44605
rect 13367 44549 13423 44605
rect 13509 44549 13565 44605
rect 13651 44549 13707 44605
rect 13793 44549 13849 44605
rect 13935 44549 13991 44605
rect 14077 44549 14133 44605
rect 14219 44549 14275 44605
rect 14361 44549 14417 44605
rect 14503 44549 14559 44605
rect 14645 44549 14701 44605
rect 14787 44549 14843 44605
rect 161 44407 217 44463
rect 303 44407 359 44463
rect 445 44407 501 44463
rect 587 44407 643 44463
rect 729 44407 785 44463
rect 871 44407 927 44463
rect 1013 44407 1069 44463
rect 1155 44407 1211 44463
rect 1297 44407 1353 44463
rect 1439 44407 1495 44463
rect 1581 44407 1637 44463
rect 1723 44407 1779 44463
rect 1865 44407 1921 44463
rect 2007 44407 2063 44463
rect 2149 44407 2205 44463
rect 2291 44407 2347 44463
rect 2433 44407 2489 44463
rect 2575 44407 2631 44463
rect 2717 44407 2773 44463
rect 2859 44407 2915 44463
rect 3001 44407 3057 44463
rect 3143 44407 3199 44463
rect 3285 44407 3341 44463
rect 3427 44407 3483 44463
rect 3569 44407 3625 44463
rect 3711 44407 3767 44463
rect 3853 44407 3909 44463
rect 3995 44407 4051 44463
rect 4137 44407 4193 44463
rect 4279 44407 4335 44463
rect 4421 44407 4477 44463
rect 4563 44407 4619 44463
rect 4705 44407 4761 44463
rect 4847 44407 4903 44463
rect 4989 44407 5045 44463
rect 5131 44407 5187 44463
rect 5273 44407 5329 44463
rect 5415 44407 5471 44463
rect 5557 44407 5613 44463
rect 5699 44407 5755 44463
rect 5841 44407 5897 44463
rect 5983 44407 6039 44463
rect 6125 44407 6181 44463
rect 6267 44407 6323 44463
rect 6409 44407 6465 44463
rect 6551 44407 6607 44463
rect 6693 44407 6749 44463
rect 6835 44407 6891 44463
rect 6977 44407 7033 44463
rect 7119 44407 7175 44463
rect 7261 44407 7317 44463
rect 7403 44407 7459 44463
rect 7545 44407 7601 44463
rect 7687 44407 7743 44463
rect 7829 44407 7885 44463
rect 7971 44407 8027 44463
rect 8113 44407 8169 44463
rect 8255 44407 8311 44463
rect 8397 44407 8453 44463
rect 8539 44407 8595 44463
rect 8681 44407 8737 44463
rect 8823 44407 8879 44463
rect 8965 44407 9021 44463
rect 9107 44407 9163 44463
rect 9249 44407 9305 44463
rect 9391 44407 9447 44463
rect 9533 44407 9589 44463
rect 9675 44407 9731 44463
rect 9817 44407 9873 44463
rect 9959 44407 10015 44463
rect 10101 44407 10157 44463
rect 10243 44407 10299 44463
rect 10385 44407 10441 44463
rect 10527 44407 10583 44463
rect 10669 44407 10725 44463
rect 10811 44407 10867 44463
rect 10953 44407 11009 44463
rect 11095 44407 11151 44463
rect 11237 44407 11293 44463
rect 11379 44407 11435 44463
rect 11521 44407 11577 44463
rect 11663 44407 11719 44463
rect 11805 44407 11861 44463
rect 11947 44407 12003 44463
rect 12089 44407 12145 44463
rect 12231 44407 12287 44463
rect 12373 44407 12429 44463
rect 12515 44407 12571 44463
rect 12657 44407 12713 44463
rect 12799 44407 12855 44463
rect 12941 44407 12997 44463
rect 13083 44407 13139 44463
rect 13225 44407 13281 44463
rect 13367 44407 13423 44463
rect 13509 44407 13565 44463
rect 13651 44407 13707 44463
rect 13793 44407 13849 44463
rect 13935 44407 13991 44463
rect 14077 44407 14133 44463
rect 14219 44407 14275 44463
rect 14361 44407 14417 44463
rect 14503 44407 14559 44463
rect 14645 44407 14701 44463
rect 14787 44407 14843 44463
rect 161 44265 217 44321
rect 303 44265 359 44321
rect 445 44265 501 44321
rect 587 44265 643 44321
rect 729 44265 785 44321
rect 871 44265 927 44321
rect 1013 44265 1069 44321
rect 1155 44265 1211 44321
rect 1297 44265 1353 44321
rect 1439 44265 1495 44321
rect 1581 44265 1637 44321
rect 1723 44265 1779 44321
rect 1865 44265 1921 44321
rect 2007 44265 2063 44321
rect 2149 44265 2205 44321
rect 2291 44265 2347 44321
rect 2433 44265 2489 44321
rect 2575 44265 2631 44321
rect 2717 44265 2773 44321
rect 2859 44265 2915 44321
rect 3001 44265 3057 44321
rect 3143 44265 3199 44321
rect 3285 44265 3341 44321
rect 3427 44265 3483 44321
rect 3569 44265 3625 44321
rect 3711 44265 3767 44321
rect 3853 44265 3909 44321
rect 3995 44265 4051 44321
rect 4137 44265 4193 44321
rect 4279 44265 4335 44321
rect 4421 44265 4477 44321
rect 4563 44265 4619 44321
rect 4705 44265 4761 44321
rect 4847 44265 4903 44321
rect 4989 44265 5045 44321
rect 5131 44265 5187 44321
rect 5273 44265 5329 44321
rect 5415 44265 5471 44321
rect 5557 44265 5613 44321
rect 5699 44265 5755 44321
rect 5841 44265 5897 44321
rect 5983 44265 6039 44321
rect 6125 44265 6181 44321
rect 6267 44265 6323 44321
rect 6409 44265 6465 44321
rect 6551 44265 6607 44321
rect 6693 44265 6749 44321
rect 6835 44265 6891 44321
rect 6977 44265 7033 44321
rect 7119 44265 7175 44321
rect 7261 44265 7317 44321
rect 7403 44265 7459 44321
rect 7545 44265 7601 44321
rect 7687 44265 7743 44321
rect 7829 44265 7885 44321
rect 7971 44265 8027 44321
rect 8113 44265 8169 44321
rect 8255 44265 8311 44321
rect 8397 44265 8453 44321
rect 8539 44265 8595 44321
rect 8681 44265 8737 44321
rect 8823 44265 8879 44321
rect 8965 44265 9021 44321
rect 9107 44265 9163 44321
rect 9249 44265 9305 44321
rect 9391 44265 9447 44321
rect 9533 44265 9589 44321
rect 9675 44265 9731 44321
rect 9817 44265 9873 44321
rect 9959 44265 10015 44321
rect 10101 44265 10157 44321
rect 10243 44265 10299 44321
rect 10385 44265 10441 44321
rect 10527 44265 10583 44321
rect 10669 44265 10725 44321
rect 10811 44265 10867 44321
rect 10953 44265 11009 44321
rect 11095 44265 11151 44321
rect 11237 44265 11293 44321
rect 11379 44265 11435 44321
rect 11521 44265 11577 44321
rect 11663 44265 11719 44321
rect 11805 44265 11861 44321
rect 11947 44265 12003 44321
rect 12089 44265 12145 44321
rect 12231 44265 12287 44321
rect 12373 44265 12429 44321
rect 12515 44265 12571 44321
rect 12657 44265 12713 44321
rect 12799 44265 12855 44321
rect 12941 44265 12997 44321
rect 13083 44265 13139 44321
rect 13225 44265 13281 44321
rect 13367 44265 13423 44321
rect 13509 44265 13565 44321
rect 13651 44265 13707 44321
rect 13793 44265 13849 44321
rect 13935 44265 13991 44321
rect 14077 44265 14133 44321
rect 14219 44265 14275 44321
rect 14361 44265 14417 44321
rect 14503 44265 14559 44321
rect 14645 44265 14701 44321
rect 14787 44265 14843 44321
rect 161 44123 217 44179
rect 303 44123 359 44179
rect 445 44123 501 44179
rect 587 44123 643 44179
rect 729 44123 785 44179
rect 871 44123 927 44179
rect 1013 44123 1069 44179
rect 1155 44123 1211 44179
rect 1297 44123 1353 44179
rect 1439 44123 1495 44179
rect 1581 44123 1637 44179
rect 1723 44123 1779 44179
rect 1865 44123 1921 44179
rect 2007 44123 2063 44179
rect 2149 44123 2205 44179
rect 2291 44123 2347 44179
rect 2433 44123 2489 44179
rect 2575 44123 2631 44179
rect 2717 44123 2773 44179
rect 2859 44123 2915 44179
rect 3001 44123 3057 44179
rect 3143 44123 3199 44179
rect 3285 44123 3341 44179
rect 3427 44123 3483 44179
rect 3569 44123 3625 44179
rect 3711 44123 3767 44179
rect 3853 44123 3909 44179
rect 3995 44123 4051 44179
rect 4137 44123 4193 44179
rect 4279 44123 4335 44179
rect 4421 44123 4477 44179
rect 4563 44123 4619 44179
rect 4705 44123 4761 44179
rect 4847 44123 4903 44179
rect 4989 44123 5045 44179
rect 5131 44123 5187 44179
rect 5273 44123 5329 44179
rect 5415 44123 5471 44179
rect 5557 44123 5613 44179
rect 5699 44123 5755 44179
rect 5841 44123 5897 44179
rect 5983 44123 6039 44179
rect 6125 44123 6181 44179
rect 6267 44123 6323 44179
rect 6409 44123 6465 44179
rect 6551 44123 6607 44179
rect 6693 44123 6749 44179
rect 6835 44123 6891 44179
rect 6977 44123 7033 44179
rect 7119 44123 7175 44179
rect 7261 44123 7317 44179
rect 7403 44123 7459 44179
rect 7545 44123 7601 44179
rect 7687 44123 7743 44179
rect 7829 44123 7885 44179
rect 7971 44123 8027 44179
rect 8113 44123 8169 44179
rect 8255 44123 8311 44179
rect 8397 44123 8453 44179
rect 8539 44123 8595 44179
rect 8681 44123 8737 44179
rect 8823 44123 8879 44179
rect 8965 44123 9021 44179
rect 9107 44123 9163 44179
rect 9249 44123 9305 44179
rect 9391 44123 9447 44179
rect 9533 44123 9589 44179
rect 9675 44123 9731 44179
rect 9817 44123 9873 44179
rect 9959 44123 10015 44179
rect 10101 44123 10157 44179
rect 10243 44123 10299 44179
rect 10385 44123 10441 44179
rect 10527 44123 10583 44179
rect 10669 44123 10725 44179
rect 10811 44123 10867 44179
rect 10953 44123 11009 44179
rect 11095 44123 11151 44179
rect 11237 44123 11293 44179
rect 11379 44123 11435 44179
rect 11521 44123 11577 44179
rect 11663 44123 11719 44179
rect 11805 44123 11861 44179
rect 11947 44123 12003 44179
rect 12089 44123 12145 44179
rect 12231 44123 12287 44179
rect 12373 44123 12429 44179
rect 12515 44123 12571 44179
rect 12657 44123 12713 44179
rect 12799 44123 12855 44179
rect 12941 44123 12997 44179
rect 13083 44123 13139 44179
rect 13225 44123 13281 44179
rect 13367 44123 13423 44179
rect 13509 44123 13565 44179
rect 13651 44123 13707 44179
rect 13793 44123 13849 44179
rect 13935 44123 13991 44179
rect 14077 44123 14133 44179
rect 14219 44123 14275 44179
rect 14361 44123 14417 44179
rect 14503 44123 14559 44179
rect 14645 44123 14701 44179
rect 14787 44123 14843 44179
rect 161 43981 217 44037
rect 303 43981 359 44037
rect 445 43981 501 44037
rect 587 43981 643 44037
rect 729 43981 785 44037
rect 871 43981 927 44037
rect 1013 43981 1069 44037
rect 1155 43981 1211 44037
rect 1297 43981 1353 44037
rect 1439 43981 1495 44037
rect 1581 43981 1637 44037
rect 1723 43981 1779 44037
rect 1865 43981 1921 44037
rect 2007 43981 2063 44037
rect 2149 43981 2205 44037
rect 2291 43981 2347 44037
rect 2433 43981 2489 44037
rect 2575 43981 2631 44037
rect 2717 43981 2773 44037
rect 2859 43981 2915 44037
rect 3001 43981 3057 44037
rect 3143 43981 3199 44037
rect 3285 43981 3341 44037
rect 3427 43981 3483 44037
rect 3569 43981 3625 44037
rect 3711 43981 3767 44037
rect 3853 43981 3909 44037
rect 3995 43981 4051 44037
rect 4137 43981 4193 44037
rect 4279 43981 4335 44037
rect 4421 43981 4477 44037
rect 4563 43981 4619 44037
rect 4705 43981 4761 44037
rect 4847 43981 4903 44037
rect 4989 43981 5045 44037
rect 5131 43981 5187 44037
rect 5273 43981 5329 44037
rect 5415 43981 5471 44037
rect 5557 43981 5613 44037
rect 5699 43981 5755 44037
rect 5841 43981 5897 44037
rect 5983 43981 6039 44037
rect 6125 43981 6181 44037
rect 6267 43981 6323 44037
rect 6409 43981 6465 44037
rect 6551 43981 6607 44037
rect 6693 43981 6749 44037
rect 6835 43981 6891 44037
rect 6977 43981 7033 44037
rect 7119 43981 7175 44037
rect 7261 43981 7317 44037
rect 7403 43981 7459 44037
rect 7545 43981 7601 44037
rect 7687 43981 7743 44037
rect 7829 43981 7885 44037
rect 7971 43981 8027 44037
rect 8113 43981 8169 44037
rect 8255 43981 8311 44037
rect 8397 43981 8453 44037
rect 8539 43981 8595 44037
rect 8681 43981 8737 44037
rect 8823 43981 8879 44037
rect 8965 43981 9021 44037
rect 9107 43981 9163 44037
rect 9249 43981 9305 44037
rect 9391 43981 9447 44037
rect 9533 43981 9589 44037
rect 9675 43981 9731 44037
rect 9817 43981 9873 44037
rect 9959 43981 10015 44037
rect 10101 43981 10157 44037
rect 10243 43981 10299 44037
rect 10385 43981 10441 44037
rect 10527 43981 10583 44037
rect 10669 43981 10725 44037
rect 10811 43981 10867 44037
rect 10953 43981 11009 44037
rect 11095 43981 11151 44037
rect 11237 43981 11293 44037
rect 11379 43981 11435 44037
rect 11521 43981 11577 44037
rect 11663 43981 11719 44037
rect 11805 43981 11861 44037
rect 11947 43981 12003 44037
rect 12089 43981 12145 44037
rect 12231 43981 12287 44037
rect 12373 43981 12429 44037
rect 12515 43981 12571 44037
rect 12657 43981 12713 44037
rect 12799 43981 12855 44037
rect 12941 43981 12997 44037
rect 13083 43981 13139 44037
rect 13225 43981 13281 44037
rect 13367 43981 13423 44037
rect 13509 43981 13565 44037
rect 13651 43981 13707 44037
rect 13793 43981 13849 44037
rect 13935 43981 13991 44037
rect 14077 43981 14133 44037
rect 14219 43981 14275 44037
rect 14361 43981 14417 44037
rect 14503 43981 14559 44037
rect 14645 43981 14701 44037
rect 14787 43981 14843 44037
rect 161 43839 217 43895
rect 303 43839 359 43895
rect 445 43839 501 43895
rect 587 43839 643 43895
rect 729 43839 785 43895
rect 871 43839 927 43895
rect 1013 43839 1069 43895
rect 1155 43839 1211 43895
rect 1297 43839 1353 43895
rect 1439 43839 1495 43895
rect 1581 43839 1637 43895
rect 1723 43839 1779 43895
rect 1865 43839 1921 43895
rect 2007 43839 2063 43895
rect 2149 43839 2205 43895
rect 2291 43839 2347 43895
rect 2433 43839 2489 43895
rect 2575 43839 2631 43895
rect 2717 43839 2773 43895
rect 2859 43839 2915 43895
rect 3001 43839 3057 43895
rect 3143 43839 3199 43895
rect 3285 43839 3341 43895
rect 3427 43839 3483 43895
rect 3569 43839 3625 43895
rect 3711 43839 3767 43895
rect 3853 43839 3909 43895
rect 3995 43839 4051 43895
rect 4137 43839 4193 43895
rect 4279 43839 4335 43895
rect 4421 43839 4477 43895
rect 4563 43839 4619 43895
rect 4705 43839 4761 43895
rect 4847 43839 4903 43895
rect 4989 43839 5045 43895
rect 5131 43839 5187 43895
rect 5273 43839 5329 43895
rect 5415 43839 5471 43895
rect 5557 43839 5613 43895
rect 5699 43839 5755 43895
rect 5841 43839 5897 43895
rect 5983 43839 6039 43895
rect 6125 43839 6181 43895
rect 6267 43839 6323 43895
rect 6409 43839 6465 43895
rect 6551 43839 6607 43895
rect 6693 43839 6749 43895
rect 6835 43839 6891 43895
rect 6977 43839 7033 43895
rect 7119 43839 7175 43895
rect 7261 43839 7317 43895
rect 7403 43839 7459 43895
rect 7545 43839 7601 43895
rect 7687 43839 7743 43895
rect 7829 43839 7885 43895
rect 7971 43839 8027 43895
rect 8113 43839 8169 43895
rect 8255 43839 8311 43895
rect 8397 43839 8453 43895
rect 8539 43839 8595 43895
rect 8681 43839 8737 43895
rect 8823 43839 8879 43895
rect 8965 43839 9021 43895
rect 9107 43839 9163 43895
rect 9249 43839 9305 43895
rect 9391 43839 9447 43895
rect 9533 43839 9589 43895
rect 9675 43839 9731 43895
rect 9817 43839 9873 43895
rect 9959 43839 10015 43895
rect 10101 43839 10157 43895
rect 10243 43839 10299 43895
rect 10385 43839 10441 43895
rect 10527 43839 10583 43895
rect 10669 43839 10725 43895
rect 10811 43839 10867 43895
rect 10953 43839 11009 43895
rect 11095 43839 11151 43895
rect 11237 43839 11293 43895
rect 11379 43839 11435 43895
rect 11521 43839 11577 43895
rect 11663 43839 11719 43895
rect 11805 43839 11861 43895
rect 11947 43839 12003 43895
rect 12089 43839 12145 43895
rect 12231 43839 12287 43895
rect 12373 43839 12429 43895
rect 12515 43839 12571 43895
rect 12657 43839 12713 43895
rect 12799 43839 12855 43895
rect 12941 43839 12997 43895
rect 13083 43839 13139 43895
rect 13225 43839 13281 43895
rect 13367 43839 13423 43895
rect 13509 43839 13565 43895
rect 13651 43839 13707 43895
rect 13793 43839 13849 43895
rect 13935 43839 13991 43895
rect 14077 43839 14133 43895
rect 14219 43839 14275 43895
rect 14361 43839 14417 43895
rect 14503 43839 14559 43895
rect 14645 43839 14701 43895
rect 14787 43839 14843 43895
rect 161 43697 217 43753
rect 303 43697 359 43753
rect 445 43697 501 43753
rect 587 43697 643 43753
rect 729 43697 785 43753
rect 871 43697 927 43753
rect 1013 43697 1069 43753
rect 1155 43697 1211 43753
rect 1297 43697 1353 43753
rect 1439 43697 1495 43753
rect 1581 43697 1637 43753
rect 1723 43697 1779 43753
rect 1865 43697 1921 43753
rect 2007 43697 2063 43753
rect 2149 43697 2205 43753
rect 2291 43697 2347 43753
rect 2433 43697 2489 43753
rect 2575 43697 2631 43753
rect 2717 43697 2773 43753
rect 2859 43697 2915 43753
rect 3001 43697 3057 43753
rect 3143 43697 3199 43753
rect 3285 43697 3341 43753
rect 3427 43697 3483 43753
rect 3569 43697 3625 43753
rect 3711 43697 3767 43753
rect 3853 43697 3909 43753
rect 3995 43697 4051 43753
rect 4137 43697 4193 43753
rect 4279 43697 4335 43753
rect 4421 43697 4477 43753
rect 4563 43697 4619 43753
rect 4705 43697 4761 43753
rect 4847 43697 4903 43753
rect 4989 43697 5045 43753
rect 5131 43697 5187 43753
rect 5273 43697 5329 43753
rect 5415 43697 5471 43753
rect 5557 43697 5613 43753
rect 5699 43697 5755 43753
rect 5841 43697 5897 43753
rect 5983 43697 6039 43753
rect 6125 43697 6181 43753
rect 6267 43697 6323 43753
rect 6409 43697 6465 43753
rect 6551 43697 6607 43753
rect 6693 43697 6749 43753
rect 6835 43697 6891 43753
rect 6977 43697 7033 43753
rect 7119 43697 7175 43753
rect 7261 43697 7317 43753
rect 7403 43697 7459 43753
rect 7545 43697 7601 43753
rect 7687 43697 7743 43753
rect 7829 43697 7885 43753
rect 7971 43697 8027 43753
rect 8113 43697 8169 43753
rect 8255 43697 8311 43753
rect 8397 43697 8453 43753
rect 8539 43697 8595 43753
rect 8681 43697 8737 43753
rect 8823 43697 8879 43753
rect 8965 43697 9021 43753
rect 9107 43697 9163 43753
rect 9249 43697 9305 43753
rect 9391 43697 9447 43753
rect 9533 43697 9589 43753
rect 9675 43697 9731 43753
rect 9817 43697 9873 43753
rect 9959 43697 10015 43753
rect 10101 43697 10157 43753
rect 10243 43697 10299 43753
rect 10385 43697 10441 43753
rect 10527 43697 10583 43753
rect 10669 43697 10725 43753
rect 10811 43697 10867 43753
rect 10953 43697 11009 43753
rect 11095 43697 11151 43753
rect 11237 43697 11293 43753
rect 11379 43697 11435 43753
rect 11521 43697 11577 43753
rect 11663 43697 11719 43753
rect 11805 43697 11861 43753
rect 11947 43697 12003 43753
rect 12089 43697 12145 43753
rect 12231 43697 12287 43753
rect 12373 43697 12429 43753
rect 12515 43697 12571 43753
rect 12657 43697 12713 43753
rect 12799 43697 12855 43753
rect 12941 43697 12997 43753
rect 13083 43697 13139 43753
rect 13225 43697 13281 43753
rect 13367 43697 13423 43753
rect 13509 43697 13565 43753
rect 13651 43697 13707 43753
rect 13793 43697 13849 43753
rect 13935 43697 13991 43753
rect 14077 43697 14133 43753
rect 14219 43697 14275 43753
rect 14361 43697 14417 43753
rect 14503 43697 14559 43753
rect 14645 43697 14701 43753
rect 14787 43697 14843 43753
rect 161 43555 217 43611
rect 303 43555 359 43611
rect 445 43555 501 43611
rect 587 43555 643 43611
rect 729 43555 785 43611
rect 871 43555 927 43611
rect 1013 43555 1069 43611
rect 1155 43555 1211 43611
rect 1297 43555 1353 43611
rect 1439 43555 1495 43611
rect 1581 43555 1637 43611
rect 1723 43555 1779 43611
rect 1865 43555 1921 43611
rect 2007 43555 2063 43611
rect 2149 43555 2205 43611
rect 2291 43555 2347 43611
rect 2433 43555 2489 43611
rect 2575 43555 2631 43611
rect 2717 43555 2773 43611
rect 2859 43555 2915 43611
rect 3001 43555 3057 43611
rect 3143 43555 3199 43611
rect 3285 43555 3341 43611
rect 3427 43555 3483 43611
rect 3569 43555 3625 43611
rect 3711 43555 3767 43611
rect 3853 43555 3909 43611
rect 3995 43555 4051 43611
rect 4137 43555 4193 43611
rect 4279 43555 4335 43611
rect 4421 43555 4477 43611
rect 4563 43555 4619 43611
rect 4705 43555 4761 43611
rect 4847 43555 4903 43611
rect 4989 43555 5045 43611
rect 5131 43555 5187 43611
rect 5273 43555 5329 43611
rect 5415 43555 5471 43611
rect 5557 43555 5613 43611
rect 5699 43555 5755 43611
rect 5841 43555 5897 43611
rect 5983 43555 6039 43611
rect 6125 43555 6181 43611
rect 6267 43555 6323 43611
rect 6409 43555 6465 43611
rect 6551 43555 6607 43611
rect 6693 43555 6749 43611
rect 6835 43555 6891 43611
rect 6977 43555 7033 43611
rect 7119 43555 7175 43611
rect 7261 43555 7317 43611
rect 7403 43555 7459 43611
rect 7545 43555 7601 43611
rect 7687 43555 7743 43611
rect 7829 43555 7885 43611
rect 7971 43555 8027 43611
rect 8113 43555 8169 43611
rect 8255 43555 8311 43611
rect 8397 43555 8453 43611
rect 8539 43555 8595 43611
rect 8681 43555 8737 43611
rect 8823 43555 8879 43611
rect 8965 43555 9021 43611
rect 9107 43555 9163 43611
rect 9249 43555 9305 43611
rect 9391 43555 9447 43611
rect 9533 43555 9589 43611
rect 9675 43555 9731 43611
rect 9817 43555 9873 43611
rect 9959 43555 10015 43611
rect 10101 43555 10157 43611
rect 10243 43555 10299 43611
rect 10385 43555 10441 43611
rect 10527 43555 10583 43611
rect 10669 43555 10725 43611
rect 10811 43555 10867 43611
rect 10953 43555 11009 43611
rect 11095 43555 11151 43611
rect 11237 43555 11293 43611
rect 11379 43555 11435 43611
rect 11521 43555 11577 43611
rect 11663 43555 11719 43611
rect 11805 43555 11861 43611
rect 11947 43555 12003 43611
rect 12089 43555 12145 43611
rect 12231 43555 12287 43611
rect 12373 43555 12429 43611
rect 12515 43555 12571 43611
rect 12657 43555 12713 43611
rect 12799 43555 12855 43611
rect 12941 43555 12997 43611
rect 13083 43555 13139 43611
rect 13225 43555 13281 43611
rect 13367 43555 13423 43611
rect 13509 43555 13565 43611
rect 13651 43555 13707 43611
rect 13793 43555 13849 43611
rect 13935 43555 13991 43611
rect 14077 43555 14133 43611
rect 14219 43555 14275 43611
rect 14361 43555 14417 43611
rect 14503 43555 14559 43611
rect 14645 43555 14701 43611
rect 14787 43555 14843 43611
rect 161 43413 217 43469
rect 303 43413 359 43469
rect 445 43413 501 43469
rect 587 43413 643 43469
rect 729 43413 785 43469
rect 871 43413 927 43469
rect 1013 43413 1069 43469
rect 1155 43413 1211 43469
rect 1297 43413 1353 43469
rect 1439 43413 1495 43469
rect 1581 43413 1637 43469
rect 1723 43413 1779 43469
rect 1865 43413 1921 43469
rect 2007 43413 2063 43469
rect 2149 43413 2205 43469
rect 2291 43413 2347 43469
rect 2433 43413 2489 43469
rect 2575 43413 2631 43469
rect 2717 43413 2773 43469
rect 2859 43413 2915 43469
rect 3001 43413 3057 43469
rect 3143 43413 3199 43469
rect 3285 43413 3341 43469
rect 3427 43413 3483 43469
rect 3569 43413 3625 43469
rect 3711 43413 3767 43469
rect 3853 43413 3909 43469
rect 3995 43413 4051 43469
rect 4137 43413 4193 43469
rect 4279 43413 4335 43469
rect 4421 43413 4477 43469
rect 4563 43413 4619 43469
rect 4705 43413 4761 43469
rect 4847 43413 4903 43469
rect 4989 43413 5045 43469
rect 5131 43413 5187 43469
rect 5273 43413 5329 43469
rect 5415 43413 5471 43469
rect 5557 43413 5613 43469
rect 5699 43413 5755 43469
rect 5841 43413 5897 43469
rect 5983 43413 6039 43469
rect 6125 43413 6181 43469
rect 6267 43413 6323 43469
rect 6409 43413 6465 43469
rect 6551 43413 6607 43469
rect 6693 43413 6749 43469
rect 6835 43413 6891 43469
rect 6977 43413 7033 43469
rect 7119 43413 7175 43469
rect 7261 43413 7317 43469
rect 7403 43413 7459 43469
rect 7545 43413 7601 43469
rect 7687 43413 7743 43469
rect 7829 43413 7885 43469
rect 7971 43413 8027 43469
rect 8113 43413 8169 43469
rect 8255 43413 8311 43469
rect 8397 43413 8453 43469
rect 8539 43413 8595 43469
rect 8681 43413 8737 43469
rect 8823 43413 8879 43469
rect 8965 43413 9021 43469
rect 9107 43413 9163 43469
rect 9249 43413 9305 43469
rect 9391 43413 9447 43469
rect 9533 43413 9589 43469
rect 9675 43413 9731 43469
rect 9817 43413 9873 43469
rect 9959 43413 10015 43469
rect 10101 43413 10157 43469
rect 10243 43413 10299 43469
rect 10385 43413 10441 43469
rect 10527 43413 10583 43469
rect 10669 43413 10725 43469
rect 10811 43413 10867 43469
rect 10953 43413 11009 43469
rect 11095 43413 11151 43469
rect 11237 43413 11293 43469
rect 11379 43413 11435 43469
rect 11521 43413 11577 43469
rect 11663 43413 11719 43469
rect 11805 43413 11861 43469
rect 11947 43413 12003 43469
rect 12089 43413 12145 43469
rect 12231 43413 12287 43469
rect 12373 43413 12429 43469
rect 12515 43413 12571 43469
rect 12657 43413 12713 43469
rect 12799 43413 12855 43469
rect 12941 43413 12997 43469
rect 13083 43413 13139 43469
rect 13225 43413 13281 43469
rect 13367 43413 13423 43469
rect 13509 43413 13565 43469
rect 13651 43413 13707 43469
rect 13793 43413 13849 43469
rect 13935 43413 13991 43469
rect 14077 43413 14133 43469
rect 14219 43413 14275 43469
rect 14361 43413 14417 43469
rect 14503 43413 14559 43469
rect 14645 43413 14701 43469
rect 14787 43413 14843 43469
rect 161 43271 217 43327
rect 303 43271 359 43327
rect 445 43271 501 43327
rect 587 43271 643 43327
rect 729 43271 785 43327
rect 871 43271 927 43327
rect 1013 43271 1069 43327
rect 1155 43271 1211 43327
rect 1297 43271 1353 43327
rect 1439 43271 1495 43327
rect 1581 43271 1637 43327
rect 1723 43271 1779 43327
rect 1865 43271 1921 43327
rect 2007 43271 2063 43327
rect 2149 43271 2205 43327
rect 2291 43271 2347 43327
rect 2433 43271 2489 43327
rect 2575 43271 2631 43327
rect 2717 43271 2773 43327
rect 2859 43271 2915 43327
rect 3001 43271 3057 43327
rect 3143 43271 3199 43327
rect 3285 43271 3341 43327
rect 3427 43271 3483 43327
rect 3569 43271 3625 43327
rect 3711 43271 3767 43327
rect 3853 43271 3909 43327
rect 3995 43271 4051 43327
rect 4137 43271 4193 43327
rect 4279 43271 4335 43327
rect 4421 43271 4477 43327
rect 4563 43271 4619 43327
rect 4705 43271 4761 43327
rect 4847 43271 4903 43327
rect 4989 43271 5045 43327
rect 5131 43271 5187 43327
rect 5273 43271 5329 43327
rect 5415 43271 5471 43327
rect 5557 43271 5613 43327
rect 5699 43271 5755 43327
rect 5841 43271 5897 43327
rect 5983 43271 6039 43327
rect 6125 43271 6181 43327
rect 6267 43271 6323 43327
rect 6409 43271 6465 43327
rect 6551 43271 6607 43327
rect 6693 43271 6749 43327
rect 6835 43271 6891 43327
rect 6977 43271 7033 43327
rect 7119 43271 7175 43327
rect 7261 43271 7317 43327
rect 7403 43271 7459 43327
rect 7545 43271 7601 43327
rect 7687 43271 7743 43327
rect 7829 43271 7885 43327
rect 7971 43271 8027 43327
rect 8113 43271 8169 43327
rect 8255 43271 8311 43327
rect 8397 43271 8453 43327
rect 8539 43271 8595 43327
rect 8681 43271 8737 43327
rect 8823 43271 8879 43327
rect 8965 43271 9021 43327
rect 9107 43271 9163 43327
rect 9249 43271 9305 43327
rect 9391 43271 9447 43327
rect 9533 43271 9589 43327
rect 9675 43271 9731 43327
rect 9817 43271 9873 43327
rect 9959 43271 10015 43327
rect 10101 43271 10157 43327
rect 10243 43271 10299 43327
rect 10385 43271 10441 43327
rect 10527 43271 10583 43327
rect 10669 43271 10725 43327
rect 10811 43271 10867 43327
rect 10953 43271 11009 43327
rect 11095 43271 11151 43327
rect 11237 43271 11293 43327
rect 11379 43271 11435 43327
rect 11521 43271 11577 43327
rect 11663 43271 11719 43327
rect 11805 43271 11861 43327
rect 11947 43271 12003 43327
rect 12089 43271 12145 43327
rect 12231 43271 12287 43327
rect 12373 43271 12429 43327
rect 12515 43271 12571 43327
rect 12657 43271 12713 43327
rect 12799 43271 12855 43327
rect 12941 43271 12997 43327
rect 13083 43271 13139 43327
rect 13225 43271 13281 43327
rect 13367 43271 13423 43327
rect 13509 43271 13565 43327
rect 13651 43271 13707 43327
rect 13793 43271 13849 43327
rect 13935 43271 13991 43327
rect 14077 43271 14133 43327
rect 14219 43271 14275 43327
rect 14361 43271 14417 43327
rect 14503 43271 14559 43327
rect 14645 43271 14701 43327
rect 14787 43271 14843 43327
rect 161 43129 217 43185
rect 303 43129 359 43185
rect 445 43129 501 43185
rect 587 43129 643 43185
rect 729 43129 785 43185
rect 871 43129 927 43185
rect 1013 43129 1069 43185
rect 1155 43129 1211 43185
rect 1297 43129 1353 43185
rect 1439 43129 1495 43185
rect 1581 43129 1637 43185
rect 1723 43129 1779 43185
rect 1865 43129 1921 43185
rect 2007 43129 2063 43185
rect 2149 43129 2205 43185
rect 2291 43129 2347 43185
rect 2433 43129 2489 43185
rect 2575 43129 2631 43185
rect 2717 43129 2773 43185
rect 2859 43129 2915 43185
rect 3001 43129 3057 43185
rect 3143 43129 3199 43185
rect 3285 43129 3341 43185
rect 3427 43129 3483 43185
rect 3569 43129 3625 43185
rect 3711 43129 3767 43185
rect 3853 43129 3909 43185
rect 3995 43129 4051 43185
rect 4137 43129 4193 43185
rect 4279 43129 4335 43185
rect 4421 43129 4477 43185
rect 4563 43129 4619 43185
rect 4705 43129 4761 43185
rect 4847 43129 4903 43185
rect 4989 43129 5045 43185
rect 5131 43129 5187 43185
rect 5273 43129 5329 43185
rect 5415 43129 5471 43185
rect 5557 43129 5613 43185
rect 5699 43129 5755 43185
rect 5841 43129 5897 43185
rect 5983 43129 6039 43185
rect 6125 43129 6181 43185
rect 6267 43129 6323 43185
rect 6409 43129 6465 43185
rect 6551 43129 6607 43185
rect 6693 43129 6749 43185
rect 6835 43129 6891 43185
rect 6977 43129 7033 43185
rect 7119 43129 7175 43185
rect 7261 43129 7317 43185
rect 7403 43129 7459 43185
rect 7545 43129 7601 43185
rect 7687 43129 7743 43185
rect 7829 43129 7885 43185
rect 7971 43129 8027 43185
rect 8113 43129 8169 43185
rect 8255 43129 8311 43185
rect 8397 43129 8453 43185
rect 8539 43129 8595 43185
rect 8681 43129 8737 43185
rect 8823 43129 8879 43185
rect 8965 43129 9021 43185
rect 9107 43129 9163 43185
rect 9249 43129 9305 43185
rect 9391 43129 9447 43185
rect 9533 43129 9589 43185
rect 9675 43129 9731 43185
rect 9817 43129 9873 43185
rect 9959 43129 10015 43185
rect 10101 43129 10157 43185
rect 10243 43129 10299 43185
rect 10385 43129 10441 43185
rect 10527 43129 10583 43185
rect 10669 43129 10725 43185
rect 10811 43129 10867 43185
rect 10953 43129 11009 43185
rect 11095 43129 11151 43185
rect 11237 43129 11293 43185
rect 11379 43129 11435 43185
rect 11521 43129 11577 43185
rect 11663 43129 11719 43185
rect 11805 43129 11861 43185
rect 11947 43129 12003 43185
rect 12089 43129 12145 43185
rect 12231 43129 12287 43185
rect 12373 43129 12429 43185
rect 12515 43129 12571 43185
rect 12657 43129 12713 43185
rect 12799 43129 12855 43185
rect 12941 43129 12997 43185
rect 13083 43129 13139 43185
rect 13225 43129 13281 43185
rect 13367 43129 13423 43185
rect 13509 43129 13565 43185
rect 13651 43129 13707 43185
rect 13793 43129 13849 43185
rect 13935 43129 13991 43185
rect 14077 43129 14133 43185
rect 14219 43129 14275 43185
rect 14361 43129 14417 43185
rect 14503 43129 14559 43185
rect 14645 43129 14701 43185
rect 14787 43129 14843 43185
rect 161 42987 217 43043
rect 303 42987 359 43043
rect 445 42987 501 43043
rect 587 42987 643 43043
rect 729 42987 785 43043
rect 871 42987 927 43043
rect 1013 42987 1069 43043
rect 1155 42987 1211 43043
rect 1297 42987 1353 43043
rect 1439 42987 1495 43043
rect 1581 42987 1637 43043
rect 1723 42987 1779 43043
rect 1865 42987 1921 43043
rect 2007 42987 2063 43043
rect 2149 42987 2205 43043
rect 2291 42987 2347 43043
rect 2433 42987 2489 43043
rect 2575 42987 2631 43043
rect 2717 42987 2773 43043
rect 2859 42987 2915 43043
rect 3001 42987 3057 43043
rect 3143 42987 3199 43043
rect 3285 42987 3341 43043
rect 3427 42987 3483 43043
rect 3569 42987 3625 43043
rect 3711 42987 3767 43043
rect 3853 42987 3909 43043
rect 3995 42987 4051 43043
rect 4137 42987 4193 43043
rect 4279 42987 4335 43043
rect 4421 42987 4477 43043
rect 4563 42987 4619 43043
rect 4705 42987 4761 43043
rect 4847 42987 4903 43043
rect 4989 42987 5045 43043
rect 5131 42987 5187 43043
rect 5273 42987 5329 43043
rect 5415 42987 5471 43043
rect 5557 42987 5613 43043
rect 5699 42987 5755 43043
rect 5841 42987 5897 43043
rect 5983 42987 6039 43043
rect 6125 42987 6181 43043
rect 6267 42987 6323 43043
rect 6409 42987 6465 43043
rect 6551 42987 6607 43043
rect 6693 42987 6749 43043
rect 6835 42987 6891 43043
rect 6977 42987 7033 43043
rect 7119 42987 7175 43043
rect 7261 42987 7317 43043
rect 7403 42987 7459 43043
rect 7545 42987 7601 43043
rect 7687 42987 7743 43043
rect 7829 42987 7885 43043
rect 7971 42987 8027 43043
rect 8113 42987 8169 43043
rect 8255 42987 8311 43043
rect 8397 42987 8453 43043
rect 8539 42987 8595 43043
rect 8681 42987 8737 43043
rect 8823 42987 8879 43043
rect 8965 42987 9021 43043
rect 9107 42987 9163 43043
rect 9249 42987 9305 43043
rect 9391 42987 9447 43043
rect 9533 42987 9589 43043
rect 9675 42987 9731 43043
rect 9817 42987 9873 43043
rect 9959 42987 10015 43043
rect 10101 42987 10157 43043
rect 10243 42987 10299 43043
rect 10385 42987 10441 43043
rect 10527 42987 10583 43043
rect 10669 42987 10725 43043
rect 10811 42987 10867 43043
rect 10953 42987 11009 43043
rect 11095 42987 11151 43043
rect 11237 42987 11293 43043
rect 11379 42987 11435 43043
rect 11521 42987 11577 43043
rect 11663 42987 11719 43043
rect 11805 42987 11861 43043
rect 11947 42987 12003 43043
rect 12089 42987 12145 43043
rect 12231 42987 12287 43043
rect 12373 42987 12429 43043
rect 12515 42987 12571 43043
rect 12657 42987 12713 43043
rect 12799 42987 12855 43043
rect 12941 42987 12997 43043
rect 13083 42987 13139 43043
rect 13225 42987 13281 43043
rect 13367 42987 13423 43043
rect 13509 42987 13565 43043
rect 13651 42987 13707 43043
rect 13793 42987 13849 43043
rect 13935 42987 13991 43043
rect 14077 42987 14133 43043
rect 14219 42987 14275 43043
rect 14361 42987 14417 43043
rect 14503 42987 14559 43043
rect 14645 42987 14701 43043
rect 14787 42987 14843 43043
rect 161 42845 217 42901
rect 303 42845 359 42901
rect 445 42845 501 42901
rect 587 42845 643 42901
rect 729 42845 785 42901
rect 871 42845 927 42901
rect 1013 42845 1069 42901
rect 1155 42845 1211 42901
rect 1297 42845 1353 42901
rect 1439 42845 1495 42901
rect 1581 42845 1637 42901
rect 1723 42845 1779 42901
rect 1865 42845 1921 42901
rect 2007 42845 2063 42901
rect 2149 42845 2205 42901
rect 2291 42845 2347 42901
rect 2433 42845 2489 42901
rect 2575 42845 2631 42901
rect 2717 42845 2773 42901
rect 2859 42845 2915 42901
rect 3001 42845 3057 42901
rect 3143 42845 3199 42901
rect 3285 42845 3341 42901
rect 3427 42845 3483 42901
rect 3569 42845 3625 42901
rect 3711 42845 3767 42901
rect 3853 42845 3909 42901
rect 3995 42845 4051 42901
rect 4137 42845 4193 42901
rect 4279 42845 4335 42901
rect 4421 42845 4477 42901
rect 4563 42845 4619 42901
rect 4705 42845 4761 42901
rect 4847 42845 4903 42901
rect 4989 42845 5045 42901
rect 5131 42845 5187 42901
rect 5273 42845 5329 42901
rect 5415 42845 5471 42901
rect 5557 42845 5613 42901
rect 5699 42845 5755 42901
rect 5841 42845 5897 42901
rect 5983 42845 6039 42901
rect 6125 42845 6181 42901
rect 6267 42845 6323 42901
rect 6409 42845 6465 42901
rect 6551 42845 6607 42901
rect 6693 42845 6749 42901
rect 6835 42845 6891 42901
rect 6977 42845 7033 42901
rect 7119 42845 7175 42901
rect 7261 42845 7317 42901
rect 7403 42845 7459 42901
rect 7545 42845 7601 42901
rect 7687 42845 7743 42901
rect 7829 42845 7885 42901
rect 7971 42845 8027 42901
rect 8113 42845 8169 42901
rect 8255 42845 8311 42901
rect 8397 42845 8453 42901
rect 8539 42845 8595 42901
rect 8681 42845 8737 42901
rect 8823 42845 8879 42901
rect 8965 42845 9021 42901
rect 9107 42845 9163 42901
rect 9249 42845 9305 42901
rect 9391 42845 9447 42901
rect 9533 42845 9589 42901
rect 9675 42845 9731 42901
rect 9817 42845 9873 42901
rect 9959 42845 10015 42901
rect 10101 42845 10157 42901
rect 10243 42845 10299 42901
rect 10385 42845 10441 42901
rect 10527 42845 10583 42901
rect 10669 42845 10725 42901
rect 10811 42845 10867 42901
rect 10953 42845 11009 42901
rect 11095 42845 11151 42901
rect 11237 42845 11293 42901
rect 11379 42845 11435 42901
rect 11521 42845 11577 42901
rect 11663 42845 11719 42901
rect 11805 42845 11861 42901
rect 11947 42845 12003 42901
rect 12089 42845 12145 42901
rect 12231 42845 12287 42901
rect 12373 42845 12429 42901
rect 12515 42845 12571 42901
rect 12657 42845 12713 42901
rect 12799 42845 12855 42901
rect 12941 42845 12997 42901
rect 13083 42845 13139 42901
rect 13225 42845 13281 42901
rect 13367 42845 13423 42901
rect 13509 42845 13565 42901
rect 13651 42845 13707 42901
rect 13793 42845 13849 42901
rect 13935 42845 13991 42901
rect 14077 42845 14133 42901
rect 14219 42845 14275 42901
rect 14361 42845 14417 42901
rect 14503 42845 14559 42901
rect 14645 42845 14701 42901
rect 14787 42845 14843 42901
rect 161 42507 217 42563
rect 303 42507 359 42563
rect 445 42507 501 42563
rect 587 42507 643 42563
rect 729 42507 785 42563
rect 871 42507 927 42563
rect 1013 42507 1069 42563
rect 1155 42507 1211 42563
rect 1297 42507 1353 42563
rect 1439 42507 1495 42563
rect 1581 42507 1637 42563
rect 1723 42507 1779 42563
rect 1865 42507 1921 42563
rect 2007 42507 2063 42563
rect 2149 42507 2205 42563
rect 2291 42507 2347 42563
rect 2433 42507 2489 42563
rect 2575 42507 2631 42563
rect 2717 42507 2773 42563
rect 2859 42507 2915 42563
rect 3001 42507 3057 42563
rect 3143 42507 3199 42563
rect 3285 42507 3341 42563
rect 3427 42507 3483 42563
rect 3569 42507 3625 42563
rect 3711 42507 3767 42563
rect 3853 42507 3909 42563
rect 3995 42507 4051 42563
rect 4137 42507 4193 42563
rect 4279 42507 4335 42563
rect 4421 42507 4477 42563
rect 4563 42507 4619 42563
rect 4705 42507 4761 42563
rect 4847 42507 4903 42563
rect 4989 42507 5045 42563
rect 5131 42507 5187 42563
rect 5273 42507 5329 42563
rect 5415 42507 5471 42563
rect 5557 42507 5613 42563
rect 5699 42507 5755 42563
rect 5841 42507 5897 42563
rect 5983 42507 6039 42563
rect 6125 42507 6181 42563
rect 6267 42507 6323 42563
rect 6409 42507 6465 42563
rect 6551 42507 6607 42563
rect 6693 42507 6749 42563
rect 6835 42507 6891 42563
rect 6977 42507 7033 42563
rect 7119 42507 7175 42563
rect 7261 42507 7317 42563
rect 7403 42507 7459 42563
rect 7545 42507 7601 42563
rect 7687 42507 7743 42563
rect 7829 42507 7885 42563
rect 7971 42507 8027 42563
rect 8113 42507 8169 42563
rect 8255 42507 8311 42563
rect 8397 42507 8453 42563
rect 8539 42507 8595 42563
rect 8681 42507 8737 42563
rect 8823 42507 8879 42563
rect 8965 42507 9021 42563
rect 9107 42507 9163 42563
rect 9249 42507 9305 42563
rect 9391 42507 9447 42563
rect 9533 42507 9589 42563
rect 9675 42507 9731 42563
rect 9817 42507 9873 42563
rect 9959 42507 10015 42563
rect 10101 42507 10157 42563
rect 10243 42507 10299 42563
rect 10385 42507 10441 42563
rect 10527 42507 10583 42563
rect 10669 42507 10725 42563
rect 10811 42507 10867 42563
rect 10953 42507 11009 42563
rect 11095 42507 11151 42563
rect 11237 42507 11293 42563
rect 11379 42507 11435 42563
rect 11521 42507 11577 42563
rect 11663 42507 11719 42563
rect 11805 42507 11861 42563
rect 11947 42507 12003 42563
rect 12089 42507 12145 42563
rect 12231 42507 12287 42563
rect 12373 42507 12429 42563
rect 12515 42507 12571 42563
rect 12657 42507 12713 42563
rect 12799 42507 12855 42563
rect 12941 42507 12997 42563
rect 13083 42507 13139 42563
rect 13225 42507 13281 42563
rect 13367 42507 13423 42563
rect 13509 42507 13565 42563
rect 13651 42507 13707 42563
rect 13793 42507 13849 42563
rect 13935 42507 13991 42563
rect 14077 42507 14133 42563
rect 14219 42507 14275 42563
rect 14361 42507 14417 42563
rect 14503 42507 14559 42563
rect 14645 42507 14701 42563
rect 14787 42507 14843 42563
rect 161 42365 217 42421
rect 303 42365 359 42421
rect 445 42365 501 42421
rect 587 42365 643 42421
rect 729 42365 785 42421
rect 871 42365 927 42421
rect 1013 42365 1069 42421
rect 1155 42365 1211 42421
rect 1297 42365 1353 42421
rect 1439 42365 1495 42421
rect 1581 42365 1637 42421
rect 1723 42365 1779 42421
rect 1865 42365 1921 42421
rect 2007 42365 2063 42421
rect 2149 42365 2205 42421
rect 2291 42365 2347 42421
rect 2433 42365 2489 42421
rect 2575 42365 2631 42421
rect 2717 42365 2773 42421
rect 2859 42365 2915 42421
rect 3001 42365 3057 42421
rect 3143 42365 3199 42421
rect 3285 42365 3341 42421
rect 3427 42365 3483 42421
rect 3569 42365 3625 42421
rect 3711 42365 3767 42421
rect 3853 42365 3909 42421
rect 3995 42365 4051 42421
rect 4137 42365 4193 42421
rect 4279 42365 4335 42421
rect 4421 42365 4477 42421
rect 4563 42365 4619 42421
rect 4705 42365 4761 42421
rect 4847 42365 4903 42421
rect 4989 42365 5045 42421
rect 5131 42365 5187 42421
rect 5273 42365 5329 42421
rect 5415 42365 5471 42421
rect 5557 42365 5613 42421
rect 5699 42365 5755 42421
rect 5841 42365 5897 42421
rect 5983 42365 6039 42421
rect 6125 42365 6181 42421
rect 6267 42365 6323 42421
rect 6409 42365 6465 42421
rect 6551 42365 6607 42421
rect 6693 42365 6749 42421
rect 6835 42365 6891 42421
rect 6977 42365 7033 42421
rect 7119 42365 7175 42421
rect 7261 42365 7317 42421
rect 7403 42365 7459 42421
rect 7545 42365 7601 42421
rect 7687 42365 7743 42421
rect 7829 42365 7885 42421
rect 7971 42365 8027 42421
rect 8113 42365 8169 42421
rect 8255 42365 8311 42421
rect 8397 42365 8453 42421
rect 8539 42365 8595 42421
rect 8681 42365 8737 42421
rect 8823 42365 8879 42421
rect 8965 42365 9021 42421
rect 9107 42365 9163 42421
rect 9249 42365 9305 42421
rect 9391 42365 9447 42421
rect 9533 42365 9589 42421
rect 9675 42365 9731 42421
rect 9817 42365 9873 42421
rect 9959 42365 10015 42421
rect 10101 42365 10157 42421
rect 10243 42365 10299 42421
rect 10385 42365 10441 42421
rect 10527 42365 10583 42421
rect 10669 42365 10725 42421
rect 10811 42365 10867 42421
rect 10953 42365 11009 42421
rect 11095 42365 11151 42421
rect 11237 42365 11293 42421
rect 11379 42365 11435 42421
rect 11521 42365 11577 42421
rect 11663 42365 11719 42421
rect 11805 42365 11861 42421
rect 11947 42365 12003 42421
rect 12089 42365 12145 42421
rect 12231 42365 12287 42421
rect 12373 42365 12429 42421
rect 12515 42365 12571 42421
rect 12657 42365 12713 42421
rect 12799 42365 12855 42421
rect 12941 42365 12997 42421
rect 13083 42365 13139 42421
rect 13225 42365 13281 42421
rect 13367 42365 13423 42421
rect 13509 42365 13565 42421
rect 13651 42365 13707 42421
rect 13793 42365 13849 42421
rect 13935 42365 13991 42421
rect 14077 42365 14133 42421
rect 14219 42365 14275 42421
rect 14361 42365 14417 42421
rect 14503 42365 14559 42421
rect 14645 42365 14701 42421
rect 14787 42365 14843 42421
rect 161 42223 217 42279
rect 303 42223 359 42279
rect 445 42223 501 42279
rect 587 42223 643 42279
rect 729 42223 785 42279
rect 871 42223 927 42279
rect 1013 42223 1069 42279
rect 1155 42223 1211 42279
rect 1297 42223 1353 42279
rect 1439 42223 1495 42279
rect 1581 42223 1637 42279
rect 1723 42223 1779 42279
rect 1865 42223 1921 42279
rect 2007 42223 2063 42279
rect 2149 42223 2205 42279
rect 2291 42223 2347 42279
rect 2433 42223 2489 42279
rect 2575 42223 2631 42279
rect 2717 42223 2773 42279
rect 2859 42223 2915 42279
rect 3001 42223 3057 42279
rect 3143 42223 3199 42279
rect 3285 42223 3341 42279
rect 3427 42223 3483 42279
rect 3569 42223 3625 42279
rect 3711 42223 3767 42279
rect 3853 42223 3909 42279
rect 3995 42223 4051 42279
rect 4137 42223 4193 42279
rect 4279 42223 4335 42279
rect 4421 42223 4477 42279
rect 4563 42223 4619 42279
rect 4705 42223 4761 42279
rect 4847 42223 4903 42279
rect 4989 42223 5045 42279
rect 5131 42223 5187 42279
rect 5273 42223 5329 42279
rect 5415 42223 5471 42279
rect 5557 42223 5613 42279
rect 5699 42223 5755 42279
rect 5841 42223 5897 42279
rect 5983 42223 6039 42279
rect 6125 42223 6181 42279
rect 6267 42223 6323 42279
rect 6409 42223 6465 42279
rect 6551 42223 6607 42279
rect 6693 42223 6749 42279
rect 6835 42223 6891 42279
rect 6977 42223 7033 42279
rect 7119 42223 7175 42279
rect 7261 42223 7317 42279
rect 7403 42223 7459 42279
rect 7545 42223 7601 42279
rect 7687 42223 7743 42279
rect 7829 42223 7885 42279
rect 7971 42223 8027 42279
rect 8113 42223 8169 42279
rect 8255 42223 8311 42279
rect 8397 42223 8453 42279
rect 8539 42223 8595 42279
rect 8681 42223 8737 42279
rect 8823 42223 8879 42279
rect 8965 42223 9021 42279
rect 9107 42223 9163 42279
rect 9249 42223 9305 42279
rect 9391 42223 9447 42279
rect 9533 42223 9589 42279
rect 9675 42223 9731 42279
rect 9817 42223 9873 42279
rect 9959 42223 10015 42279
rect 10101 42223 10157 42279
rect 10243 42223 10299 42279
rect 10385 42223 10441 42279
rect 10527 42223 10583 42279
rect 10669 42223 10725 42279
rect 10811 42223 10867 42279
rect 10953 42223 11009 42279
rect 11095 42223 11151 42279
rect 11237 42223 11293 42279
rect 11379 42223 11435 42279
rect 11521 42223 11577 42279
rect 11663 42223 11719 42279
rect 11805 42223 11861 42279
rect 11947 42223 12003 42279
rect 12089 42223 12145 42279
rect 12231 42223 12287 42279
rect 12373 42223 12429 42279
rect 12515 42223 12571 42279
rect 12657 42223 12713 42279
rect 12799 42223 12855 42279
rect 12941 42223 12997 42279
rect 13083 42223 13139 42279
rect 13225 42223 13281 42279
rect 13367 42223 13423 42279
rect 13509 42223 13565 42279
rect 13651 42223 13707 42279
rect 13793 42223 13849 42279
rect 13935 42223 13991 42279
rect 14077 42223 14133 42279
rect 14219 42223 14275 42279
rect 14361 42223 14417 42279
rect 14503 42223 14559 42279
rect 14645 42223 14701 42279
rect 14787 42223 14843 42279
rect 161 42081 217 42137
rect 303 42081 359 42137
rect 445 42081 501 42137
rect 587 42081 643 42137
rect 729 42081 785 42137
rect 871 42081 927 42137
rect 1013 42081 1069 42137
rect 1155 42081 1211 42137
rect 1297 42081 1353 42137
rect 1439 42081 1495 42137
rect 1581 42081 1637 42137
rect 1723 42081 1779 42137
rect 1865 42081 1921 42137
rect 2007 42081 2063 42137
rect 2149 42081 2205 42137
rect 2291 42081 2347 42137
rect 2433 42081 2489 42137
rect 2575 42081 2631 42137
rect 2717 42081 2773 42137
rect 2859 42081 2915 42137
rect 3001 42081 3057 42137
rect 3143 42081 3199 42137
rect 3285 42081 3341 42137
rect 3427 42081 3483 42137
rect 3569 42081 3625 42137
rect 3711 42081 3767 42137
rect 3853 42081 3909 42137
rect 3995 42081 4051 42137
rect 4137 42081 4193 42137
rect 4279 42081 4335 42137
rect 4421 42081 4477 42137
rect 4563 42081 4619 42137
rect 4705 42081 4761 42137
rect 4847 42081 4903 42137
rect 4989 42081 5045 42137
rect 5131 42081 5187 42137
rect 5273 42081 5329 42137
rect 5415 42081 5471 42137
rect 5557 42081 5613 42137
rect 5699 42081 5755 42137
rect 5841 42081 5897 42137
rect 5983 42081 6039 42137
rect 6125 42081 6181 42137
rect 6267 42081 6323 42137
rect 6409 42081 6465 42137
rect 6551 42081 6607 42137
rect 6693 42081 6749 42137
rect 6835 42081 6891 42137
rect 6977 42081 7033 42137
rect 7119 42081 7175 42137
rect 7261 42081 7317 42137
rect 7403 42081 7459 42137
rect 7545 42081 7601 42137
rect 7687 42081 7743 42137
rect 7829 42081 7885 42137
rect 7971 42081 8027 42137
rect 8113 42081 8169 42137
rect 8255 42081 8311 42137
rect 8397 42081 8453 42137
rect 8539 42081 8595 42137
rect 8681 42081 8737 42137
rect 8823 42081 8879 42137
rect 8965 42081 9021 42137
rect 9107 42081 9163 42137
rect 9249 42081 9305 42137
rect 9391 42081 9447 42137
rect 9533 42081 9589 42137
rect 9675 42081 9731 42137
rect 9817 42081 9873 42137
rect 9959 42081 10015 42137
rect 10101 42081 10157 42137
rect 10243 42081 10299 42137
rect 10385 42081 10441 42137
rect 10527 42081 10583 42137
rect 10669 42081 10725 42137
rect 10811 42081 10867 42137
rect 10953 42081 11009 42137
rect 11095 42081 11151 42137
rect 11237 42081 11293 42137
rect 11379 42081 11435 42137
rect 11521 42081 11577 42137
rect 11663 42081 11719 42137
rect 11805 42081 11861 42137
rect 11947 42081 12003 42137
rect 12089 42081 12145 42137
rect 12231 42081 12287 42137
rect 12373 42081 12429 42137
rect 12515 42081 12571 42137
rect 12657 42081 12713 42137
rect 12799 42081 12855 42137
rect 12941 42081 12997 42137
rect 13083 42081 13139 42137
rect 13225 42081 13281 42137
rect 13367 42081 13423 42137
rect 13509 42081 13565 42137
rect 13651 42081 13707 42137
rect 13793 42081 13849 42137
rect 13935 42081 13991 42137
rect 14077 42081 14133 42137
rect 14219 42081 14275 42137
rect 14361 42081 14417 42137
rect 14503 42081 14559 42137
rect 14645 42081 14701 42137
rect 14787 42081 14843 42137
rect 161 41939 217 41995
rect 303 41939 359 41995
rect 445 41939 501 41995
rect 587 41939 643 41995
rect 729 41939 785 41995
rect 871 41939 927 41995
rect 1013 41939 1069 41995
rect 1155 41939 1211 41995
rect 1297 41939 1353 41995
rect 1439 41939 1495 41995
rect 1581 41939 1637 41995
rect 1723 41939 1779 41995
rect 1865 41939 1921 41995
rect 2007 41939 2063 41995
rect 2149 41939 2205 41995
rect 2291 41939 2347 41995
rect 2433 41939 2489 41995
rect 2575 41939 2631 41995
rect 2717 41939 2773 41995
rect 2859 41939 2915 41995
rect 3001 41939 3057 41995
rect 3143 41939 3199 41995
rect 3285 41939 3341 41995
rect 3427 41939 3483 41995
rect 3569 41939 3625 41995
rect 3711 41939 3767 41995
rect 3853 41939 3909 41995
rect 3995 41939 4051 41995
rect 4137 41939 4193 41995
rect 4279 41939 4335 41995
rect 4421 41939 4477 41995
rect 4563 41939 4619 41995
rect 4705 41939 4761 41995
rect 4847 41939 4903 41995
rect 4989 41939 5045 41995
rect 5131 41939 5187 41995
rect 5273 41939 5329 41995
rect 5415 41939 5471 41995
rect 5557 41939 5613 41995
rect 5699 41939 5755 41995
rect 5841 41939 5897 41995
rect 5983 41939 6039 41995
rect 6125 41939 6181 41995
rect 6267 41939 6323 41995
rect 6409 41939 6465 41995
rect 6551 41939 6607 41995
rect 6693 41939 6749 41995
rect 6835 41939 6891 41995
rect 6977 41939 7033 41995
rect 7119 41939 7175 41995
rect 7261 41939 7317 41995
rect 7403 41939 7459 41995
rect 7545 41939 7601 41995
rect 7687 41939 7743 41995
rect 7829 41939 7885 41995
rect 7971 41939 8027 41995
rect 8113 41939 8169 41995
rect 8255 41939 8311 41995
rect 8397 41939 8453 41995
rect 8539 41939 8595 41995
rect 8681 41939 8737 41995
rect 8823 41939 8879 41995
rect 8965 41939 9021 41995
rect 9107 41939 9163 41995
rect 9249 41939 9305 41995
rect 9391 41939 9447 41995
rect 9533 41939 9589 41995
rect 9675 41939 9731 41995
rect 9817 41939 9873 41995
rect 9959 41939 10015 41995
rect 10101 41939 10157 41995
rect 10243 41939 10299 41995
rect 10385 41939 10441 41995
rect 10527 41939 10583 41995
rect 10669 41939 10725 41995
rect 10811 41939 10867 41995
rect 10953 41939 11009 41995
rect 11095 41939 11151 41995
rect 11237 41939 11293 41995
rect 11379 41939 11435 41995
rect 11521 41939 11577 41995
rect 11663 41939 11719 41995
rect 11805 41939 11861 41995
rect 11947 41939 12003 41995
rect 12089 41939 12145 41995
rect 12231 41939 12287 41995
rect 12373 41939 12429 41995
rect 12515 41939 12571 41995
rect 12657 41939 12713 41995
rect 12799 41939 12855 41995
rect 12941 41939 12997 41995
rect 13083 41939 13139 41995
rect 13225 41939 13281 41995
rect 13367 41939 13423 41995
rect 13509 41939 13565 41995
rect 13651 41939 13707 41995
rect 13793 41939 13849 41995
rect 13935 41939 13991 41995
rect 14077 41939 14133 41995
rect 14219 41939 14275 41995
rect 14361 41939 14417 41995
rect 14503 41939 14559 41995
rect 14645 41939 14701 41995
rect 14787 41939 14843 41995
rect 161 41797 217 41853
rect 303 41797 359 41853
rect 445 41797 501 41853
rect 587 41797 643 41853
rect 729 41797 785 41853
rect 871 41797 927 41853
rect 1013 41797 1069 41853
rect 1155 41797 1211 41853
rect 1297 41797 1353 41853
rect 1439 41797 1495 41853
rect 1581 41797 1637 41853
rect 1723 41797 1779 41853
rect 1865 41797 1921 41853
rect 2007 41797 2063 41853
rect 2149 41797 2205 41853
rect 2291 41797 2347 41853
rect 2433 41797 2489 41853
rect 2575 41797 2631 41853
rect 2717 41797 2773 41853
rect 2859 41797 2915 41853
rect 3001 41797 3057 41853
rect 3143 41797 3199 41853
rect 3285 41797 3341 41853
rect 3427 41797 3483 41853
rect 3569 41797 3625 41853
rect 3711 41797 3767 41853
rect 3853 41797 3909 41853
rect 3995 41797 4051 41853
rect 4137 41797 4193 41853
rect 4279 41797 4335 41853
rect 4421 41797 4477 41853
rect 4563 41797 4619 41853
rect 4705 41797 4761 41853
rect 4847 41797 4903 41853
rect 4989 41797 5045 41853
rect 5131 41797 5187 41853
rect 5273 41797 5329 41853
rect 5415 41797 5471 41853
rect 5557 41797 5613 41853
rect 5699 41797 5755 41853
rect 5841 41797 5897 41853
rect 5983 41797 6039 41853
rect 6125 41797 6181 41853
rect 6267 41797 6323 41853
rect 6409 41797 6465 41853
rect 6551 41797 6607 41853
rect 6693 41797 6749 41853
rect 6835 41797 6891 41853
rect 6977 41797 7033 41853
rect 7119 41797 7175 41853
rect 7261 41797 7317 41853
rect 7403 41797 7459 41853
rect 7545 41797 7601 41853
rect 7687 41797 7743 41853
rect 7829 41797 7885 41853
rect 7971 41797 8027 41853
rect 8113 41797 8169 41853
rect 8255 41797 8311 41853
rect 8397 41797 8453 41853
rect 8539 41797 8595 41853
rect 8681 41797 8737 41853
rect 8823 41797 8879 41853
rect 8965 41797 9021 41853
rect 9107 41797 9163 41853
rect 9249 41797 9305 41853
rect 9391 41797 9447 41853
rect 9533 41797 9589 41853
rect 9675 41797 9731 41853
rect 9817 41797 9873 41853
rect 9959 41797 10015 41853
rect 10101 41797 10157 41853
rect 10243 41797 10299 41853
rect 10385 41797 10441 41853
rect 10527 41797 10583 41853
rect 10669 41797 10725 41853
rect 10811 41797 10867 41853
rect 10953 41797 11009 41853
rect 11095 41797 11151 41853
rect 11237 41797 11293 41853
rect 11379 41797 11435 41853
rect 11521 41797 11577 41853
rect 11663 41797 11719 41853
rect 11805 41797 11861 41853
rect 11947 41797 12003 41853
rect 12089 41797 12145 41853
rect 12231 41797 12287 41853
rect 12373 41797 12429 41853
rect 12515 41797 12571 41853
rect 12657 41797 12713 41853
rect 12799 41797 12855 41853
rect 12941 41797 12997 41853
rect 13083 41797 13139 41853
rect 13225 41797 13281 41853
rect 13367 41797 13423 41853
rect 13509 41797 13565 41853
rect 13651 41797 13707 41853
rect 13793 41797 13849 41853
rect 13935 41797 13991 41853
rect 14077 41797 14133 41853
rect 14219 41797 14275 41853
rect 14361 41797 14417 41853
rect 14503 41797 14559 41853
rect 14645 41797 14701 41853
rect 14787 41797 14843 41853
rect 161 41655 217 41711
rect 303 41655 359 41711
rect 445 41655 501 41711
rect 587 41655 643 41711
rect 729 41655 785 41711
rect 871 41655 927 41711
rect 1013 41655 1069 41711
rect 1155 41655 1211 41711
rect 1297 41655 1353 41711
rect 1439 41655 1495 41711
rect 1581 41655 1637 41711
rect 1723 41655 1779 41711
rect 1865 41655 1921 41711
rect 2007 41655 2063 41711
rect 2149 41655 2205 41711
rect 2291 41655 2347 41711
rect 2433 41655 2489 41711
rect 2575 41655 2631 41711
rect 2717 41655 2773 41711
rect 2859 41655 2915 41711
rect 3001 41655 3057 41711
rect 3143 41655 3199 41711
rect 3285 41655 3341 41711
rect 3427 41655 3483 41711
rect 3569 41655 3625 41711
rect 3711 41655 3767 41711
rect 3853 41655 3909 41711
rect 3995 41655 4051 41711
rect 4137 41655 4193 41711
rect 4279 41655 4335 41711
rect 4421 41655 4477 41711
rect 4563 41655 4619 41711
rect 4705 41655 4761 41711
rect 4847 41655 4903 41711
rect 4989 41655 5045 41711
rect 5131 41655 5187 41711
rect 5273 41655 5329 41711
rect 5415 41655 5471 41711
rect 5557 41655 5613 41711
rect 5699 41655 5755 41711
rect 5841 41655 5897 41711
rect 5983 41655 6039 41711
rect 6125 41655 6181 41711
rect 6267 41655 6323 41711
rect 6409 41655 6465 41711
rect 6551 41655 6607 41711
rect 6693 41655 6749 41711
rect 6835 41655 6891 41711
rect 6977 41655 7033 41711
rect 7119 41655 7175 41711
rect 7261 41655 7317 41711
rect 7403 41655 7459 41711
rect 7545 41655 7601 41711
rect 7687 41655 7743 41711
rect 7829 41655 7885 41711
rect 7971 41655 8027 41711
rect 8113 41655 8169 41711
rect 8255 41655 8311 41711
rect 8397 41655 8453 41711
rect 8539 41655 8595 41711
rect 8681 41655 8737 41711
rect 8823 41655 8879 41711
rect 8965 41655 9021 41711
rect 9107 41655 9163 41711
rect 9249 41655 9305 41711
rect 9391 41655 9447 41711
rect 9533 41655 9589 41711
rect 9675 41655 9731 41711
rect 9817 41655 9873 41711
rect 9959 41655 10015 41711
rect 10101 41655 10157 41711
rect 10243 41655 10299 41711
rect 10385 41655 10441 41711
rect 10527 41655 10583 41711
rect 10669 41655 10725 41711
rect 10811 41655 10867 41711
rect 10953 41655 11009 41711
rect 11095 41655 11151 41711
rect 11237 41655 11293 41711
rect 11379 41655 11435 41711
rect 11521 41655 11577 41711
rect 11663 41655 11719 41711
rect 11805 41655 11861 41711
rect 11947 41655 12003 41711
rect 12089 41655 12145 41711
rect 12231 41655 12287 41711
rect 12373 41655 12429 41711
rect 12515 41655 12571 41711
rect 12657 41655 12713 41711
rect 12799 41655 12855 41711
rect 12941 41655 12997 41711
rect 13083 41655 13139 41711
rect 13225 41655 13281 41711
rect 13367 41655 13423 41711
rect 13509 41655 13565 41711
rect 13651 41655 13707 41711
rect 13793 41655 13849 41711
rect 13935 41655 13991 41711
rect 14077 41655 14133 41711
rect 14219 41655 14275 41711
rect 14361 41655 14417 41711
rect 14503 41655 14559 41711
rect 14645 41655 14701 41711
rect 14787 41655 14843 41711
rect 161 41513 217 41569
rect 303 41513 359 41569
rect 445 41513 501 41569
rect 587 41513 643 41569
rect 729 41513 785 41569
rect 871 41513 927 41569
rect 1013 41513 1069 41569
rect 1155 41513 1211 41569
rect 1297 41513 1353 41569
rect 1439 41513 1495 41569
rect 1581 41513 1637 41569
rect 1723 41513 1779 41569
rect 1865 41513 1921 41569
rect 2007 41513 2063 41569
rect 2149 41513 2205 41569
rect 2291 41513 2347 41569
rect 2433 41513 2489 41569
rect 2575 41513 2631 41569
rect 2717 41513 2773 41569
rect 2859 41513 2915 41569
rect 3001 41513 3057 41569
rect 3143 41513 3199 41569
rect 3285 41513 3341 41569
rect 3427 41513 3483 41569
rect 3569 41513 3625 41569
rect 3711 41513 3767 41569
rect 3853 41513 3909 41569
rect 3995 41513 4051 41569
rect 4137 41513 4193 41569
rect 4279 41513 4335 41569
rect 4421 41513 4477 41569
rect 4563 41513 4619 41569
rect 4705 41513 4761 41569
rect 4847 41513 4903 41569
rect 4989 41513 5045 41569
rect 5131 41513 5187 41569
rect 5273 41513 5329 41569
rect 5415 41513 5471 41569
rect 5557 41513 5613 41569
rect 5699 41513 5755 41569
rect 5841 41513 5897 41569
rect 5983 41513 6039 41569
rect 6125 41513 6181 41569
rect 6267 41513 6323 41569
rect 6409 41513 6465 41569
rect 6551 41513 6607 41569
rect 6693 41513 6749 41569
rect 6835 41513 6891 41569
rect 6977 41513 7033 41569
rect 7119 41513 7175 41569
rect 7261 41513 7317 41569
rect 7403 41513 7459 41569
rect 7545 41513 7601 41569
rect 7687 41513 7743 41569
rect 7829 41513 7885 41569
rect 7971 41513 8027 41569
rect 8113 41513 8169 41569
rect 8255 41513 8311 41569
rect 8397 41513 8453 41569
rect 8539 41513 8595 41569
rect 8681 41513 8737 41569
rect 8823 41513 8879 41569
rect 8965 41513 9021 41569
rect 9107 41513 9163 41569
rect 9249 41513 9305 41569
rect 9391 41513 9447 41569
rect 9533 41513 9589 41569
rect 9675 41513 9731 41569
rect 9817 41513 9873 41569
rect 9959 41513 10015 41569
rect 10101 41513 10157 41569
rect 10243 41513 10299 41569
rect 10385 41513 10441 41569
rect 10527 41513 10583 41569
rect 10669 41513 10725 41569
rect 10811 41513 10867 41569
rect 10953 41513 11009 41569
rect 11095 41513 11151 41569
rect 11237 41513 11293 41569
rect 11379 41513 11435 41569
rect 11521 41513 11577 41569
rect 11663 41513 11719 41569
rect 11805 41513 11861 41569
rect 11947 41513 12003 41569
rect 12089 41513 12145 41569
rect 12231 41513 12287 41569
rect 12373 41513 12429 41569
rect 12515 41513 12571 41569
rect 12657 41513 12713 41569
rect 12799 41513 12855 41569
rect 12941 41513 12997 41569
rect 13083 41513 13139 41569
rect 13225 41513 13281 41569
rect 13367 41513 13423 41569
rect 13509 41513 13565 41569
rect 13651 41513 13707 41569
rect 13793 41513 13849 41569
rect 13935 41513 13991 41569
rect 14077 41513 14133 41569
rect 14219 41513 14275 41569
rect 14361 41513 14417 41569
rect 14503 41513 14559 41569
rect 14645 41513 14701 41569
rect 14787 41513 14843 41569
rect 161 41371 217 41427
rect 303 41371 359 41427
rect 445 41371 501 41427
rect 587 41371 643 41427
rect 729 41371 785 41427
rect 871 41371 927 41427
rect 1013 41371 1069 41427
rect 1155 41371 1211 41427
rect 1297 41371 1353 41427
rect 1439 41371 1495 41427
rect 1581 41371 1637 41427
rect 1723 41371 1779 41427
rect 1865 41371 1921 41427
rect 2007 41371 2063 41427
rect 2149 41371 2205 41427
rect 2291 41371 2347 41427
rect 2433 41371 2489 41427
rect 2575 41371 2631 41427
rect 2717 41371 2773 41427
rect 2859 41371 2915 41427
rect 3001 41371 3057 41427
rect 3143 41371 3199 41427
rect 3285 41371 3341 41427
rect 3427 41371 3483 41427
rect 3569 41371 3625 41427
rect 3711 41371 3767 41427
rect 3853 41371 3909 41427
rect 3995 41371 4051 41427
rect 4137 41371 4193 41427
rect 4279 41371 4335 41427
rect 4421 41371 4477 41427
rect 4563 41371 4619 41427
rect 4705 41371 4761 41427
rect 4847 41371 4903 41427
rect 4989 41371 5045 41427
rect 5131 41371 5187 41427
rect 5273 41371 5329 41427
rect 5415 41371 5471 41427
rect 5557 41371 5613 41427
rect 5699 41371 5755 41427
rect 5841 41371 5897 41427
rect 5983 41371 6039 41427
rect 6125 41371 6181 41427
rect 6267 41371 6323 41427
rect 6409 41371 6465 41427
rect 6551 41371 6607 41427
rect 6693 41371 6749 41427
rect 6835 41371 6891 41427
rect 6977 41371 7033 41427
rect 7119 41371 7175 41427
rect 7261 41371 7317 41427
rect 7403 41371 7459 41427
rect 7545 41371 7601 41427
rect 7687 41371 7743 41427
rect 7829 41371 7885 41427
rect 7971 41371 8027 41427
rect 8113 41371 8169 41427
rect 8255 41371 8311 41427
rect 8397 41371 8453 41427
rect 8539 41371 8595 41427
rect 8681 41371 8737 41427
rect 8823 41371 8879 41427
rect 8965 41371 9021 41427
rect 9107 41371 9163 41427
rect 9249 41371 9305 41427
rect 9391 41371 9447 41427
rect 9533 41371 9589 41427
rect 9675 41371 9731 41427
rect 9817 41371 9873 41427
rect 9959 41371 10015 41427
rect 10101 41371 10157 41427
rect 10243 41371 10299 41427
rect 10385 41371 10441 41427
rect 10527 41371 10583 41427
rect 10669 41371 10725 41427
rect 10811 41371 10867 41427
rect 10953 41371 11009 41427
rect 11095 41371 11151 41427
rect 11237 41371 11293 41427
rect 11379 41371 11435 41427
rect 11521 41371 11577 41427
rect 11663 41371 11719 41427
rect 11805 41371 11861 41427
rect 11947 41371 12003 41427
rect 12089 41371 12145 41427
rect 12231 41371 12287 41427
rect 12373 41371 12429 41427
rect 12515 41371 12571 41427
rect 12657 41371 12713 41427
rect 12799 41371 12855 41427
rect 12941 41371 12997 41427
rect 13083 41371 13139 41427
rect 13225 41371 13281 41427
rect 13367 41371 13423 41427
rect 13509 41371 13565 41427
rect 13651 41371 13707 41427
rect 13793 41371 13849 41427
rect 13935 41371 13991 41427
rect 14077 41371 14133 41427
rect 14219 41371 14275 41427
rect 14361 41371 14417 41427
rect 14503 41371 14559 41427
rect 14645 41371 14701 41427
rect 14787 41371 14843 41427
rect 161 41229 217 41285
rect 303 41229 359 41285
rect 445 41229 501 41285
rect 587 41229 643 41285
rect 729 41229 785 41285
rect 871 41229 927 41285
rect 1013 41229 1069 41285
rect 1155 41229 1211 41285
rect 1297 41229 1353 41285
rect 1439 41229 1495 41285
rect 1581 41229 1637 41285
rect 1723 41229 1779 41285
rect 1865 41229 1921 41285
rect 2007 41229 2063 41285
rect 2149 41229 2205 41285
rect 2291 41229 2347 41285
rect 2433 41229 2489 41285
rect 2575 41229 2631 41285
rect 2717 41229 2773 41285
rect 2859 41229 2915 41285
rect 3001 41229 3057 41285
rect 3143 41229 3199 41285
rect 3285 41229 3341 41285
rect 3427 41229 3483 41285
rect 3569 41229 3625 41285
rect 3711 41229 3767 41285
rect 3853 41229 3909 41285
rect 3995 41229 4051 41285
rect 4137 41229 4193 41285
rect 4279 41229 4335 41285
rect 4421 41229 4477 41285
rect 4563 41229 4619 41285
rect 4705 41229 4761 41285
rect 4847 41229 4903 41285
rect 4989 41229 5045 41285
rect 5131 41229 5187 41285
rect 5273 41229 5329 41285
rect 5415 41229 5471 41285
rect 5557 41229 5613 41285
rect 5699 41229 5755 41285
rect 5841 41229 5897 41285
rect 5983 41229 6039 41285
rect 6125 41229 6181 41285
rect 6267 41229 6323 41285
rect 6409 41229 6465 41285
rect 6551 41229 6607 41285
rect 6693 41229 6749 41285
rect 6835 41229 6891 41285
rect 6977 41229 7033 41285
rect 7119 41229 7175 41285
rect 7261 41229 7317 41285
rect 7403 41229 7459 41285
rect 7545 41229 7601 41285
rect 7687 41229 7743 41285
rect 7829 41229 7885 41285
rect 7971 41229 8027 41285
rect 8113 41229 8169 41285
rect 8255 41229 8311 41285
rect 8397 41229 8453 41285
rect 8539 41229 8595 41285
rect 8681 41229 8737 41285
rect 8823 41229 8879 41285
rect 8965 41229 9021 41285
rect 9107 41229 9163 41285
rect 9249 41229 9305 41285
rect 9391 41229 9447 41285
rect 9533 41229 9589 41285
rect 9675 41229 9731 41285
rect 9817 41229 9873 41285
rect 9959 41229 10015 41285
rect 10101 41229 10157 41285
rect 10243 41229 10299 41285
rect 10385 41229 10441 41285
rect 10527 41229 10583 41285
rect 10669 41229 10725 41285
rect 10811 41229 10867 41285
rect 10953 41229 11009 41285
rect 11095 41229 11151 41285
rect 11237 41229 11293 41285
rect 11379 41229 11435 41285
rect 11521 41229 11577 41285
rect 11663 41229 11719 41285
rect 11805 41229 11861 41285
rect 11947 41229 12003 41285
rect 12089 41229 12145 41285
rect 12231 41229 12287 41285
rect 12373 41229 12429 41285
rect 12515 41229 12571 41285
rect 12657 41229 12713 41285
rect 12799 41229 12855 41285
rect 12941 41229 12997 41285
rect 13083 41229 13139 41285
rect 13225 41229 13281 41285
rect 13367 41229 13423 41285
rect 13509 41229 13565 41285
rect 13651 41229 13707 41285
rect 13793 41229 13849 41285
rect 13935 41229 13991 41285
rect 14077 41229 14133 41285
rect 14219 41229 14275 41285
rect 14361 41229 14417 41285
rect 14503 41229 14559 41285
rect 14645 41229 14701 41285
rect 14787 41229 14843 41285
rect 161 40907 217 40963
rect 303 40907 359 40963
rect 445 40907 501 40963
rect 587 40907 643 40963
rect 729 40907 785 40963
rect 871 40907 927 40963
rect 1013 40907 1069 40963
rect 1155 40907 1211 40963
rect 1297 40907 1353 40963
rect 1439 40907 1495 40963
rect 1581 40907 1637 40963
rect 1723 40907 1779 40963
rect 1865 40907 1921 40963
rect 2007 40907 2063 40963
rect 2149 40907 2205 40963
rect 2291 40907 2347 40963
rect 2433 40907 2489 40963
rect 2575 40907 2631 40963
rect 2717 40907 2773 40963
rect 2859 40907 2915 40963
rect 3001 40907 3057 40963
rect 3143 40907 3199 40963
rect 3285 40907 3341 40963
rect 3427 40907 3483 40963
rect 3569 40907 3625 40963
rect 3711 40907 3767 40963
rect 3853 40907 3909 40963
rect 3995 40907 4051 40963
rect 4137 40907 4193 40963
rect 4279 40907 4335 40963
rect 4421 40907 4477 40963
rect 4563 40907 4619 40963
rect 4705 40907 4761 40963
rect 4847 40907 4903 40963
rect 4989 40907 5045 40963
rect 5131 40907 5187 40963
rect 5273 40907 5329 40963
rect 5415 40907 5471 40963
rect 5557 40907 5613 40963
rect 5699 40907 5755 40963
rect 5841 40907 5897 40963
rect 5983 40907 6039 40963
rect 6125 40907 6181 40963
rect 6267 40907 6323 40963
rect 6409 40907 6465 40963
rect 6551 40907 6607 40963
rect 6693 40907 6749 40963
rect 6835 40907 6891 40963
rect 6977 40907 7033 40963
rect 7119 40907 7175 40963
rect 7261 40907 7317 40963
rect 7403 40907 7459 40963
rect 7545 40907 7601 40963
rect 7687 40907 7743 40963
rect 7829 40907 7885 40963
rect 7971 40907 8027 40963
rect 8113 40907 8169 40963
rect 8255 40907 8311 40963
rect 8397 40907 8453 40963
rect 8539 40907 8595 40963
rect 8681 40907 8737 40963
rect 8823 40907 8879 40963
rect 8965 40907 9021 40963
rect 9107 40907 9163 40963
rect 9249 40907 9305 40963
rect 9391 40907 9447 40963
rect 9533 40907 9589 40963
rect 9675 40907 9731 40963
rect 9817 40907 9873 40963
rect 9959 40907 10015 40963
rect 10101 40907 10157 40963
rect 10243 40907 10299 40963
rect 10385 40907 10441 40963
rect 10527 40907 10583 40963
rect 10669 40907 10725 40963
rect 10811 40907 10867 40963
rect 10953 40907 11009 40963
rect 11095 40907 11151 40963
rect 11237 40907 11293 40963
rect 11379 40907 11435 40963
rect 11521 40907 11577 40963
rect 11663 40907 11719 40963
rect 11805 40907 11861 40963
rect 11947 40907 12003 40963
rect 12089 40907 12145 40963
rect 12231 40907 12287 40963
rect 12373 40907 12429 40963
rect 12515 40907 12571 40963
rect 12657 40907 12713 40963
rect 12799 40907 12855 40963
rect 12941 40907 12997 40963
rect 13083 40907 13139 40963
rect 13225 40907 13281 40963
rect 13367 40907 13423 40963
rect 13509 40907 13565 40963
rect 13651 40907 13707 40963
rect 13793 40907 13849 40963
rect 13935 40907 13991 40963
rect 14077 40907 14133 40963
rect 14219 40907 14275 40963
rect 14361 40907 14417 40963
rect 14503 40907 14559 40963
rect 14645 40907 14701 40963
rect 14787 40907 14843 40963
rect 161 40765 217 40821
rect 303 40765 359 40821
rect 445 40765 501 40821
rect 587 40765 643 40821
rect 729 40765 785 40821
rect 871 40765 927 40821
rect 1013 40765 1069 40821
rect 1155 40765 1211 40821
rect 1297 40765 1353 40821
rect 1439 40765 1495 40821
rect 1581 40765 1637 40821
rect 1723 40765 1779 40821
rect 1865 40765 1921 40821
rect 2007 40765 2063 40821
rect 2149 40765 2205 40821
rect 2291 40765 2347 40821
rect 2433 40765 2489 40821
rect 2575 40765 2631 40821
rect 2717 40765 2773 40821
rect 2859 40765 2915 40821
rect 3001 40765 3057 40821
rect 3143 40765 3199 40821
rect 3285 40765 3341 40821
rect 3427 40765 3483 40821
rect 3569 40765 3625 40821
rect 3711 40765 3767 40821
rect 3853 40765 3909 40821
rect 3995 40765 4051 40821
rect 4137 40765 4193 40821
rect 4279 40765 4335 40821
rect 4421 40765 4477 40821
rect 4563 40765 4619 40821
rect 4705 40765 4761 40821
rect 4847 40765 4903 40821
rect 4989 40765 5045 40821
rect 5131 40765 5187 40821
rect 5273 40765 5329 40821
rect 5415 40765 5471 40821
rect 5557 40765 5613 40821
rect 5699 40765 5755 40821
rect 5841 40765 5897 40821
rect 5983 40765 6039 40821
rect 6125 40765 6181 40821
rect 6267 40765 6323 40821
rect 6409 40765 6465 40821
rect 6551 40765 6607 40821
rect 6693 40765 6749 40821
rect 6835 40765 6891 40821
rect 6977 40765 7033 40821
rect 7119 40765 7175 40821
rect 7261 40765 7317 40821
rect 7403 40765 7459 40821
rect 7545 40765 7601 40821
rect 7687 40765 7743 40821
rect 7829 40765 7885 40821
rect 7971 40765 8027 40821
rect 8113 40765 8169 40821
rect 8255 40765 8311 40821
rect 8397 40765 8453 40821
rect 8539 40765 8595 40821
rect 8681 40765 8737 40821
rect 8823 40765 8879 40821
rect 8965 40765 9021 40821
rect 9107 40765 9163 40821
rect 9249 40765 9305 40821
rect 9391 40765 9447 40821
rect 9533 40765 9589 40821
rect 9675 40765 9731 40821
rect 9817 40765 9873 40821
rect 9959 40765 10015 40821
rect 10101 40765 10157 40821
rect 10243 40765 10299 40821
rect 10385 40765 10441 40821
rect 10527 40765 10583 40821
rect 10669 40765 10725 40821
rect 10811 40765 10867 40821
rect 10953 40765 11009 40821
rect 11095 40765 11151 40821
rect 11237 40765 11293 40821
rect 11379 40765 11435 40821
rect 11521 40765 11577 40821
rect 11663 40765 11719 40821
rect 11805 40765 11861 40821
rect 11947 40765 12003 40821
rect 12089 40765 12145 40821
rect 12231 40765 12287 40821
rect 12373 40765 12429 40821
rect 12515 40765 12571 40821
rect 12657 40765 12713 40821
rect 12799 40765 12855 40821
rect 12941 40765 12997 40821
rect 13083 40765 13139 40821
rect 13225 40765 13281 40821
rect 13367 40765 13423 40821
rect 13509 40765 13565 40821
rect 13651 40765 13707 40821
rect 13793 40765 13849 40821
rect 13935 40765 13991 40821
rect 14077 40765 14133 40821
rect 14219 40765 14275 40821
rect 14361 40765 14417 40821
rect 14503 40765 14559 40821
rect 14645 40765 14701 40821
rect 14787 40765 14843 40821
rect 161 40623 217 40679
rect 303 40623 359 40679
rect 445 40623 501 40679
rect 587 40623 643 40679
rect 729 40623 785 40679
rect 871 40623 927 40679
rect 1013 40623 1069 40679
rect 1155 40623 1211 40679
rect 1297 40623 1353 40679
rect 1439 40623 1495 40679
rect 1581 40623 1637 40679
rect 1723 40623 1779 40679
rect 1865 40623 1921 40679
rect 2007 40623 2063 40679
rect 2149 40623 2205 40679
rect 2291 40623 2347 40679
rect 2433 40623 2489 40679
rect 2575 40623 2631 40679
rect 2717 40623 2773 40679
rect 2859 40623 2915 40679
rect 3001 40623 3057 40679
rect 3143 40623 3199 40679
rect 3285 40623 3341 40679
rect 3427 40623 3483 40679
rect 3569 40623 3625 40679
rect 3711 40623 3767 40679
rect 3853 40623 3909 40679
rect 3995 40623 4051 40679
rect 4137 40623 4193 40679
rect 4279 40623 4335 40679
rect 4421 40623 4477 40679
rect 4563 40623 4619 40679
rect 4705 40623 4761 40679
rect 4847 40623 4903 40679
rect 4989 40623 5045 40679
rect 5131 40623 5187 40679
rect 5273 40623 5329 40679
rect 5415 40623 5471 40679
rect 5557 40623 5613 40679
rect 5699 40623 5755 40679
rect 5841 40623 5897 40679
rect 5983 40623 6039 40679
rect 6125 40623 6181 40679
rect 6267 40623 6323 40679
rect 6409 40623 6465 40679
rect 6551 40623 6607 40679
rect 6693 40623 6749 40679
rect 6835 40623 6891 40679
rect 6977 40623 7033 40679
rect 7119 40623 7175 40679
rect 7261 40623 7317 40679
rect 7403 40623 7459 40679
rect 7545 40623 7601 40679
rect 7687 40623 7743 40679
rect 7829 40623 7885 40679
rect 7971 40623 8027 40679
rect 8113 40623 8169 40679
rect 8255 40623 8311 40679
rect 8397 40623 8453 40679
rect 8539 40623 8595 40679
rect 8681 40623 8737 40679
rect 8823 40623 8879 40679
rect 8965 40623 9021 40679
rect 9107 40623 9163 40679
rect 9249 40623 9305 40679
rect 9391 40623 9447 40679
rect 9533 40623 9589 40679
rect 9675 40623 9731 40679
rect 9817 40623 9873 40679
rect 9959 40623 10015 40679
rect 10101 40623 10157 40679
rect 10243 40623 10299 40679
rect 10385 40623 10441 40679
rect 10527 40623 10583 40679
rect 10669 40623 10725 40679
rect 10811 40623 10867 40679
rect 10953 40623 11009 40679
rect 11095 40623 11151 40679
rect 11237 40623 11293 40679
rect 11379 40623 11435 40679
rect 11521 40623 11577 40679
rect 11663 40623 11719 40679
rect 11805 40623 11861 40679
rect 11947 40623 12003 40679
rect 12089 40623 12145 40679
rect 12231 40623 12287 40679
rect 12373 40623 12429 40679
rect 12515 40623 12571 40679
rect 12657 40623 12713 40679
rect 12799 40623 12855 40679
rect 12941 40623 12997 40679
rect 13083 40623 13139 40679
rect 13225 40623 13281 40679
rect 13367 40623 13423 40679
rect 13509 40623 13565 40679
rect 13651 40623 13707 40679
rect 13793 40623 13849 40679
rect 13935 40623 13991 40679
rect 14077 40623 14133 40679
rect 14219 40623 14275 40679
rect 14361 40623 14417 40679
rect 14503 40623 14559 40679
rect 14645 40623 14701 40679
rect 14787 40623 14843 40679
rect 161 40481 217 40537
rect 303 40481 359 40537
rect 445 40481 501 40537
rect 587 40481 643 40537
rect 729 40481 785 40537
rect 871 40481 927 40537
rect 1013 40481 1069 40537
rect 1155 40481 1211 40537
rect 1297 40481 1353 40537
rect 1439 40481 1495 40537
rect 1581 40481 1637 40537
rect 1723 40481 1779 40537
rect 1865 40481 1921 40537
rect 2007 40481 2063 40537
rect 2149 40481 2205 40537
rect 2291 40481 2347 40537
rect 2433 40481 2489 40537
rect 2575 40481 2631 40537
rect 2717 40481 2773 40537
rect 2859 40481 2915 40537
rect 3001 40481 3057 40537
rect 3143 40481 3199 40537
rect 3285 40481 3341 40537
rect 3427 40481 3483 40537
rect 3569 40481 3625 40537
rect 3711 40481 3767 40537
rect 3853 40481 3909 40537
rect 3995 40481 4051 40537
rect 4137 40481 4193 40537
rect 4279 40481 4335 40537
rect 4421 40481 4477 40537
rect 4563 40481 4619 40537
rect 4705 40481 4761 40537
rect 4847 40481 4903 40537
rect 4989 40481 5045 40537
rect 5131 40481 5187 40537
rect 5273 40481 5329 40537
rect 5415 40481 5471 40537
rect 5557 40481 5613 40537
rect 5699 40481 5755 40537
rect 5841 40481 5897 40537
rect 5983 40481 6039 40537
rect 6125 40481 6181 40537
rect 6267 40481 6323 40537
rect 6409 40481 6465 40537
rect 6551 40481 6607 40537
rect 6693 40481 6749 40537
rect 6835 40481 6891 40537
rect 6977 40481 7033 40537
rect 7119 40481 7175 40537
rect 7261 40481 7317 40537
rect 7403 40481 7459 40537
rect 7545 40481 7601 40537
rect 7687 40481 7743 40537
rect 7829 40481 7885 40537
rect 7971 40481 8027 40537
rect 8113 40481 8169 40537
rect 8255 40481 8311 40537
rect 8397 40481 8453 40537
rect 8539 40481 8595 40537
rect 8681 40481 8737 40537
rect 8823 40481 8879 40537
rect 8965 40481 9021 40537
rect 9107 40481 9163 40537
rect 9249 40481 9305 40537
rect 9391 40481 9447 40537
rect 9533 40481 9589 40537
rect 9675 40481 9731 40537
rect 9817 40481 9873 40537
rect 9959 40481 10015 40537
rect 10101 40481 10157 40537
rect 10243 40481 10299 40537
rect 10385 40481 10441 40537
rect 10527 40481 10583 40537
rect 10669 40481 10725 40537
rect 10811 40481 10867 40537
rect 10953 40481 11009 40537
rect 11095 40481 11151 40537
rect 11237 40481 11293 40537
rect 11379 40481 11435 40537
rect 11521 40481 11577 40537
rect 11663 40481 11719 40537
rect 11805 40481 11861 40537
rect 11947 40481 12003 40537
rect 12089 40481 12145 40537
rect 12231 40481 12287 40537
rect 12373 40481 12429 40537
rect 12515 40481 12571 40537
rect 12657 40481 12713 40537
rect 12799 40481 12855 40537
rect 12941 40481 12997 40537
rect 13083 40481 13139 40537
rect 13225 40481 13281 40537
rect 13367 40481 13423 40537
rect 13509 40481 13565 40537
rect 13651 40481 13707 40537
rect 13793 40481 13849 40537
rect 13935 40481 13991 40537
rect 14077 40481 14133 40537
rect 14219 40481 14275 40537
rect 14361 40481 14417 40537
rect 14503 40481 14559 40537
rect 14645 40481 14701 40537
rect 14787 40481 14843 40537
rect 161 40339 217 40395
rect 303 40339 359 40395
rect 445 40339 501 40395
rect 587 40339 643 40395
rect 729 40339 785 40395
rect 871 40339 927 40395
rect 1013 40339 1069 40395
rect 1155 40339 1211 40395
rect 1297 40339 1353 40395
rect 1439 40339 1495 40395
rect 1581 40339 1637 40395
rect 1723 40339 1779 40395
rect 1865 40339 1921 40395
rect 2007 40339 2063 40395
rect 2149 40339 2205 40395
rect 2291 40339 2347 40395
rect 2433 40339 2489 40395
rect 2575 40339 2631 40395
rect 2717 40339 2773 40395
rect 2859 40339 2915 40395
rect 3001 40339 3057 40395
rect 3143 40339 3199 40395
rect 3285 40339 3341 40395
rect 3427 40339 3483 40395
rect 3569 40339 3625 40395
rect 3711 40339 3767 40395
rect 3853 40339 3909 40395
rect 3995 40339 4051 40395
rect 4137 40339 4193 40395
rect 4279 40339 4335 40395
rect 4421 40339 4477 40395
rect 4563 40339 4619 40395
rect 4705 40339 4761 40395
rect 4847 40339 4903 40395
rect 4989 40339 5045 40395
rect 5131 40339 5187 40395
rect 5273 40339 5329 40395
rect 5415 40339 5471 40395
rect 5557 40339 5613 40395
rect 5699 40339 5755 40395
rect 5841 40339 5897 40395
rect 5983 40339 6039 40395
rect 6125 40339 6181 40395
rect 6267 40339 6323 40395
rect 6409 40339 6465 40395
rect 6551 40339 6607 40395
rect 6693 40339 6749 40395
rect 6835 40339 6891 40395
rect 6977 40339 7033 40395
rect 7119 40339 7175 40395
rect 7261 40339 7317 40395
rect 7403 40339 7459 40395
rect 7545 40339 7601 40395
rect 7687 40339 7743 40395
rect 7829 40339 7885 40395
rect 7971 40339 8027 40395
rect 8113 40339 8169 40395
rect 8255 40339 8311 40395
rect 8397 40339 8453 40395
rect 8539 40339 8595 40395
rect 8681 40339 8737 40395
rect 8823 40339 8879 40395
rect 8965 40339 9021 40395
rect 9107 40339 9163 40395
rect 9249 40339 9305 40395
rect 9391 40339 9447 40395
rect 9533 40339 9589 40395
rect 9675 40339 9731 40395
rect 9817 40339 9873 40395
rect 9959 40339 10015 40395
rect 10101 40339 10157 40395
rect 10243 40339 10299 40395
rect 10385 40339 10441 40395
rect 10527 40339 10583 40395
rect 10669 40339 10725 40395
rect 10811 40339 10867 40395
rect 10953 40339 11009 40395
rect 11095 40339 11151 40395
rect 11237 40339 11293 40395
rect 11379 40339 11435 40395
rect 11521 40339 11577 40395
rect 11663 40339 11719 40395
rect 11805 40339 11861 40395
rect 11947 40339 12003 40395
rect 12089 40339 12145 40395
rect 12231 40339 12287 40395
rect 12373 40339 12429 40395
rect 12515 40339 12571 40395
rect 12657 40339 12713 40395
rect 12799 40339 12855 40395
rect 12941 40339 12997 40395
rect 13083 40339 13139 40395
rect 13225 40339 13281 40395
rect 13367 40339 13423 40395
rect 13509 40339 13565 40395
rect 13651 40339 13707 40395
rect 13793 40339 13849 40395
rect 13935 40339 13991 40395
rect 14077 40339 14133 40395
rect 14219 40339 14275 40395
rect 14361 40339 14417 40395
rect 14503 40339 14559 40395
rect 14645 40339 14701 40395
rect 14787 40339 14843 40395
rect 161 40197 217 40253
rect 303 40197 359 40253
rect 445 40197 501 40253
rect 587 40197 643 40253
rect 729 40197 785 40253
rect 871 40197 927 40253
rect 1013 40197 1069 40253
rect 1155 40197 1211 40253
rect 1297 40197 1353 40253
rect 1439 40197 1495 40253
rect 1581 40197 1637 40253
rect 1723 40197 1779 40253
rect 1865 40197 1921 40253
rect 2007 40197 2063 40253
rect 2149 40197 2205 40253
rect 2291 40197 2347 40253
rect 2433 40197 2489 40253
rect 2575 40197 2631 40253
rect 2717 40197 2773 40253
rect 2859 40197 2915 40253
rect 3001 40197 3057 40253
rect 3143 40197 3199 40253
rect 3285 40197 3341 40253
rect 3427 40197 3483 40253
rect 3569 40197 3625 40253
rect 3711 40197 3767 40253
rect 3853 40197 3909 40253
rect 3995 40197 4051 40253
rect 4137 40197 4193 40253
rect 4279 40197 4335 40253
rect 4421 40197 4477 40253
rect 4563 40197 4619 40253
rect 4705 40197 4761 40253
rect 4847 40197 4903 40253
rect 4989 40197 5045 40253
rect 5131 40197 5187 40253
rect 5273 40197 5329 40253
rect 5415 40197 5471 40253
rect 5557 40197 5613 40253
rect 5699 40197 5755 40253
rect 5841 40197 5897 40253
rect 5983 40197 6039 40253
rect 6125 40197 6181 40253
rect 6267 40197 6323 40253
rect 6409 40197 6465 40253
rect 6551 40197 6607 40253
rect 6693 40197 6749 40253
rect 6835 40197 6891 40253
rect 6977 40197 7033 40253
rect 7119 40197 7175 40253
rect 7261 40197 7317 40253
rect 7403 40197 7459 40253
rect 7545 40197 7601 40253
rect 7687 40197 7743 40253
rect 7829 40197 7885 40253
rect 7971 40197 8027 40253
rect 8113 40197 8169 40253
rect 8255 40197 8311 40253
rect 8397 40197 8453 40253
rect 8539 40197 8595 40253
rect 8681 40197 8737 40253
rect 8823 40197 8879 40253
rect 8965 40197 9021 40253
rect 9107 40197 9163 40253
rect 9249 40197 9305 40253
rect 9391 40197 9447 40253
rect 9533 40197 9589 40253
rect 9675 40197 9731 40253
rect 9817 40197 9873 40253
rect 9959 40197 10015 40253
rect 10101 40197 10157 40253
rect 10243 40197 10299 40253
rect 10385 40197 10441 40253
rect 10527 40197 10583 40253
rect 10669 40197 10725 40253
rect 10811 40197 10867 40253
rect 10953 40197 11009 40253
rect 11095 40197 11151 40253
rect 11237 40197 11293 40253
rect 11379 40197 11435 40253
rect 11521 40197 11577 40253
rect 11663 40197 11719 40253
rect 11805 40197 11861 40253
rect 11947 40197 12003 40253
rect 12089 40197 12145 40253
rect 12231 40197 12287 40253
rect 12373 40197 12429 40253
rect 12515 40197 12571 40253
rect 12657 40197 12713 40253
rect 12799 40197 12855 40253
rect 12941 40197 12997 40253
rect 13083 40197 13139 40253
rect 13225 40197 13281 40253
rect 13367 40197 13423 40253
rect 13509 40197 13565 40253
rect 13651 40197 13707 40253
rect 13793 40197 13849 40253
rect 13935 40197 13991 40253
rect 14077 40197 14133 40253
rect 14219 40197 14275 40253
rect 14361 40197 14417 40253
rect 14503 40197 14559 40253
rect 14645 40197 14701 40253
rect 14787 40197 14843 40253
rect 161 40055 217 40111
rect 303 40055 359 40111
rect 445 40055 501 40111
rect 587 40055 643 40111
rect 729 40055 785 40111
rect 871 40055 927 40111
rect 1013 40055 1069 40111
rect 1155 40055 1211 40111
rect 1297 40055 1353 40111
rect 1439 40055 1495 40111
rect 1581 40055 1637 40111
rect 1723 40055 1779 40111
rect 1865 40055 1921 40111
rect 2007 40055 2063 40111
rect 2149 40055 2205 40111
rect 2291 40055 2347 40111
rect 2433 40055 2489 40111
rect 2575 40055 2631 40111
rect 2717 40055 2773 40111
rect 2859 40055 2915 40111
rect 3001 40055 3057 40111
rect 3143 40055 3199 40111
rect 3285 40055 3341 40111
rect 3427 40055 3483 40111
rect 3569 40055 3625 40111
rect 3711 40055 3767 40111
rect 3853 40055 3909 40111
rect 3995 40055 4051 40111
rect 4137 40055 4193 40111
rect 4279 40055 4335 40111
rect 4421 40055 4477 40111
rect 4563 40055 4619 40111
rect 4705 40055 4761 40111
rect 4847 40055 4903 40111
rect 4989 40055 5045 40111
rect 5131 40055 5187 40111
rect 5273 40055 5329 40111
rect 5415 40055 5471 40111
rect 5557 40055 5613 40111
rect 5699 40055 5755 40111
rect 5841 40055 5897 40111
rect 5983 40055 6039 40111
rect 6125 40055 6181 40111
rect 6267 40055 6323 40111
rect 6409 40055 6465 40111
rect 6551 40055 6607 40111
rect 6693 40055 6749 40111
rect 6835 40055 6891 40111
rect 6977 40055 7033 40111
rect 7119 40055 7175 40111
rect 7261 40055 7317 40111
rect 7403 40055 7459 40111
rect 7545 40055 7601 40111
rect 7687 40055 7743 40111
rect 7829 40055 7885 40111
rect 7971 40055 8027 40111
rect 8113 40055 8169 40111
rect 8255 40055 8311 40111
rect 8397 40055 8453 40111
rect 8539 40055 8595 40111
rect 8681 40055 8737 40111
rect 8823 40055 8879 40111
rect 8965 40055 9021 40111
rect 9107 40055 9163 40111
rect 9249 40055 9305 40111
rect 9391 40055 9447 40111
rect 9533 40055 9589 40111
rect 9675 40055 9731 40111
rect 9817 40055 9873 40111
rect 9959 40055 10015 40111
rect 10101 40055 10157 40111
rect 10243 40055 10299 40111
rect 10385 40055 10441 40111
rect 10527 40055 10583 40111
rect 10669 40055 10725 40111
rect 10811 40055 10867 40111
rect 10953 40055 11009 40111
rect 11095 40055 11151 40111
rect 11237 40055 11293 40111
rect 11379 40055 11435 40111
rect 11521 40055 11577 40111
rect 11663 40055 11719 40111
rect 11805 40055 11861 40111
rect 11947 40055 12003 40111
rect 12089 40055 12145 40111
rect 12231 40055 12287 40111
rect 12373 40055 12429 40111
rect 12515 40055 12571 40111
rect 12657 40055 12713 40111
rect 12799 40055 12855 40111
rect 12941 40055 12997 40111
rect 13083 40055 13139 40111
rect 13225 40055 13281 40111
rect 13367 40055 13423 40111
rect 13509 40055 13565 40111
rect 13651 40055 13707 40111
rect 13793 40055 13849 40111
rect 13935 40055 13991 40111
rect 14077 40055 14133 40111
rect 14219 40055 14275 40111
rect 14361 40055 14417 40111
rect 14503 40055 14559 40111
rect 14645 40055 14701 40111
rect 14787 40055 14843 40111
rect 161 39913 217 39969
rect 303 39913 359 39969
rect 445 39913 501 39969
rect 587 39913 643 39969
rect 729 39913 785 39969
rect 871 39913 927 39969
rect 1013 39913 1069 39969
rect 1155 39913 1211 39969
rect 1297 39913 1353 39969
rect 1439 39913 1495 39969
rect 1581 39913 1637 39969
rect 1723 39913 1779 39969
rect 1865 39913 1921 39969
rect 2007 39913 2063 39969
rect 2149 39913 2205 39969
rect 2291 39913 2347 39969
rect 2433 39913 2489 39969
rect 2575 39913 2631 39969
rect 2717 39913 2773 39969
rect 2859 39913 2915 39969
rect 3001 39913 3057 39969
rect 3143 39913 3199 39969
rect 3285 39913 3341 39969
rect 3427 39913 3483 39969
rect 3569 39913 3625 39969
rect 3711 39913 3767 39969
rect 3853 39913 3909 39969
rect 3995 39913 4051 39969
rect 4137 39913 4193 39969
rect 4279 39913 4335 39969
rect 4421 39913 4477 39969
rect 4563 39913 4619 39969
rect 4705 39913 4761 39969
rect 4847 39913 4903 39969
rect 4989 39913 5045 39969
rect 5131 39913 5187 39969
rect 5273 39913 5329 39969
rect 5415 39913 5471 39969
rect 5557 39913 5613 39969
rect 5699 39913 5755 39969
rect 5841 39913 5897 39969
rect 5983 39913 6039 39969
rect 6125 39913 6181 39969
rect 6267 39913 6323 39969
rect 6409 39913 6465 39969
rect 6551 39913 6607 39969
rect 6693 39913 6749 39969
rect 6835 39913 6891 39969
rect 6977 39913 7033 39969
rect 7119 39913 7175 39969
rect 7261 39913 7317 39969
rect 7403 39913 7459 39969
rect 7545 39913 7601 39969
rect 7687 39913 7743 39969
rect 7829 39913 7885 39969
rect 7971 39913 8027 39969
rect 8113 39913 8169 39969
rect 8255 39913 8311 39969
rect 8397 39913 8453 39969
rect 8539 39913 8595 39969
rect 8681 39913 8737 39969
rect 8823 39913 8879 39969
rect 8965 39913 9021 39969
rect 9107 39913 9163 39969
rect 9249 39913 9305 39969
rect 9391 39913 9447 39969
rect 9533 39913 9589 39969
rect 9675 39913 9731 39969
rect 9817 39913 9873 39969
rect 9959 39913 10015 39969
rect 10101 39913 10157 39969
rect 10243 39913 10299 39969
rect 10385 39913 10441 39969
rect 10527 39913 10583 39969
rect 10669 39913 10725 39969
rect 10811 39913 10867 39969
rect 10953 39913 11009 39969
rect 11095 39913 11151 39969
rect 11237 39913 11293 39969
rect 11379 39913 11435 39969
rect 11521 39913 11577 39969
rect 11663 39913 11719 39969
rect 11805 39913 11861 39969
rect 11947 39913 12003 39969
rect 12089 39913 12145 39969
rect 12231 39913 12287 39969
rect 12373 39913 12429 39969
rect 12515 39913 12571 39969
rect 12657 39913 12713 39969
rect 12799 39913 12855 39969
rect 12941 39913 12997 39969
rect 13083 39913 13139 39969
rect 13225 39913 13281 39969
rect 13367 39913 13423 39969
rect 13509 39913 13565 39969
rect 13651 39913 13707 39969
rect 13793 39913 13849 39969
rect 13935 39913 13991 39969
rect 14077 39913 14133 39969
rect 14219 39913 14275 39969
rect 14361 39913 14417 39969
rect 14503 39913 14559 39969
rect 14645 39913 14701 39969
rect 14787 39913 14843 39969
rect 161 39771 217 39827
rect 303 39771 359 39827
rect 445 39771 501 39827
rect 587 39771 643 39827
rect 729 39771 785 39827
rect 871 39771 927 39827
rect 1013 39771 1069 39827
rect 1155 39771 1211 39827
rect 1297 39771 1353 39827
rect 1439 39771 1495 39827
rect 1581 39771 1637 39827
rect 1723 39771 1779 39827
rect 1865 39771 1921 39827
rect 2007 39771 2063 39827
rect 2149 39771 2205 39827
rect 2291 39771 2347 39827
rect 2433 39771 2489 39827
rect 2575 39771 2631 39827
rect 2717 39771 2773 39827
rect 2859 39771 2915 39827
rect 3001 39771 3057 39827
rect 3143 39771 3199 39827
rect 3285 39771 3341 39827
rect 3427 39771 3483 39827
rect 3569 39771 3625 39827
rect 3711 39771 3767 39827
rect 3853 39771 3909 39827
rect 3995 39771 4051 39827
rect 4137 39771 4193 39827
rect 4279 39771 4335 39827
rect 4421 39771 4477 39827
rect 4563 39771 4619 39827
rect 4705 39771 4761 39827
rect 4847 39771 4903 39827
rect 4989 39771 5045 39827
rect 5131 39771 5187 39827
rect 5273 39771 5329 39827
rect 5415 39771 5471 39827
rect 5557 39771 5613 39827
rect 5699 39771 5755 39827
rect 5841 39771 5897 39827
rect 5983 39771 6039 39827
rect 6125 39771 6181 39827
rect 6267 39771 6323 39827
rect 6409 39771 6465 39827
rect 6551 39771 6607 39827
rect 6693 39771 6749 39827
rect 6835 39771 6891 39827
rect 6977 39771 7033 39827
rect 7119 39771 7175 39827
rect 7261 39771 7317 39827
rect 7403 39771 7459 39827
rect 7545 39771 7601 39827
rect 7687 39771 7743 39827
rect 7829 39771 7885 39827
rect 7971 39771 8027 39827
rect 8113 39771 8169 39827
rect 8255 39771 8311 39827
rect 8397 39771 8453 39827
rect 8539 39771 8595 39827
rect 8681 39771 8737 39827
rect 8823 39771 8879 39827
rect 8965 39771 9021 39827
rect 9107 39771 9163 39827
rect 9249 39771 9305 39827
rect 9391 39771 9447 39827
rect 9533 39771 9589 39827
rect 9675 39771 9731 39827
rect 9817 39771 9873 39827
rect 9959 39771 10015 39827
rect 10101 39771 10157 39827
rect 10243 39771 10299 39827
rect 10385 39771 10441 39827
rect 10527 39771 10583 39827
rect 10669 39771 10725 39827
rect 10811 39771 10867 39827
rect 10953 39771 11009 39827
rect 11095 39771 11151 39827
rect 11237 39771 11293 39827
rect 11379 39771 11435 39827
rect 11521 39771 11577 39827
rect 11663 39771 11719 39827
rect 11805 39771 11861 39827
rect 11947 39771 12003 39827
rect 12089 39771 12145 39827
rect 12231 39771 12287 39827
rect 12373 39771 12429 39827
rect 12515 39771 12571 39827
rect 12657 39771 12713 39827
rect 12799 39771 12855 39827
rect 12941 39771 12997 39827
rect 13083 39771 13139 39827
rect 13225 39771 13281 39827
rect 13367 39771 13423 39827
rect 13509 39771 13565 39827
rect 13651 39771 13707 39827
rect 13793 39771 13849 39827
rect 13935 39771 13991 39827
rect 14077 39771 14133 39827
rect 14219 39771 14275 39827
rect 14361 39771 14417 39827
rect 14503 39771 14559 39827
rect 14645 39771 14701 39827
rect 14787 39771 14843 39827
rect 161 39629 217 39685
rect 303 39629 359 39685
rect 445 39629 501 39685
rect 587 39629 643 39685
rect 729 39629 785 39685
rect 871 39629 927 39685
rect 1013 39629 1069 39685
rect 1155 39629 1211 39685
rect 1297 39629 1353 39685
rect 1439 39629 1495 39685
rect 1581 39629 1637 39685
rect 1723 39629 1779 39685
rect 1865 39629 1921 39685
rect 2007 39629 2063 39685
rect 2149 39629 2205 39685
rect 2291 39629 2347 39685
rect 2433 39629 2489 39685
rect 2575 39629 2631 39685
rect 2717 39629 2773 39685
rect 2859 39629 2915 39685
rect 3001 39629 3057 39685
rect 3143 39629 3199 39685
rect 3285 39629 3341 39685
rect 3427 39629 3483 39685
rect 3569 39629 3625 39685
rect 3711 39629 3767 39685
rect 3853 39629 3909 39685
rect 3995 39629 4051 39685
rect 4137 39629 4193 39685
rect 4279 39629 4335 39685
rect 4421 39629 4477 39685
rect 4563 39629 4619 39685
rect 4705 39629 4761 39685
rect 4847 39629 4903 39685
rect 4989 39629 5045 39685
rect 5131 39629 5187 39685
rect 5273 39629 5329 39685
rect 5415 39629 5471 39685
rect 5557 39629 5613 39685
rect 5699 39629 5755 39685
rect 5841 39629 5897 39685
rect 5983 39629 6039 39685
rect 6125 39629 6181 39685
rect 6267 39629 6323 39685
rect 6409 39629 6465 39685
rect 6551 39629 6607 39685
rect 6693 39629 6749 39685
rect 6835 39629 6891 39685
rect 6977 39629 7033 39685
rect 7119 39629 7175 39685
rect 7261 39629 7317 39685
rect 7403 39629 7459 39685
rect 7545 39629 7601 39685
rect 7687 39629 7743 39685
rect 7829 39629 7885 39685
rect 7971 39629 8027 39685
rect 8113 39629 8169 39685
rect 8255 39629 8311 39685
rect 8397 39629 8453 39685
rect 8539 39629 8595 39685
rect 8681 39629 8737 39685
rect 8823 39629 8879 39685
rect 8965 39629 9021 39685
rect 9107 39629 9163 39685
rect 9249 39629 9305 39685
rect 9391 39629 9447 39685
rect 9533 39629 9589 39685
rect 9675 39629 9731 39685
rect 9817 39629 9873 39685
rect 9959 39629 10015 39685
rect 10101 39629 10157 39685
rect 10243 39629 10299 39685
rect 10385 39629 10441 39685
rect 10527 39629 10583 39685
rect 10669 39629 10725 39685
rect 10811 39629 10867 39685
rect 10953 39629 11009 39685
rect 11095 39629 11151 39685
rect 11237 39629 11293 39685
rect 11379 39629 11435 39685
rect 11521 39629 11577 39685
rect 11663 39629 11719 39685
rect 11805 39629 11861 39685
rect 11947 39629 12003 39685
rect 12089 39629 12145 39685
rect 12231 39629 12287 39685
rect 12373 39629 12429 39685
rect 12515 39629 12571 39685
rect 12657 39629 12713 39685
rect 12799 39629 12855 39685
rect 12941 39629 12997 39685
rect 13083 39629 13139 39685
rect 13225 39629 13281 39685
rect 13367 39629 13423 39685
rect 13509 39629 13565 39685
rect 13651 39629 13707 39685
rect 13793 39629 13849 39685
rect 13935 39629 13991 39685
rect 14077 39629 14133 39685
rect 14219 39629 14275 39685
rect 14361 39629 14417 39685
rect 14503 39629 14559 39685
rect 14645 39629 14701 39685
rect 14787 39629 14843 39685
rect 161 39286 217 39342
rect 303 39286 359 39342
rect 445 39286 501 39342
rect 587 39286 643 39342
rect 729 39286 785 39342
rect 871 39286 927 39342
rect 1013 39286 1069 39342
rect 1155 39286 1211 39342
rect 1297 39286 1353 39342
rect 1439 39286 1495 39342
rect 1581 39286 1637 39342
rect 1723 39286 1779 39342
rect 1865 39286 1921 39342
rect 2007 39286 2063 39342
rect 2149 39286 2205 39342
rect 2291 39286 2347 39342
rect 2433 39286 2489 39342
rect 2575 39286 2631 39342
rect 2717 39286 2773 39342
rect 2859 39286 2915 39342
rect 3001 39286 3057 39342
rect 3143 39286 3199 39342
rect 3285 39286 3341 39342
rect 3427 39286 3483 39342
rect 3569 39286 3625 39342
rect 3711 39286 3767 39342
rect 3853 39286 3909 39342
rect 3995 39286 4051 39342
rect 4137 39286 4193 39342
rect 4279 39286 4335 39342
rect 4421 39286 4477 39342
rect 4563 39286 4619 39342
rect 4705 39286 4761 39342
rect 4847 39286 4903 39342
rect 4989 39286 5045 39342
rect 5131 39286 5187 39342
rect 5273 39286 5329 39342
rect 5415 39286 5471 39342
rect 5557 39286 5613 39342
rect 5699 39286 5755 39342
rect 5841 39286 5897 39342
rect 5983 39286 6039 39342
rect 6125 39286 6181 39342
rect 6267 39286 6323 39342
rect 6409 39286 6465 39342
rect 6551 39286 6607 39342
rect 6693 39286 6749 39342
rect 6835 39286 6891 39342
rect 6977 39286 7033 39342
rect 7119 39286 7175 39342
rect 7261 39286 7317 39342
rect 7403 39286 7459 39342
rect 7545 39286 7601 39342
rect 7687 39286 7743 39342
rect 7829 39286 7885 39342
rect 7971 39286 8027 39342
rect 8113 39286 8169 39342
rect 8255 39286 8311 39342
rect 8397 39286 8453 39342
rect 8539 39286 8595 39342
rect 8681 39286 8737 39342
rect 8823 39286 8879 39342
rect 8965 39286 9021 39342
rect 9107 39286 9163 39342
rect 9249 39286 9305 39342
rect 9391 39286 9447 39342
rect 9533 39286 9589 39342
rect 9675 39286 9731 39342
rect 9817 39286 9873 39342
rect 9959 39286 10015 39342
rect 10101 39286 10157 39342
rect 10243 39286 10299 39342
rect 10385 39286 10441 39342
rect 10527 39286 10583 39342
rect 10669 39286 10725 39342
rect 10811 39286 10867 39342
rect 10953 39286 11009 39342
rect 11095 39286 11151 39342
rect 11237 39286 11293 39342
rect 11379 39286 11435 39342
rect 11521 39286 11577 39342
rect 11663 39286 11719 39342
rect 11805 39286 11861 39342
rect 11947 39286 12003 39342
rect 12089 39286 12145 39342
rect 12231 39286 12287 39342
rect 12373 39286 12429 39342
rect 12515 39286 12571 39342
rect 12657 39286 12713 39342
rect 12799 39286 12855 39342
rect 12941 39286 12997 39342
rect 13083 39286 13139 39342
rect 13225 39286 13281 39342
rect 13367 39286 13423 39342
rect 13509 39286 13565 39342
rect 13651 39286 13707 39342
rect 13793 39286 13849 39342
rect 13935 39286 13991 39342
rect 14077 39286 14133 39342
rect 14219 39286 14275 39342
rect 14361 39286 14417 39342
rect 14503 39286 14559 39342
rect 14645 39286 14701 39342
rect 14787 39286 14843 39342
rect 161 39144 217 39200
rect 303 39144 359 39200
rect 445 39144 501 39200
rect 587 39144 643 39200
rect 729 39144 785 39200
rect 871 39144 927 39200
rect 1013 39144 1069 39200
rect 1155 39144 1211 39200
rect 1297 39144 1353 39200
rect 1439 39144 1495 39200
rect 1581 39144 1637 39200
rect 1723 39144 1779 39200
rect 1865 39144 1921 39200
rect 2007 39144 2063 39200
rect 2149 39144 2205 39200
rect 2291 39144 2347 39200
rect 2433 39144 2489 39200
rect 2575 39144 2631 39200
rect 2717 39144 2773 39200
rect 2859 39144 2915 39200
rect 3001 39144 3057 39200
rect 3143 39144 3199 39200
rect 3285 39144 3341 39200
rect 3427 39144 3483 39200
rect 3569 39144 3625 39200
rect 3711 39144 3767 39200
rect 3853 39144 3909 39200
rect 3995 39144 4051 39200
rect 4137 39144 4193 39200
rect 4279 39144 4335 39200
rect 4421 39144 4477 39200
rect 4563 39144 4619 39200
rect 4705 39144 4761 39200
rect 4847 39144 4903 39200
rect 4989 39144 5045 39200
rect 5131 39144 5187 39200
rect 5273 39144 5329 39200
rect 5415 39144 5471 39200
rect 5557 39144 5613 39200
rect 5699 39144 5755 39200
rect 5841 39144 5897 39200
rect 5983 39144 6039 39200
rect 6125 39144 6181 39200
rect 6267 39144 6323 39200
rect 6409 39144 6465 39200
rect 6551 39144 6607 39200
rect 6693 39144 6749 39200
rect 6835 39144 6891 39200
rect 6977 39144 7033 39200
rect 7119 39144 7175 39200
rect 7261 39144 7317 39200
rect 7403 39144 7459 39200
rect 7545 39144 7601 39200
rect 7687 39144 7743 39200
rect 7829 39144 7885 39200
rect 7971 39144 8027 39200
rect 8113 39144 8169 39200
rect 8255 39144 8311 39200
rect 8397 39144 8453 39200
rect 8539 39144 8595 39200
rect 8681 39144 8737 39200
rect 8823 39144 8879 39200
rect 8965 39144 9021 39200
rect 9107 39144 9163 39200
rect 9249 39144 9305 39200
rect 9391 39144 9447 39200
rect 9533 39144 9589 39200
rect 9675 39144 9731 39200
rect 9817 39144 9873 39200
rect 9959 39144 10015 39200
rect 10101 39144 10157 39200
rect 10243 39144 10299 39200
rect 10385 39144 10441 39200
rect 10527 39144 10583 39200
rect 10669 39144 10725 39200
rect 10811 39144 10867 39200
rect 10953 39144 11009 39200
rect 11095 39144 11151 39200
rect 11237 39144 11293 39200
rect 11379 39144 11435 39200
rect 11521 39144 11577 39200
rect 11663 39144 11719 39200
rect 11805 39144 11861 39200
rect 11947 39144 12003 39200
rect 12089 39144 12145 39200
rect 12231 39144 12287 39200
rect 12373 39144 12429 39200
rect 12515 39144 12571 39200
rect 12657 39144 12713 39200
rect 12799 39144 12855 39200
rect 12941 39144 12997 39200
rect 13083 39144 13139 39200
rect 13225 39144 13281 39200
rect 13367 39144 13423 39200
rect 13509 39144 13565 39200
rect 13651 39144 13707 39200
rect 13793 39144 13849 39200
rect 13935 39144 13991 39200
rect 14077 39144 14133 39200
rect 14219 39144 14275 39200
rect 14361 39144 14417 39200
rect 14503 39144 14559 39200
rect 14645 39144 14701 39200
rect 14787 39144 14843 39200
rect 161 39002 217 39058
rect 303 39002 359 39058
rect 445 39002 501 39058
rect 587 39002 643 39058
rect 729 39002 785 39058
rect 871 39002 927 39058
rect 1013 39002 1069 39058
rect 1155 39002 1211 39058
rect 1297 39002 1353 39058
rect 1439 39002 1495 39058
rect 1581 39002 1637 39058
rect 1723 39002 1779 39058
rect 1865 39002 1921 39058
rect 2007 39002 2063 39058
rect 2149 39002 2205 39058
rect 2291 39002 2347 39058
rect 2433 39002 2489 39058
rect 2575 39002 2631 39058
rect 2717 39002 2773 39058
rect 2859 39002 2915 39058
rect 3001 39002 3057 39058
rect 3143 39002 3199 39058
rect 3285 39002 3341 39058
rect 3427 39002 3483 39058
rect 3569 39002 3625 39058
rect 3711 39002 3767 39058
rect 3853 39002 3909 39058
rect 3995 39002 4051 39058
rect 4137 39002 4193 39058
rect 4279 39002 4335 39058
rect 4421 39002 4477 39058
rect 4563 39002 4619 39058
rect 4705 39002 4761 39058
rect 4847 39002 4903 39058
rect 4989 39002 5045 39058
rect 5131 39002 5187 39058
rect 5273 39002 5329 39058
rect 5415 39002 5471 39058
rect 5557 39002 5613 39058
rect 5699 39002 5755 39058
rect 5841 39002 5897 39058
rect 5983 39002 6039 39058
rect 6125 39002 6181 39058
rect 6267 39002 6323 39058
rect 6409 39002 6465 39058
rect 6551 39002 6607 39058
rect 6693 39002 6749 39058
rect 6835 39002 6891 39058
rect 6977 39002 7033 39058
rect 7119 39002 7175 39058
rect 7261 39002 7317 39058
rect 7403 39002 7459 39058
rect 7545 39002 7601 39058
rect 7687 39002 7743 39058
rect 7829 39002 7885 39058
rect 7971 39002 8027 39058
rect 8113 39002 8169 39058
rect 8255 39002 8311 39058
rect 8397 39002 8453 39058
rect 8539 39002 8595 39058
rect 8681 39002 8737 39058
rect 8823 39002 8879 39058
rect 8965 39002 9021 39058
rect 9107 39002 9163 39058
rect 9249 39002 9305 39058
rect 9391 39002 9447 39058
rect 9533 39002 9589 39058
rect 9675 39002 9731 39058
rect 9817 39002 9873 39058
rect 9959 39002 10015 39058
rect 10101 39002 10157 39058
rect 10243 39002 10299 39058
rect 10385 39002 10441 39058
rect 10527 39002 10583 39058
rect 10669 39002 10725 39058
rect 10811 39002 10867 39058
rect 10953 39002 11009 39058
rect 11095 39002 11151 39058
rect 11237 39002 11293 39058
rect 11379 39002 11435 39058
rect 11521 39002 11577 39058
rect 11663 39002 11719 39058
rect 11805 39002 11861 39058
rect 11947 39002 12003 39058
rect 12089 39002 12145 39058
rect 12231 39002 12287 39058
rect 12373 39002 12429 39058
rect 12515 39002 12571 39058
rect 12657 39002 12713 39058
rect 12799 39002 12855 39058
rect 12941 39002 12997 39058
rect 13083 39002 13139 39058
rect 13225 39002 13281 39058
rect 13367 39002 13423 39058
rect 13509 39002 13565 39058
rect 13651 39002 13707 39058
rect 13793 39002 13849 39058
rect 13935 39002 13991 39058
rect 14077 39002 14133 39058
rect 14219 39002 14275 39058
rect 14361 39002 14417 39058
rect 14503 39002 14559 39058
rect 14645 39002 14701 39058
rect 14787 39002 14843 39058
rect 161 38860 217 38916
rect 303 38860 359 38916
rect 445 38860 501 38916
rect 587 38860 643 38916
rect 729 38860 785 38916
rect 871 38860 927 38916
rect 1013 38860 1069 38916
rect 1155 38860 1211 38916
rect 1297 38860 1353 38916
rect 1439 38860 1495 38916
rect 1581 38860 1637 38916
rect 1723 38860 1779 38916
rect 1865 38860 1921 38916
rect 2007 38860 2063 38916
rect 2149 38860 2205 38916
rect 2291 38860 2347 38916
rect 2433 38860 2489 38916
rect 2575 38860 2631 38916
rect 2717 38860 2773 38916
rect 2859 38860 2915 38916
rect 3001 38860 3057 38916
rect 3143 38860 3199 38916
rect 3285 38860 3341 38916
rect 3427 38860 3483 38916
rect 3569 38860 3625 38916
rect 3711 38860 3767 38916
rect 3853 38860 3909 38916
rect 3995 38860 4051 38916
rect 4137 38860 4193 38916
rect 4279 38860 4335 38916
rect 4421 38860 4477 38916
rect 4563 38860 4619 38916
rect 4705 38860 4761 38916
rect 4847 38860 4903 38916
rect 4989 38860 5045 38916
rect 5131 38860 5187 38916
rect 5273 38860 5329 38916
rect 5415 38860 5471 38916
rect 5557 38860 5613 38916
rect 5699 38860 5755 38916
rect 5841 38860 5897 38916
rect 5983 38860 6039 38916
rect 6125 38860 6181 38916
rect 6267 38860 6323 38916
rect 6409 38860 6465 38916
rect 6551 38860 6607 38916
rect 6693 38860 6749 38916
rect 6835 38860 6891 38916
rect 6977 38860 7033 38916
rect 7119 38860 7175 38916
rect 7261 38860 7317 38916
rect 7403 38860 7459 38916
rect 7545 38860 7601 38916
rect 7687 38860 7743 38916
rect 7829 38860 7885 38916
rect 7971 38860 8027 38916
rect 8113 38860 8169 38916
rect 8255 38860 8311 38916
rect 8397 38860 8453 38916
rect 8539 38860 8595 38916
rect 8681 38860 8737 38916
rect 8823 38860 8879 38916
rect 8965 38860 9021 38916
rect 9107 38860 9163 38916
rect 9249 38860 9305 38916
rect 9391 38860 9447 38916
rect 9533 38860 9589 38916
rect 9675 38860 9731 38916
rect 9817 38860 9873 38916
rect 9959 38860 10015 38916
rect 10101 38860 10157 38916
rect 10243 38860 10299 38916
rect 10385 38860 10441 38916
rect 10527 38860 10583 38916
rect 10669 38860 10725 38916
rect 10811 38860 10867 38916
rect 10953 38860 11009 38916
rect 11095 38860 11151 38916
rect 11237 38860 11293 38916
rect 11379 38860 11435 38916
rect 11521 38860 11577 38916
rect 11663 38860 11719 38916
rect 11805 38860 11861 38916
rect 11947 38860 12003 38916
rect 12089 38860 12145 38916
rect 12231 38860 12287 38916
rect 12373 38860 12429 38916
rect 12515 38860 12571 38916
rect 12657 38860 12713 38916
rect 12799 38860 12855 38916
rect 12941 38860 12997 38916
rect 13083 38860 13139 38916
rect 13225 38860 13281 38916
rect 13367 38860 13423 38916
rect 13509 38860 13565 38916
rect 13651 38860 13707 38916
rect 13793 38860 13849 38916
rect 13935 38860 13991 38916
rect 14077 38860 14133 38916
rect 14219 38860 14275 38916
rect 14361 38860 14417 38916
rect 14503 38860 14559 38916
rect 14645 38860 14701 38916
rect 14787 38860 14843 38916
rect 161 38718 217 38774
rect 303 38718 359 38774
rect 445 38718 501 38774
rect 587 38718 643 38774
rect 729 38718 785 38774
rect 871 38718 927 38774
rect 1013 38718 1069 38774
rect 1155 38718 1211 38774
rect 1297 38718 1353 38774
rect 1439 38718 1495 38774
rect 1581 38718 1637 38774
rect 1723 38718 1779 38774
rect 1865 38718 1921 38774
rect 2007 38718 2063 38774
rect 2149 38718 2205 38774
rect 2291 38718 2347 38774
rect 2433 38718 2489 38774
rect 2575 38718 2631 38774
rect 2717 38718 2773 38774
rect 2859 38718 2915 38774
rect 3001 38718 3057 38774
rect 3143 38718 3199 38774
rect 3285 38718 3341 38774
rect 3427 38718 3483 38774
rect 3569 38718 3625 38774
rect 3711 38718 3767 38774
rect 3853 38718 3909 38774
rect 3995 38718 4051 38774
rect 4137 38718 4193 38774
rect 4279 38718 4335 38774
rect 4421 38718 4477 38774
rect 4563 38718 4619 38774
rect 4705 38718 4761 38774
rect 4847 38718 4903 38774
rect 4989 38718 5045 38774
rect 5131 38718 5187 38774
rect 5273 38718 5329 38774
rect 5415 38718 5471 38774
rect 5557 38718 5613 38774
rect 5699 38718 5755 38774
rect 5841 38718 5897 38774
rect 5983 38718 6039 38774
rect 6125 38718 6181 38774
rect 6267 38718 6323 38774
rect 6409 38718 6465 38774
rect 6551 38718 6607 38774
rect 6693 38718 6749 38774
rect 6835 38718 6891 38774
rect 6977 38718 7033 38774
rect 7119 38718 7175 38774
rect 7261 38718 7317 38774
rect 7403 38718 7459 38774
rect 7545 38718 7601 38774
rect 7687 38718 7743 38774
rect 7829 38718 7885 38774
rect 7971 38718 8027 38774
rect 8113 38718 8169 38774
rect 8255 38718 8311 38774
rect 8397 38718 8453 38774
rect 8539 38718 8595 38774
rect 8681 38718 8737 38774
rect 8823 38718 8879 38774
rect 8965 38718 9021 38774
rect 9107 38718 9163 38774
rect 9249 38718 9305 38774
rect 9391 38718 9447 38774
rect 9533 38718 9589 38774
rect 9675 38718 9731 38774
rect 9817 38718 9873 38774
rect 9959 38718 10015 38774
rect 10101 38718 10157 38774
rect 10243 38718 10299 38774
rect 10385 38718 10441 38774
rect 10527 38718 10583 38774
rect 10669 38718 10725 38774
rect 10811 38718 10867 38774
rect 10953 38718 11009 38774
rect 11095 38718 11151 38774
rect 11237 38718 11293 38774
rect 11379 38718 11435 38774
rect 11521 38718 11577 38774
rect 11663 38718 11719 38774
rect 11805 38718 11861 38774
rect 11947 38718 12003 38774
rect 12089 38718 12145 38774
rect 12231 38718 12287 38774
rect 12373 38718 12429 38774
rect 12515 38718 12571 38774
rect 12657 38718 12713 38774
rect 12799 38718 12855 38774
rect 12941 38718 12997 38774
rect 13083 38718 13139 38774
rect 13225 38718 13281 38774
rect 13367 38718 13423 38774
rect 13509 38718 13565 38774
rect 13651 38718 13707 38774
rect 13793 38718 13849 38774
rect 13935 38718 13991 38774
rect 14077 38718 14133 38774
rect 14219 38718 14275 38774
rect 14361 38718 14417 38774
rect 14503 38718 14559 38774
rect 14645 38718 14701 38774
rect 14787 38718 14843 38774
rect 161 38576 217 38632
rect 303 38576 359 38632
rect 445 38576 501 38632
rect 587 38576 643 38632
rect 729 38576 785 38632
rect 871 38576 927 38632
rect 1013 38576 1069 38632
rect 1155 38576 1211 38632
rect 1297 38576 1353 38632
rect 1439 38576 1495 38632
rect 1581 38576 1637 38632
rect 1723 38576 1779 38632
rect 1865 38576 1921 38632
rect 2007 38576 2063 38632
rect 2149 38576 2205 38632
rect 2291 38576 2347 38632
rect 2433 38576 2489 38632
rect 2575 38576 2631 38632
rect 2717 38576 2773 38632
rect 2859 38576 2915 38632
rect 3001 38576 3057 38632
rect 3143 38576 3199 38632
rect 3285 38576 3341 38632
rect 3427 38576 3483 38632
rect 3569 38576 3625 38632
rect 3711 38576 3767 38632
rect 3853 38576 3909 38632
rect 3995 38576 4051 38632
rect 4137 38576 4193 38632
rect 4279 38576 4335 38632
rect 4421 38576 4477 38632
rect 4563 38576 4619 38632
rect 4705 38576 4761 38632
rect 4847 38576 4903 38632
rect 4989 38576 5045 38632
rect 5131 38576 5187 38632
rect 5273 38576 5329 38632
rect 5415 38576 5471 38632
rect 5557 38576 5613 38632
rect 5699 38576 5755 38632
rect 5841 38576 5897 38632
rect 5983 38576 6039 38632
rect 6125 38576 6181 38632
rect 6267 38576 6323 38632
rect 6409 38576 6465 38632
rect 6551 38576 6607 38632
rect 6693 38576 6749 38632
rect 6835 38576 6891 38632
rect 6977 38576 7033 38632
rect 7119 38576 7175 38632
rect 7261 38576 7317 38632
rect 7403 38576 7459 38632
rect 7545 38576 7601 38632
rect 7687 38576 7743 38632
rect 7829 38576 7885 38632
rect 7971 38576 8027 38632
rect 8113 38576 8169 38632
rect 8255 38576 8311 38632
rect 8397 38576 8453 38632
rect 8539 38576 8595 38632
rect 8681 38576 8737 38632
rect 8823 38576 8879 38632
rect 8965 38576 9021 38632
rect 9107 38576 9163 38632
rect 9249 38576 9305 38632
rect 9391 38576 9447 38632
rect 9533 38576 9589 38632
rect 9675 38576 9731 38632
rect 9817 38576 9873 38632
rect 9959 38576 10015 38632
rect 10101 38576 10157 38632
rect 10243 38576 10299 38632
rect 10385 38576 10441 38632
rect 10527 38576 10583 38632
rect 10669 38576 10725 38632
rect 10811 38576 10867 38632
rect 10953 38576 11009 38632
rect 11095 38576 11151 38632
rect 11237 38576 11293 38632
rect 11379 38576 11435 38632
rect 11521 38576 11577 38632
rect 11663 38576 11719 38632
rect 11805 38576 11861 38632
rect 11947 38576 12003 38632
rect 12089 38576 12145 38632
rect 12231 38576 12287 38632
rect 12373 38576 12429 38632
rect 12515 38576 12571 38632
rect 12657 38576 12713 38632
rect 12799 38576 12855 38632
rect 12941 38576 12997 38632
rect 13083 38576 13139 38632
rect 13225 38576 13281 38632
rect 13367 38576 13423 38632
rect 13509 38576 13565 38632
rect 13651 38576 13707 38632
rect 13793 38576 13849 38632
rect 13935 38576 13991 38632
rect 14077 38576 14133 38632
rect 14219 38576 14275 38632
rect 14361 38576 14417 38632
rect 14503 38576 14559 38632
rect 14645 38576 14701 38632
rect 14787 38576 14843 38632
rect 161 38434 217 38490
rect 303 38434 359 38490
rect 445 38434 501 38490
rect 587 38434 643 38490
rect 729 38434 785 38490
rect 871 38434 927 38490
rect 1013 38434 1069 38490
rect 1155 38434 1211 38490
rect 1297 38434 1353 38490
rect 1439 38434 1495 38490
rect 1581 38434 1637 38490
rect 1723 38434 1779 38490
rect 1865 38434 1921 38490
rect 2007 38434 2063 38490
rect 2149 38434 2205 38490
rect 2291 38434 2347 38490
rect 2433 38434 2489 38490
rect 2575 38434 2631 38490
rect 2717 38434 2773 38490
rect 2859 38434 2915 38490
rect 3001 38434 3057 38490
rect 3143 38434 3199 38490
rect 3285 38434 3341 38490
rect 3427 38434 3483 38490
rect 3569 38434 3625 38490
rect 3711 38434 3767 38490
rect 3853 38434 3909 38490
rect 3995 38434 4051 38490
rect 4137 38434 4193 38490
rect 4279 38434 4335 38490
rect 4421 38434 4477 38490
rect 4563 38434 4619 38490
rect 4705 38434 4761 38490
rect 4847 38434 4903 38490
rect 4989 38434 5045 38490
rect 5131 38434 5187 38490
rect 5273 38434 5329 38490
rect 5415 38434 5471 38490
rect 5557 38434 5613 38490
rect 5699 38434 5755 38490
rect 5841 38434 5897 38490
rect 5983 38434 6039 38490
rect 6125 38434 6181 38490
rect 6267 38434 6323 38490
rect 6409 38434 6465 38490
rect 6551 38434 6607 38490
rect 6693 38434 6749 38490
rect 6835 38434 6891 38490
rect 6977 38434 7033 38490
rect 7119 38434 7175 38490
rect 7261 38434 7317 38490
rect 7403 38434 7459 38490
rect 7545 38434 7601 38490
rect 7687 38434 7743 38490
rect 7829 38434 7885 38490
rect 7971 38434 8027 38490
rect 8113 38434 8169 38490
rect 8255 38434 8311 38490
rect 8397 38434 8453 38490
rect 8539 38434 8595 38490
rect 8681 38434 8737 38490
rect 8823 38434 8879 38490
rect 8965 38434 9021 38490
rect 9107 38434 9163 38490
rect 9249 38434 9305 38490
rect 9391 38434 9447 38490
rect 9533 38434 9589 38490
rect 9675 38434 9731 38490
rect 9817 38434 9873 38490
rect 9959 38434 10015 38490
rect 10101 38434 10157 38490
rect 10243 38434 10299 38490
rect 10385 38434 10441 38490
rect 10527 38434 10583 38490
rect 10669 38434 10725 38490
rect 10811 38434 10867 38490
rect 10953 38434 11009 38490
rect 11095 38434 11151 38490
rect 11237 38434 11293 38490
rect 11379 38434 11435 38490
rect 11521 38434 11577 38490
rect 11663 38434 11719 38490
rect 11805 38434 11861 38490
rect 11947 38434 12003 38490
rect 12089 38434 12145 38490
rect 12231 38434 12287 38490
rect 12373 38434 12429 38490
rect 12515 38434 12571 38490
rect 12657 38434 12713 38490
rect 12799 38434 12855 38490
rect 12941 38434 12997 38490
rect 13083 38434 13139 38490
rect 13225 38434 13281 38490
rect 13367 38434 13423 38490
rect 13509 38434 13565 38490
rect 13651 38434 13707 38490
rect 13793 38434 13849 38490
rect 13935 38434 13991 38490
rect 14077 38434 14133 38490
rect 14219 38434 14275 38490
rect 14361 38434 14417 38490
rect 14503 38434 14559 38490
rect 14645 38434 14701 38490
rect 14787 38434 14843 38490
rect 161 38292 217 38348
rect 303 38292 359 38348
rect 445 38292 501 38348
rect 587 38292 643 38348
rect 729 38292 785 38348
rect 871 38292 927 38348
rect 1013 38292 1069 38348
rect 1155 38292 1211 38348
rect 1297 38292 1353 38348
rect 1439 38292 1495 38348
rect 1581 38292 1637 38348
rect 1723 38292 1779 38348
rect 1865 38292 1921 38348
rect 2007 38292 2063 38348
rect 2149 38292 2205 38348
rect 2291 38292 2347 38348
rect 2433 38292 2489 38348
rect 2575 38292 2631 38348
rect 2717 38292 2773 38348
rect 2859 38292 2915 38348
rect 3001 38292 3057 38348
rect 3143 38292 3199 38348
rect 3285 38292 3341 38348
rect 3427 38292 3483 38348
rect 3569 38292 3625 38348
rect 3711 38292 3767 38348
rect 3853 38292 3909 38348
rect 3995 38292 4051 38348
rect 4137 38292 4193 38348
rect 4279 38292 4335 38348
rect 4421 38292 4477 38348
rect 4563 38292 4619 38348
rect 4705 38292 4761 38348
rect 4847 38292 4903 38348
rect 4989 38292 5045 38348
rect 5131 38292 5187 38348
rect 5273 38292 5329 38348
rect 5415 38292 5471 38348
rect 5557 38292 5613 38348
rect 5699 38292 5755 38348
rect 5841 38292 5897 38348
rect 5983 38292 6039 38348
rect 6125 38292 6181 38348
rect 6267 38292 6323 38348
rect 6409 38292 6465 38348
rect 6551 38292 6607 38348
rect 6693 38292 6749 38348
rect 6835 38292 6891 38348
rect 6977 38292 7033 38348
rect 7119 38292 7175 38348
rect 7261 38292 7317 38348
rect 7403 38292 7459 38348
rect 7545 38292 7601 38348
rect 7687 38292 7743 38348
rect 7829 38292 7885 38348
rect 7971 38292 8027 38348
rect 8113 38292 8169 38348
rect 8255 38292 8311 38348
rect 8397 38292 8453 38348
rect 8539 38292 8595 38348
rect 8681 38292 8737 38348
rect 8823 38292 8879 38348
rect 8965 38292 9021 38348
rect 9107 38292 9163 38348
rect 9249 38292 9305 38348
rect 9391 38292 9447 38348
rect 9533 38292 9589 38348
rect 9675 38292 9731 38348
rect 9817 38292 9873 38348
rect 9959 38292 10015 38348
rect 10101 38292 10157 38348
rect 10243 38292 10299 38348
rect 10385 38292 10441 38348
rect 10527 38292 10583 38348
rect 10669 38292 10725 38348
rect 10811 38292 10867 38348
rect 10953 38292 11009 38348
rect 11095 38292 11151 38348
rect 11237 38292 11293 38348
rect 11379 38292 11435 38348
rect 11521 38292 11577 38348
rect 11663 38292 11719 38348
rect 11805 38292 11861 38348
rect 11947 38292 12003 38348
rect 12089 38292 12145 38348
rect 12231 38292 12287 38348
rect 12373 38292 12429 38348
rect 12515 38292 12571 38348
rect 12657 38292 12713 38348
rect 12799 38292 12855 38348
rect 12941 38292 12997 38348
rect 13083 38292 13139 38348
rect 13225 38292 13281 38348
rect 13367 38292 13423 38348
rect 13509 38292 13565 38348
rect 13651 38292 13707 38348
rect 13793 38292 13849 38348
rect 13935 38292 13991 38348
rect 14077 38292 14133 38348
rect 14219 38292 14275 38348
rect 14361 38292 14417 38348
rect 14503 38292 14559 38348
rect 14645 38292 14701 38348
rect 14787 38292 14843 38348
rect 161 38150 217 38206
rect 303 38150 359 38206
rect 445 38150 501 38206
rect 587 38150 643 38206
rect 729 38150 785 38206
rect 871 38150 927 38206
rect 1013 38150 1069 38206
rect 1155 38150 1211 38206
rect 1297 38150 1353 38206
rect 1439 38150 1495 38206
rect 1581 38150 1637 38206
rect 1723 38150 1779 38206
rect 1865 38150 1921 38206
rect 2007 38150 2063 38206
rect 2149 38150 2205 38206
rect 2291 38150 2347 38206
rect 2433 38150 2489 38206
rect 2575 38150 2631 38206
rect 2717 38150 2773 38206
rect 2859 38150 2915 38206
rect 3001 38150 3057 38206
rect 3143 38150 3199 38206
rect 3285 38150 3341 38206
rect 3427 38150 3483 38206
rect 3569 38150 3625 38206
rect 3711 38150 3767 38206
rect 3853 38150 3909 38206
rect 3995 38150 4051 38206
rect 4137 38150 4193 38206
rect 4279 38150 4335 38206
rect 4421 38150 4477 38206
rect 4563 38150 4619 38206
rect 4705 38150 4761 38206
rect 4847 38150 4903 38206
rect 4989 38150 5045 38206
rect 5131 38150 5187 38206
rect 5273 38150 5329 38206
rect 5415 38150 5471 38206
rect 5557 38150 5613 38206
rect 5699 38150 5755 38206
rect 5841 38150 5897 38206
rect 5983 38150 6039 38206
rect 6125 38150 6181 38206
rect 6267 38150 6323 38206
rect 6409 38150 6465 38206
rect 6551 38150 6607 38206
rect 6693 38150 6749 38206
rect 6835 38150 6891 38206
rect 6977 38150 7033 38206
rect 7119 38150 7175 38206
rect 7261 38150 7317 38206
rect 7403 38150 7459 38206
rect 7545 38150 7601 38206
rect 7687 38150 7743 38206
rect 7829 38150 7885 38206
rect 7971 38150 8027 38206
rect 8113 38150 8169 38206
rect 8255 38150 8311 38206
rect 8397 38150 8453 38206
rect 8539 38150 8595 38206
rect 8681 38150 8737 38206
rect 8823 38150 8879 38206
rect 8965 38150 9021 38206
rect 9107 38150 9163 38206
rect 9249 38150 9305 38206
rect 9391 38150 9447 38206
rect 9533 38150 9589 38206
rect 9675 38150 9731 38206
rect 9817 38150 9873 38206
rect 9959 38150 10015 38206
rect 10101 38150 10157 38206
rect 10243 38150 10299 38206
rect 10385 38150 10441 38206
rect 10527 38150 10583 38206
rect 10669 38150 10725 38206
rect 10811 38150 10867 38206
rect 10953 38150 11009 38206
rect 11095 38150 11151 38206
rect 11237 38150 11293 38206
rect 11379 38150 11435 38206
rect 11521 38150 11577 38206
rect 11663 38150 11719 38206
rect 11805 38150 11861 38206
rect 11947 38150 12003 38206
rect 12089 38150 12145 38206
rect 12231 38150 12287 38206
rect 12373 38150 12429 38206
rect 12515 38150 12571 38206
rect 12657 38150 12713 38206
rect 12799 38150 12855 38206
rect 12941 38150 12997 38206
rect 13083 38150 13139 38206
rect 13225 38150 13281 38206
rect 13367 38150 13423 38206
rect 13509 38150 13565 38206
rect 13651 38150 13707 38206
rect 13793 38150 13849 38206
rect 13935 38150 13991 38206
rect 14077 38150 14133 38206
rect 14219 38150 14275 38206
rect 14361 38150 14417 38206
rect 14503 38150 14559 38206
rect 14645 38150 14701 38206
rect 14787 38150 14843 38206
rect 161 38008 217 38064
rect 303 38008 359 38064
rect 445 38008 501 38064
rect 587 38008 643 38064
rect 729 38008 785 38064
rect 871 38008 927 38064
rect 1013 38008 1069 38064
rect 1155 38008 1211 38064
rect 1297 38008 1353 38064
rect 1439 38008 1495 38064
rect 1581 38008 1637 38064
rect 1723 38008 1779 38064
rect 1865 38008 1921 38064
rect 2007 38008 2063 38064
rect 2149 38008 2205 38064
rect 2291 38008 2347 38064
rect 2433 38008 2489 38064
rect 2575 38008 2631 38064
rect 2717 38008 2773 38064
rect 2859 38008 2915 38064
rect 3001 38008 3057 38064
rect 3143 38008 3199 38064
rect 3285 38008 3341 38064
rect 3427 38008 3483 38064
rect 3569 38008 3625 38064
rect 3711 38008 3767 38064
rect 3853 38008 3909 38064
rect 3995 38008 4051 38064
rect 4137 38008 4193 38064
rect 4279 38008 4335 38064
rect 4421 38008 4477 38064
rect 4563 38008 4619 38064
rect 4705 38008 4761 38064
rect 4847 38008 4903 38064
rect 4989 38008 5045 38064
rect 5131 38008 5187 38064
rect 5273 38008 5329 38064
rect 5415 38008 5471 38064
rect 5557 38008 5613 38064
rect 5699 38008 5755 38064
rect 5841 38008 5897 38064
rect 5983 38008 6039 38064
rect 6125 38008 6181 38064
rect 6267 38008 6323 38064
rect 6409 38008 6465 38064
rect 6551 38008 6607 38064
rect 6693 38008 6749 38064
rect 6835 38008 6891 38064
rect 6977 38008 7033 38064
rect 7119 38008 7175 38064
rect 7261 38008 7317 38064
rect 7403 38008 7459 38064
rect 7545 38008 7601 38064
rect 7687 38008 7743 38064
rect 7829 38008 7885 38064
rect 7971 38008 8027 38064
rect 8113 38008 8169 38064
rect 8255 38008 8311 38064
rect 8397 38008 8453 38064
rect 8539 38008 8595 38064
rect 8681 38008 8737 38064
rect 8823 38008 8879 38064
rect 8965 38008 9021 38064
rect 9107 38008 9163 38064
rect 9249 38008 9305 38064
rect 9391 38008 9447 38064
rect 9533 38008 9589 38064
rect 9675 38008 9731 38064
rect 9817 38008 9873 38064
rect 9959 38008 10015 38064
rect 10101 38008 10157 38064
rect 10243 38008 10299 38064
rect 10385 38008 10441 38064
rect 10527 38008 10583 38064
rect 10669 38008 10725 38064
rect 10811 38008 10867 38064
rect 10953 38008 11009 38064
rect 11095 38008 11151 38064
rect 11237 38008 11293 38064
rect 11379 38008 11435 38064
rect 11521 38008 11577 38064
rect 11663 38008 11719 38064
rect 11805 38008 11861 38064
rect 11947 38008 12003 38064
rect 12089 38008 12145 38064
rect 12231 38008 12287 38064
rect 12373 38008 12429 38064
rect 12515 38008 12571 38064
rect 12657 38008 12713 38064
rect 12799 38008 12855 38064
rect 12941 38008 12997 38064
rect 13083 38008 13139 38064
rect 13225 38008 13281 38064
rect 13367 38008 13423 38064
rect 13509 38008 13565 38064
rect 13651 38008 13707 38064
rect 13793 38008 13849 38064
rect 13935 38008 13991 38064
rect 14077 38008 14133 38064
rect 14219 38008 14275 38064
rect 14361 38008 14417 38064
rect 14503 38008 14559 38064
rect 14645 38008 14701 38064
rect 14787 38008 14843 38064
rect 161 37866 217 37922
rect 303 37866 359 37922
rect 445 37866 501 37922
rect 587 37866 643 37922
rect 729 37866 785 37922
rect 871 37866 927 37922
rect 1013 37866 1069 37922
rect 1155 37866 1211 37922
rect 1297 37866 1353 37922
rect 1439 37866 1495 37922
rect 1581 37866 1637 37922
rect 1723 37866 1779 37922
rect 1865 37866 1921 37922
rect 2007 37866 2063 37922
rect 2149 37866 2205 37922
rect 2291 37866 2347 37922
rect 2433 37866 2489 37922
rect 2575 37866 2631 37922
rect 2717 37866 2773 37922
rect 2859 37866 2915 37922
rect 3001 37866 3057 37922
rect 3143 37866 3199 37922
rect 3285 37866 3341 37922
rect 3427 37866 3483 37922
rect 3569 37866 3625 37922
rect 3711 37866 3767 37922
rect 3853 37866 3909 37922
rect 3995 37866 4051 37922
rect 4137 37866 4193 37922
rect 4279 37866 4335 37922
rect 4421 37866 4477 37922
rect 4563 37866 4619 37922
rect 4705 37866 4761 37922
rect 4847 37866 4903 37922
rect 4989 37866 5045 37922
rect 5131 37866 5187 37922
rect 5273 37866 5329 37922
rect 5415 37866 5471 37922
rect 5557 37866 5613 37922
rect 5699 37866 5755 37922
rect 5841 37866 5897 37922
rect 5983 37866 6039 37922
rect 6125 37866 6181 37922
rect 6267 37866 6323 37922
rect 6409 37866 6465 37922
rect 6551 37866 6607 37922
rect 6693 37866 6749 37922
rect 6835 37866 6891 37922
rect 6977 37866 7033 37922
rect 7119 37866 7175 37922
rect 7261 37866 7317 37922
rect 7403 37866 7459 37922
rect 7545 37866 7601 37922
rect 7687 37866 7743 37922
rect 7829 37866 7885 37922
rect 7971 37866 8027 37922
rect 8113 37866 8169 37922
rect 8255 37866 8311 37922
rect 8397 37866 8453 37922
rect 8539 37866 8595 37922
rect 8681 37866 8737 37922
rect 8823 37866 8879 37922
rect 8965 37866 9021 37922
rect 9107 37866 9163 37922
rect 9249 37866 9305 37922
rect 9391 37866 9447 37922
rect 9533 37866 9589 37922
rect 9675 37866 9731 37922
rect 9817 37866 9873 37922
rect 9959 37866 10015 37922
rect 10101 37866 10157 37922
rect 10243 37866 10299 37922
rect 10385 37866 10441 37922
rect 10527 37866 10583 37922
rect 10669 37866 10725 37922
rect 10811 37866 10867 37922
rect 10953 37866 11009 37922
rect 11095 37866 11151 37922
rect 11237 37866 11293 37922
rect 11379 37866 11435 37922
rect 11521 37866 11577 37922
rect 11663 37866 11719 37922
rect 11805 37866 11861 37922
rect 11947 37866 12003 37922
rect 12089 37866 12145 37922
rect 12231 37866 12287 37922
rect 12373 37866 12429 37922
rect 12515 37866 12571 37922
rect 12657 37866 12713 37922
rect 12799 37866 12855 37922
rect 12941 37866 12997 37922
rect 13083 37866 13139 37922
rect 13225 37866 13281 37922
rect 13367 37866 13423 37922
rect 13509 37866 13565 37922
rect 13651 37866 13707 37922
rect 13793 37866 13849 37922
rect 13935 37866 13991 37922
rect 14077 37866 14133 37922
rect 14219 37866 14275 37922
rect 14361 37866 14417 37922
rect 14503 37866 14559 37922
rect 14645 37866 14701 37922
rect 14787 37866 14843 37922
rect 161 37724 217 37780
rect 303 37724 359 37780
rect 445 37724 501 37780
rect 587 37724 643 37780
rect 729 37724 785 37780
rect 871 37724 927 37780
rect 1013 37724 1069 37780
rect 1155 37724 1211 37780
rect 1297 37724 1353 37780
rect 1439 37724 1495 37780
rect 1581 37724 1637 37780
rect 1723 37724 1779 37780
rect 1865 37724 1921 37780
rect 2007 37724 2063 37780
rect 2149 37724 2205 37780
rect 2291 37724 2347 37780
rect 2433 37724 2489 37780
rect 2575 37724 2631 37780
rect 2717 37724 2773 37780
rect 2859 37724 2915 37780
rect 3001 37724 3057 37780
rect 3143 37724 3199 37780
rect 3285 37724 3341 37780
rect 3427 37724 3483 37780
rect 3569 37724 3625 37780
rect 3711 37724 3767 37780
rect 3853 37724 3909 37780
rect 3995 37724 4051 37780
rect 4137 37724 4193 37780
rect 4279 37724 4335 37780
rect 4421 37724 4477 37780
rect 4563 37724 4619 37780
rect 4705 37724 4761 37780
rect 4847 37724 4903 37780
rect 4989 37724 5045 37780
rect 5131 37724 5187 37780
rect 5273 37724 5329 37780
rect 5415 37724 5471 37780
rect 5557 37724 5613 37780
rect 5699 37724 5755 37780
rect 5841 37724 5897 37780
rect 5983 37724 6039 37780
rect 6125 37724 6181 37780
rect 6267 37724 6323 37780
rect 6409 37724 6465 37780
rect 6551 37724 6607 37780
rect 6693 37724 6749 37780
rect 6835 37724 6891 37780
rect 6977 37724 7033 37780
rect 7119 37724 7175 37780
rect 7261 37724 7317 37780
rect 7403 37724 7459 37780
rect 7545 37724 7601 37780
rect 7687 37724 7743 37780
rect 7829 37724 7885 37780
rect 7971 37724 8027 37780
rect 8113 37724 8169 37780
rect 8255 37724 8311 37780
rect 8397 37724 8453 37780
rect 8539 37724 8595 37780
rect 8681 37724 8737 37780
rect 8823 37724 8879 37780
rect 8965 37724 9021 37780
rect 9107 37724 9163 37780
rect 9249 37724 9305 37780
rect 9391 37724 9447 37780
rect 9533 37724 9589 37780
rect 9675 37724 9731 37780
rect 9817 37724 9873 37780
rect 9959 37724 10015 37780
rect 10101 37724 10157 37780
rect 10243 37724 10299 37780
rect 10385 37724 10441 37780
rect 10527 37724 10583 37780
rect 10669 37724 10725 37780
rect 10811 37724 10867 37780
rect 10953 37724 11009 37780
rect 11095 37724 11151 37780
rect 11237 37724 11293 37780
rect 11379 37724 11435 37780
rect 11521 37724 11577 37780
rect 11663 37724 11719 37780
rect 11805 37724 11861 37780
rect 11947 37724 12003 37780
rect 12089 37724 12145 37780
rect 12231 37724 12287 37780
rect 12373 37724 12429 37780
rect 12515 37724 12571 37780
rect 12657 37724 12713 37780
rect 12799 37724 12855 37780
rect 12941 37724 12997 37780
rect 13083 37724 13139 37780
rect 13225 37724 13281 37780
rect 13367 37724 13423 37780
rect 13509 37724 13565 37780
rect 13651 37724 13707 37780
rect 13793 37724 13849 37780
rect 13935 37724 13991 37780
rect 14077 37724 14133 37780
rect 14219 37724 14275 37780
rect 14361 37724 14417 37780
rect 14503 37724 14559 37780
rect 14645 37724 14701 37780
rect 14787 37724 14843 37780
rect 161 37582 217 37638
rect 303 37582 359 37638
rect 445 37582 501 37638
rect 587 37582 643 37638
rect 729 37582 785 37638
rect 871 37582 927 37638
rect 1013 37582 1069 37638
rect 1155 37582 1211 37638
rect 1297 37582 1353 37638
rect 1439 37582 1495 37638
rect 1581 37582 1637 37638
rect 1723 37582 1779 37638
rect 1865 37582 1921 37638
rect 2007 37582 2063 37638
rect 2149 37582 2205 37638
rect 2291 37582 2347 37638
rect 2433 37582 2489 37638
rect 2575 37582 2631 37638
rect 2717 37582 2773 37638
rect 2859 37582 2915 37638
rect 3001 37582 3057 37638
rect 3143 37582 3199 37638
rect 3285 37582 3341 37638
rect 3427 37582 3483 37638
rect 3569 37582 3625 37638
rect 3711 37582 3767 37638
rect 3853 37582 3909 37638
rect 3995 37582 4051 37638
rect 4137 37582 4193 37638
rect 4279 37582 4335 37638
rect 4421 37582 4477 37638
rect 4563 37582 4619 37638
rect 4705 37582 4761 37638
rect 4847 37582 4903 37638
rect 4989 37582 5045 37638
rect 5131 37582 5187 37638
rect 5273 37582 5329 37638
rect 5415 37582 5471 37638
rect 5557 37582 5613 37638
rect 5699 37582 5755 37638
rect 5841 37582 5897 37638
rect 5983 37582 6039 37638
rect 6125 37582 6181 37638
rect 6267 37582 6323 37638
rect 6409 37582 6465 37638
rect 6551 37582 6607 37638
rect 6693 37582 6749 37638
rect 6835 37582 6891 37638
rect 6977 37582 7033 37638
rect 7119 37582 7175 37638
rect 7261 37582 7317 37638
rect 7403 37582 7459 37638
rect 7545 37582 7601 37638
rect 7687 37582 7743 37638
rect 7829 37582 7885 37638
rect 7971 37582 8027 37638
rect 8113 37582 8169 37638
rect 8255 37582 8311 37638
rect 8397 37582 8453 37638
rect 8539 37582 8595 37638
rect 8681 37582 8737 37638
rect 8823 37582 8879 37638
rect 8965 37582 9021 37638
rect 9107 37582 9163 37638
rect 9249 37582 9305 37638
rect 9391 37582 9447 37638
rect 9533 37582 9589 37638
rect 9675 37582 9731 37638
rect 9817 37582 9873 37638
rect 9959 37582 10015 37638
rect 10101 37582 10157 37638
rect 10243 37582 10299 37638
rect 10385 37582 10441 37638
rect 10527 37582 10583 37638
rect 10669 37582 10725 37638
rect 10811 37582 10867 37638
rect 10953 37582 11009 37638
rect 11095 37582 11151 37638
rect 11237 37582 11293 37638
rect 11379 37582 11435 37638
rect 11521 37582 11577 37638
rect 11663 37582 11719 37638
rect 11805 37582 11861 37638
rect 11947 37582 12003 37638
rect 12089 37582 12145 37638
rect 12231 37582 12287 37638
rect 12373 37582 12429 37638
rect 12515 37582 12571 37638
rect 12657 37582 12713 37638
rect 12799 37582 12855 37638
rect 12941 37582 12997 37638
rect 13083 37582 13139 37638
rect 13225 37582 13281 37638
rect 13367 37582 13423 37638
rect 13509 37582 13565 37638
rect 13651 37582 13707 37638
rect 13793 37582 13849 37638
rect 13935 37582 13991 37638
rect 14077 37582 14133 37638
rect 14219 37582 14275 37638
rect 14361 37582 14417 37638
rect 14503 37582 14559 37638
rect 14645 37582 14701 37638
rect 14787 37582 14843 37638
rect 161 37440 217 37496
rect 303 37440 359 37496
rect 445 37440 501 37496
rect 587 37440 643 37496
rect 729 37440 785 37496
rect 871 37440 927 37496
rect 1013 37440 1069 37496
rect 1155 37440 1211 37496
rect 1297 37440 1353 37496
rect 1439 37440 1495 37496
rect 1581 37440 1637 37496
rect 1723 37440 1779 37496
rect 1865 37440 1921 37496
rect 2007 37440 2063 37496
rect 2149 37440 2205 37496
rect 2291 37440 2347 37496
rect 2433 37440 2489 37496
rect 2575 37440 2631 37496
rect 2717 37440 2773 37496
rect 2859 37440 2915 37496
rect 3001 37440 3057 37496
rect 3143 37440 3199 37496
rect 3285 37440 3341 37496
rect 3427 37440 3483 37496
rect 3569 37440 3625 37496
rect 3711 37440 3767 37496
rect 3853 37440 3909 37496
rect 3995 37440 4051 37496
rect 4137 37440 4193 37496
rect 4279 37440 4335 37496
rect 4421 37440 4477 37496
rect 4563 37440 4619 37496
rect 4705 37440 4761 37496
rect 4847 37440 4903 37496
rect 4989 37440 5045 37496
rect 5131 37440 5187 37496
rect 5273 37440 5329 37496
rect 5415 37440 5471 37496
rect 5557 37440 5613 37496
rect 5699 37440 5755 37496
rect 5841 37440 5897 37496
rect 5983 37440 6039 37496
rect 6125 37440 6181 37496
rect 6267 37440 6323 37496
rect 6409 37440 6465 37496
rect 6551 37440 6607 37496
rect 6693 37440 6749 37496
rect 6835 37440 6891 37496
rect 6977 37440 7033 37496
rect 7119 37440 7175 37496
rect 7261 37440 7317 37496
rect 7403 37440 7459 37496
rect 7545 37440 7601 37496
rect 7687 37440 7743 37496
rect 7829 37440 7885 37496
rect 7971 37440 8027 37496
rect 8113 37440 8169 37496
rect 8255 37440 8311 37496
rect 8397 37440 8453 37496
rect 8539 37440 8595 37496
rect 8681 37440 8737 37496
rect 8823 37440 8879 37496
rect 8965 37440 9021 37496
rect 9107 37440 9163 37496
rect 9249 37440 9305 37496
rect 9391 37440 9447 37496
rect 9533 37440 9589 37496
rect 9675 37440 9731 37496
rect 9817 37440 9873 37496
rect 9959 37440 10015 37496
rect 10101 37440 10157 37496
rect 10243 37440 10299 37496
rect 10385 37440 10441 37496
rect 10527 37440 10583 37496
rect 10669 37440 10725 37496
rect 10811 37440 10867 37496
rect 10953 37440 11009 37496
rect 11095 37440 11151 37496
rect 11237 37440 11293 37496
rect 11379 37440 11435 37496
rect 11521 37440 11577 37496
rect 11663 37440 11719 37496
rect 11805 37440 11861 37496
rect 11947 37440 12003 37496
rect 12089 37440 12145 37496
rect 12231 37440 12287 37496
rect 12373 37440 12429 37496
rect 12515 37440 12571 37496
rect 12657 37440 12713 37496
rect 12799 37440 12855 37496
rect 12941 37440 12997 37496
rect 13083 37440 13139 37496
rect 13225 37440 13281 37496
rect 13367 37440 13423 37496
rect 13509 37440 13565 37496
rect 13651 37440 13707 37496
rect 13793 37440 13849 37496
rect 13935 37440 13991 37496
rect 14077 37440 14133 37496
rect 14219 37440 14275 37496
rect 14361 37440 14417 37496
rect 14503 37440 14559 37496
rect 14645 37440 14701 37496
rect 14787 37440 14843 37496
rect 161 37298 217 37354
rect 303 37298 359 37354
rect 445 37298 501 37354
rect 587 37298 643 37354
rect 729 37298 785 37354
rect 871 37298 927 37354
rect 1013 37298 1069 37354
rect 1155 37298 1211 37354
rect 1297 37298 1353 37354
rect 1439 37298 1495 37354
rect 1581 37298 1637 37354
rect 1723 37298 1779 37354
rect 1865 37298 1921 37354
rect 2007 37298 2063 37354
rect 2149 37298 2205 37354
rect 2291 37298 2347 37354
rect 2433 37298 2489 37354
rect 2575 37298 2631 37354
rect 2717 37298 2773 37354
rect 2859 37298 2915 37354
rect 3001 37298 3057 37354
rect 3143 37298 3199 37354
rect 3285 37298 3341 37354
rect 3427 37298 3483 37354
rect 3569 37298 3625 37354
rect 3711 37298 3767 37354
rect 3853 37298 3909 37354
rect 3995 37298 4051 37354
rect 4137 37298 4193 37354
rect 4279 37298 4335 37354
rect 4421 37298 4477 37354
rect 4563 37298 4619 37354
rect 4705 37298 4761 37354
rect 4847 37298 4903 37354
rect 4989 37298 5045 37354
rect 5131 37298 5187 37354
rect 5273 37298 5329 37354
rect 5415 37298 5471 37354
rect 5557 37298 5613 37354
rect 5699 37298 5755 37354
rect 5841 37298 5897 37354
rect 5983 37298 6039 37354
rect 6125 37298 6181 37354
rect 6267 37298 6323 37354
rect 6409 37298 6465 37354
rect 6551 37298 6607 37354
rect 6693 37298 6749 37354
rect 6835 37298 6891 37354
rect 6977 37298 7033 37354
rect 7119 37298 7175 37354
rect 7261 37298 7317 37354
rect 7403 37298 7459 37354
rect 7545 37298 7601 37354
rect 7687 37298 7743 37354
rect 7829 37298 7885 37354
rect 7971 37298 8027 37354
rect 8113 37298 8169 37354
rect 8255 37298 8311 37354
rect 8397 37298 8453 37354
rect 8539 37298 8595 37354
rect 8681 37298 8737 37354
rect 8823 37298 8879 37354
rect 8965 37298 9021 37354
rect 9107 37298 9163 37354
rect 9249 37298 9305 37354
rect 9391 37298 9447 37354
rect 9533 37298 9589 37354
rect 9675 37298 9731 37354
rect 9817 37298 9873 37354
rect 9959 37298 10015 37354
rect 10101 37298 10157 37354
rect 10243 37298 10299 37354
rect 10385 37298 10441 37354
rect 10527 37298 10583 37354
rect 10669 37298 10725 37354
rect 10811 37298 10867 37354
rect 10953 37298 11009 37354
rect 11095 37298 11151 37354
rect 11237 37298 11293 37354
rect 11379 37298 11435 37354
rect 11521 37298 11577 37354
rect 11663 37298 11719 37354
rect 11805 37298 11861 37354
rect 11947 37298 12003 37354
rect 12089 37298 12145 37354
rect 12231 37298 12287 37354
rect 12373 37298 12429 37354
rect 12515 37298 12571 37354
rect 12657 37298 12713 37354
rect 12799 37298 12855 37354
rect 12941 37298 12997 37354
rect 13083 37298 13139 37354
rect 13225 37298 13281 37354
rect 13367 37298 13423 37354
rect 13509 37298 13565 37354
rect 13651 37298 13707 37354
rect 13793 37298 13849 37354
rect 13935 37298 13991 37354
rect 14077 37298 14133 37354
rect 14219 37298 14275 37354
rect 14361 37298 14417 37354
rect 14503 37298 14559 37354
rect 14645 37298 14701 37354
rect 14787 37298 14843 37354
rect 161 37156 217 37212
rect 303 37156 359 37212
rect 445 37156 501 37212
rect 587 37156 643 37212
rect 729 37156 785 37212
rect 871 37156 927 37212
rect 1013 37156 1069 37212
rect 1155 37156 1211 37212
rect 1297 37156 1353 37212
rect 1439 37156 1495 37212
rect 1581 37156 1637 37212
rect 1723 37156 1779 37212
rect 1865 37156 1921 37212
rect 2007 37156 2063 37212
rect 2149 37156 2205 37212
rect 2291 37156 2347 37212
rect 2433 37156 2489 37212
rect 2575 37156 2631 37212
rect 2717 37156 2773 37212
rect 2859 37156 2915 37212
rect 3001 37156 3057 37212
rect 3143 37156 3199 37212
rect 3285 37156 3341 37212
rect 3427 37156 3483 37212
rect 3569 37156 3625 37212
rect 3711 37156 3767 37212
rect 3853 37156 3909 37212
rect 3995 37156 4051 37212
rect 4137 37156 4193 37212
rect 4279 37156 4335 37212
rect 4421 37156 4477 37212
rect 4563 37156 4619 37212
rect 4705 37156 4761 37212
rect 4847 37156 4903 37212
rect 4989 37156 5045 37212
rect 5131 37156 5187 37212
rect 5273 37156 5329 37212
rect 5415 37156 5471 37212
rect 5557 37156 5613 37212
rect 5699 37156 5755 37212
rect 5841 37156 5897 37212
rect 5983 37156 6039 37212
rect 6125 37156 6181 37212
rect 6267 37156 6323 37212
rect 6409 37156 6465 37212
rect 6551 37156 6607 37212
rect 6693 37156 6749 37212
rect 6835 37156 6891 37212
rect 6977 37156 7033 37212
rect 7119 37156 7175 37212
rect 7261 37156 7317 37212
rect 7403 37156 7459 37212
rect 7545 37156 7601 37212
rect 7687 37156 7743 37212
rect 7829 37156 7885 37212
rect 7971 37156 8027 37212
rect 8113 37156 8169 37212
rect 8255 37156 8311 37212
rect 8397 37156 8453 37212
rect 8539 37156 8595 37212
rect 8681 37156 8737 37212
rect 8823 37156 8879 37212
rect 8965 37156 9021 37212
rect 9107 37156 9163 37212
rect 9249 37156 9305 37212
rect 9391 37156 9447 37212
rect 9533 37156 9589 37212
rect 9675 37156 9731 37212
rect 9817 37156 9873 37212
rect 9959 37156 10015 37212
rect 10101 37156 10157 37212
rect 10243 37156 10299 37212
rect 10385 37156 10441 37212
rect 10527 37156 10583 37212
rect 10669 37156 10725 37212
rect 10811 37156 10867 37212
rect 10953 37156 11009 37212
rect 11095 37156 11151 37212
rect 11237 37156 11293 37212
rect 11379 37156 11435 37212
rect 11521 37156 11577 37212
rect 11663 37156 11719 37212
rect 11805 37156 11861 37212
rect 11947 37156 12003 37212
rect 12089 37156 12145 37212
rect 12231 37156 12287 37212
rect 12373 37156 12429 37212
rect 12515 37156 12571 37212
rect 12657 37156 12713 37212
rect 12799 37156 12855 37212
rect 12941 37156 12997 37212
rect 13083 37156 13139 37212
rect 13225 37156 13281 37212
rect 13367 37156 13423 37212
rect 13509 37156 13565 37212
rect 13651 37156 13707 37212
rect 13793 37156 13849 37212
rect 13935 37156 13991 37212
rect 14077 37156 14133 37212
rect 14219 37156 14275 37212
rect 14361 37156 14417 37212
rect 14503 37156 14559 37212
rect 14645 37156 14701 37212
rect 14787 37156 14843 37212
rect 161 37014 217 37070
rect 303 37014 359 37070
rect 445 37014 501 37070
rect 587 37014 643 37070
rect 729 37014 785 37070
rect 871 37014 927 37070
rect 1013 37014 1069 37070
rect 1155 37014 1211 37070
rect 1297 37014 1353 37070
rect 1439 37014 1495 37070
rect 1581 37014 1637 37070
rect 1723 37014 1779 37070
rect 1865 37014 1921 37070
rect 2007 37014 2063 37070
rect 2149 37014 2205 37070
rect 2291 37014 2347 37070
rect 2433 37014 2489 37070
rect 2575 37014 2631 37070
rect 2717 37014 2773 37070
rect 2859 37014 2915 37070
rect 3001 37014 3057 37070
rect 3143 37014 3199 37070
rect 3285 37014 3341 37070
rect 3427 37014 3483 37070
rect 3569 37014 3625 37070
rect 3711 37014 3767 37070
rect 3853 37014 3909 37070
rect 3995 37014 4051 37070
rect 4137 37014 4193 37070
rect 4279 37014 4335 37070
rect 4421 37014 4477 37070
rect 4563 37014 4619 37070
rect 4705 37014 4761 37070
rect 4847 37014 4903 37070
rect 4989 37014 5045 37070
rect 5131 37014 5187 37070
rect 5273 37014 5329 37070
rect 5415 37014 5471 37070
rect 5557 37014 5613 37070
rect 5699 37014 5755 37070
rect 5841 37014 5897 37070
rect 5983 37014 6039 37070
rect 6125 37014 6181 37070
rect 6267 37014 6323 37070
rect 6409 37014 6465 37070
rect 6551 37014 6607 37070
rect 6693 37014 6749 37070
rect 6835 37014 6891 37070
rect 6977 37014 7033 37070
rect 7119 37014 7175 37070
rect 7261 37014 7317 37070
rect 7403 37014 7459 37070
rect 7545 37014 7601 37070
rect 7687 37014 7743 37070
rect 7829 37014 7885 37070
rect 7971 37014 8027 37070
rect 8113 37014 8169 37070
rect 8255 37014 8311 37070
rect 8397 37014 8453 37070
rect 8539 37014 8595 37070
rect 8681 37014 8737 37070
rect 8823 37014 8879 37070
rect 8965 37014 9021 37070
rect 9107 37014 9163 37070
rect 9249 37014 9305 37070
rect 9391 37014 9447 37070
rect 9533 37014 9589 37070
rect 9675 37014 9731 37070
rect 9817 37014 9873 37070
rect 9959 37014 10015 37070
rect 10101 37014 10157 37070
rect 10243 37014 10299 37070
rect 10385 37014 10441 37070
rect 10527 37014 10583 37070
rect 10669 37014 10725 37070
rect 10811 37014 10867 37070
rect 10953 37014 11009 37070
rect 11095 37014 11151 37070
rect 11237 37014 11293 37070
rect 11379 37014 11435 37070
rect 11521 37014 11577 37070
rect 11663 37014 11719 37070
rect 11805 37014 11861 37070
rect 11947 37014 12003 37070
rect 12089 37014 12145 37070
rect 12231 37014 12287 37070
rect 12373 37014 12429 37070
rect 12515 37014 12571 37070
rect 12657 37014 12713 37070
rect 12799 37014 12855 37070
rect 12941 37014 12997 37070
rect 13083 37014 13139 37070
rect 13225 37014 13281 37070
rect 13367 37014 13423 37070
rect 13509 37014 13565 37070
rect 13651 37014 13707 37070
rect 13793 37014 13849 37070
rect 13935 37014 13991 37070
rect 14077 37014 14133 37070
rect 14219 37014 14275 37070
rect 14361 37014 14417 37070
rect 14503 37014 14559 37070
rect 14645 37014 14701 37070
rect 14787 37014 14843 37070
rect 161 36872 217 36928
rect 303 36872 359 36928
rect 445 36872 501 36928
rect 587 36872 643 36928
rect 729 36872 785 36928
rect 871 36872 927 36928
rect 1013 36872 1069 36928
rect 1155 36872 1211 36928
rect 1297 36872 1353 36928
rect 1439 36872 1495 36928
rect 1581 36872 1637 36928
rect 1723 36872 1779 36928
rect 1865 36872 1921 36928
rect 2007 36872 2063 36928
rect 2149 36872 2205 36928
rect 2291 36872 2347 36928
rect 2433 36872 2489 36928
rect 2575 36872 2631 36928
rect 2717 36872 2773 36928
rect 2859 36872 2915 36928
rect 3001 36872 3057 36928
rect 3143 36872 3199 36928
rect 3285 36872 3341 36928
rect 3427 36872 3483 36928
rect 3569 36872 3625 36928
rect 3711 36872 3767 36928
rect 3853 36872 3909 36928
rect 3995 36872 4051 36928
rect 4137 36872 4193 36928
rect 4279 36872 4335 36928
rect 4421 36872 4477 36928
rect 4563 36872 4619 36928
rect 4705 36872 4761 36928
rect 4847 36872 4903 36928
rect 4989 36872 5045 36928
rect 5131 36872 5187 36928
rect 5273 36872 5329 36928
rect 5415 36872 5471 36928
rect 5557 36872 5613 36928
rect 5699 36872 5755 36928
rect 5841 36872 5897 36928
rect 5983 36872 6039 36928
rect 6125 36872 6181 36928
rect 6267 36872 6323 36928
rect 6409 36872 6465 36928
rect 6551 36872 6607 36928
rect 6693 36872 6749 36928
rect 6835 36872 6891 36928
rect 6977 36872 7033 36928
rect 7119 36872 7175 36928
rect 7261 36872 7317 36928
rect 7403 36872 7459 36928
rect 7545 36872 7601 36928
rect 7687 36872 7743 36928
rect 7829 36872 7885 36928
rect 7971 36872 8027 36928
rect 8113 36872 8169 36928
rect 8255 36872 8311 36928
rect 8397 36872 8453 36928
rect 8539 36872 8595 36928
rect 8681 36872 8737 36928
rect 8823 36872 8879 36928
rect 8965 36872 9021 36928
rect 9107 36872 9163 36928
rect 9249 36872 9305 36928
rect 9391 36872 9447 36928
rect 9533 36872 9589 36928
rect 9675 36872 9731 36928
rect 9817 36872 9873 36928
rect 9959 36872 10015 36928
rect 10101 36872 10157 36928
rect 10243 36872 10299 36928
rect 10385 36872 10441 36928
rect 10527 36872 10583 36928
rect 10669 36872 10725 36928
rect 10811 36872 10867 36928
rect 10953 36872 11009 36928
rect 11095 36872 11151 36928
rect 11237 36872 11293 36928
rect 11379 36872 11435 36928
rect 11521 36872 11577 36928
rect 11663 36872 11719 36928
rect 11805 36872 11861 36928
rect 11947 36872 12003 36928
rect 12089 36872 12145 36928
rect 12231 36872 12287 36928
rect 12373 36872 12429 36928
rect 12515 36872 12571 36928
rect 12657 36872 12713 36928
rect 12799 36872 12855 36928
rect 12941 36872 12997 36928
rect 13083 36872 13139 36928
rect 13225 36872 13281 36928
rect 13367 36872 13423 36928
rect 13509 36872 13565 36928
rect 13651 36872 13707 36928
rect 13793 36872 13849 36928
rect 13935 36872 13991 36928
rect 14077 36872 14133 36928
rect 14219 36872 14275 36928
rect 14361 36872 14417 36928
rect 14503 36872 14559 36928
rect 14645 36872 14701 36928
rect 14787 36872 14843 36928
rect 161 36730 217 36786
rect 303 36730 359 36786
rect 445 36730 501 36786
rect 587 36730 643 36786
rect 729 36730 785 36786
rect 871 36730 927 36786
rect 1013 36730 1069 36786
rect 1155 36730 1211 36786
rect 1297 36730 1353 36786
rect 1439 36730 1495 36786
rect 1581 36730 1637 36786
rect 1723 36730 1779 36786
rect 1865 36730 1921 36786
rect 2007 36730 2063 36786
rect 2149 36730 2205 36786
rect 2291 36730 2347 36786
rect 2433 36730 2489 36786
rect 2575 36730 2631 36786
rect 2717 36730 2773 36786
rect 2859 36730 2915 36786
rect 3001 36730 3057 36786
rect 3143 36730 3199 36786
rect 3285 36730 3341 36786
rect 3427 36730 3483 36786
rect 3569 36730 3625 36786
rect 3711 36730 3767 36786
rect 3853 36730 3909 36786
rect 3995 36730 4051 36786
rect 4137 36730 4193 36786
rect 4279 36730 4335 36786
rect 4421 36730 4477 36786
rect 4563 36730 4619 36786
rect 4705 36730 4761 36786
rect 4847 36730 4903 36786
rect 4989 36730 5045 36786
rect 5131 36730 5187 36786
rect 5273 36730 5329 36786
rect 5415 36730 5471 36786
rect 5557 36730 5613 36786
rect 5699 36730 5755 36786
rect 5841 36730 5897 36786
rect 5983 36730 6039 36786
rect 6125 36730 6181 36786
rect 6267 36730 6323 36786
rect 6409 36730 6465 36786
rect 6551 36730 6607 36786
rect 6693 36730 6749 36786
rect 6835 36730 6891 36786
rect 6977 36730 7033 36786
rect 7119 36730 7175 36786
rect 7261 36730 7317 36786
rect 7403 36730 7459 36786
rect 7545 36730 7601 36786
rect 7687 36730 7743 36786
rect 7829 36730 7885 36786
rect 7971 36730 8027 36786
rect 8113 36730 8169 36786
rect 8255 36730 8311 36786
rect 8397 36730 8453 36786
rect 8539 36730 8595 36786
rect 8681 36730 8737 36786
rect 8823 36730 8879 36786
rect 8965 36730 9021 36786
rect 9107 36730 9163 36786
rect 9249 36730 9305 36786
rect 9391 36730 9447 36786
rect 9533 36730 9589 36786
rect 9675 36730 9731 36786
rect 9817 36730 9873 36786
rect 9959 36730 10015 36786
rect 10101 36730 10157 36786
rect 10243 36730 10299 36786
rect 10385 36730 10441 36786
rect 10527 36730 10583 36786
rect 10669 36730 10725 36786
rect 10811 36730 10867 36786
rect 10953 36730 11009 36786
rect 11095 36730 11151 36786
rect 11237 36730 11293 36786
rect 11379 36730 11435 36786
rect 11521 36730 11577 36786
rect 11663 36730 11719 36786
rect 11805 36730 11861 36786
rect 11947 36730 12003 36786
rect 12089 36730 12145 36786
rect 12231 36730 12287 36786
rect 12373 36730 12429 36786
rect 12515 36730 12571 36786
rect 12657 36730 12713 36786
rect 12799 36730 12855 36786
rect 12941 36730 12997 36786
rect 13083 36730 13139 36786
rect 13225 36730 13281 36786
rect 13367 36730 13423 36786
rect 13509 36730 13565 36786
rect 13651 36730 13707 36786
rect 13793 36730 13849 36786
rect 13935 36730 13991 36786
rect 14077 36730 14133 36786
rect 14219 36730 14275 36786
rect 14361 36730 14417 36786
rect 14503 36730 14559 36786
rect 14645 36730 14701 36786
rect 14787 36730 14843 36786
rect 161 36588 217 36644
rect 303 36588 359 36644
rect 445 36588 501 36644
rect 587 36588 643 36644
rect 729 36588 785 36644
rect 871 36588 927 36644
rect 1013 36588 1069 36644
rect 1155 36588 1211 36644
rect 1297 36588 1353 36644
rect 1439 36588 1495 36644
rect 1581 36588 1637 36644
rect 1723 36588 1779 36644
rect 1865 36588 1921 36644
rect 2007 36588 2063 36644
rect 2149 36588 2205 36644
rect 2291 36588 2347 36644
rect 2433 36588 2489 36644
rect 2575 36588 2631 36644
rect 2717 36588 2773 36644
rect 2859 36588 2915 36644
rect 3001 36588 3057 36644
rect 3143 36588 3199 36644
rect 3285 36588 3341 36644
rect 3427 36588 3483 36644
rect 3569 36588 3625 36644
rect 3711 36588 3767 36644
rect 3853 36588 3909 36644
rect 3995 36588 4051 36644
rect 4137 36588 4193 36644
rect 4279 36588 4335 36644
rect 4421 36588 4477 36644
rect 4563 36588 4619 36644
rect 4705 36588 4761 36644
rect 4847 36588 4903 36644
rect 4989 36588 5045 36644
rect 5131 36588 5187 36644
rect 5273 36588 5329 36644
rect 5415 36588 5471 36644
rect 5557 36588 5613 36644
rect 5699 36588 5755 36644
rect 5841 36588 5897 36644
rect 5983 36588 6039 36644
rect 6125 36588 6181 36644
rect 6267 36588 6323 36644
rect 6409 36588 6465 36644
rect 6551 36588 6607 36644
rect 6693 36588 6749 36644
rect 6835 36588 6891 36644
rect 6977 36588 7033 36644
rect 7119 36588 7175 36644
rect 7261 36588 7317 36644
rect 7403 36588 7459 36644
rect 7545 36588 7601 36644
rect 7687 36588 7743 36644
rect 7829 36588 7885 36644
rect 7971 36588 8027 36644
rect 8113 36588 8169 36644
rect 8255 36588 8311 36644
rect 8397 36588 8453 36644
rect 8539 36588 8595 36644
rect 8681 36588 8737 36644
rect 8823 36588 8879 36644
rect 8965 36588 9021 36644
rect 9107 36588 9163 36644
rect 9249 36588 9305 36644
rect 9391 36588 9447 36644
rect 9533 36588 9589 36644
rect 9675 36588 9731 36644
rect 9817 36588 9873 36644
rect 9959 36588 10015 36644
rect 10101 36588 10157 36644
rect 10243 36588 10299 36644
rect 10385 36588 10441 36644
rect 10527 36588 10583 36644
rect 10669 36588 10725 36644
rect 10811 36588 10867 36644
rect 10953 36588 11009 36644
rect 11095 36588 11151 36644
rect 11237 36588 11293 36644
rect 11379 36588 11435 36644
rect 11521 36588 11577 36644
rect 11663 36588 11719 36644
rect 11805 36588 11861 36644
rect 11947 36588 12003 36644
rect 12089 36588 12145 36644
rect 12231 36588 12287 36644
rect 12373 36588 12429 36644
rect 12515 36588 12571 36644
rect 12657 36588 12713 36644
rect 12799 36588 12855 36644
rect 12941 36588 12997 36644
rect 13083 36588 13139 36644
rect 13225 36588 13281 36644
rect 13367 36588 13423 36644
rect 13509 36588 13565 36644
rect 13651 36588 13707 36644
rect 13793 36588 13849 36644
rect 13935 36588 13991 36644
rect 14077 36588 14133 36644
rect 14219 36588 14275 36644
rect 14361 36588 14417 36644
rect 14503 36588 14559 36644
rect 14645 36588 14701 36644
rect 14787 36588 14843 36644
rect 161 36446 217 36502
rect 303 36446 359 36502
rect 445 36446 501 36502
rect 587 36446 643 36502
rect 729 36446 785 36502
rect 871 36446 927 36502
rect 1013 36446 1069 36502
rect 1155 36446 1211 36502
rect 1297 36446 1353 36502
rect 1439 36446 1495 36502
rect 1581 36446 1637 36502
rect 1723 36446 1779 36502
rect 1865 36446 1921 36502
rect 2007 36446 2063 36502
rect 2149 36446 2205 36502
rect 2291 36446 2347 36502
rect 2433 36446 2489 36502
rect 2575 36446 2631 36502
rect 2717 36446 2773 36502
rect 2859 36446 2915 36502
rect 3001 36446 3057 36502
rect 3143 36446 3199 36502
rect 3285 36446 3341 36502
rect 3427 36446 3483 36502
rect 3569 36446 3625 36502
rect 3711 36446 3767 36502
rect 3853 36446 3909 36502
rect 3995 36446 4051 36502
rect 4137 36446 4193 36502
rect 4279 36446 4335 36502
rect 4421 36446 4477 36502
rect 4563 36446 4619 36502
rect 4705 36446 4761 36502
rect 4847 36446 4903 36502
rect 4989 36446 5045 36502
rect 5131 36446 5187 36502
rect 5273 36446 5329 36502
rect 5415 36446 5471 36502
rect 5557 36446 5613 36502
rect 5699 36446 5755 36502
rect 5841 36446 5897 36502
rect 5983 36446 6039 36502
rect 6125 36446 6181 36502
rect 6267 36446 6323 36502
rect 6409 36446 6465 36502
rect 6551 36446 6607 36502
rect 6693 36446 6749 36502
rect 6835 36446 6891 36502
rect 6977 36446 7033 36502
rect 7119 36446 7175 36502
rect 7261 36446 7317 36502
rect 7403 36446 7459 36502
rect 7545 36446 7601 36502
rect 7687 36446 7743 36502
rect 7829 36446 7885 36502
rect 7971 36446 8027 36502
rect 8113 36446 8169 36502
rect 8255 36446 8311 36502
rect 8397 36446 8453 36502
rect 8539 36446 8595 36502
rect 8681 36446 8737 36502
rect 8823 36446 8879 36502
rect 8965 36446 9021 36502
rect 9107 36446 9163 36502
rect 9249 36446 9305 36502
rect 9391 36446 9447 36502
rect 9533 36446 9589 36502
rect 9675 36446 9731 36502
rect 9817 36446 9873 36502
rect 9959 36446 10015 36502
rect 10101 36446 10157 36502
rect 10243 36446 10299 36502
rect 10385 36446 10441 36502
rect 10527 36446 10583 36502
rect 10669 36446 10725 36502
rect 10811 36446 10867 36502
rect 10953 36446 11009 36502
rect 11095 36446 11151 36502
rect 11237 36446 11293 36502
rect 11379 36446 11435 36502
rect 11521 36446 11577 36502
rect 11663 36446 11719 36502
rect 11805 36446 11861 36502
rect 11947 36446 12003 36502
rect 12089 36446 12145 36502
rect 12231 36446 12287 36502
rect 12373 36446 12429 36502
rect 12515 36446 12571 36502
rect 12657 36446 12713 36502
rect 12799 36446 12855 36502
rect 12941 36446 12997 36502
rect 13083 36446 13139 36502
rect 13225 36446 13281 36502
rect 13367 36446 13423 36502
rect 13509 36446 13565 36502
rect 13651 36446 13707 36502
rect 13793 36446 13849 36502
rect 13935 36446 13991 36502
rect 14077 36446 14133 36502
rect 14219 36446 14275 36502
rect 14361 36446 14417 36502
rect 14503 36446 14559 36502
rect 14645 36446 14701 36502
rect 14787 36446 14843 36502
rect 161 36086 217 36142
rect 303 36086 359 36142
rect 445 36086 501 36142
rect 587 36086 643 36142
rect 729 36086 785 36142
rect 871 36086 927 36142
rect 1013 36086 1069 36142
rect 1155 36086 1211 36142
rect 1297 36086 1353 36142
rect 1439 36086 1495 36142
rect 1581 36086 1637 36142
rect 1723 36086 1779 36142
rect 1865 36086 1921 36142
rect 2007 36086 2063 36142
rect 2149 36086 2205 36142
rect 2291 36086 2347 36142
rect 2433 36086 2489 36142
rect 2575 36086 2631 36142
rect 2717 36086 2773 36142
rect 2859 36086 2915 36142
rect 3001 36086 3057 36142
rect 3143 36086 3199 36142
rect 3285 36086 3341 36142
rect 3427 36086 3483 36142
rect 3569 36086 3625 36142
rect 3711 36086 3767 36142
rect 3853 36086 3909 36142
rect 3995 36086 4051 36142
rect 4137 36086 4193 36142
rect 4279 36086 4335 36142
rect 4421 36086 4477 36142
rect 4563 36086 4619 36142
rect 4705 36086 4761 36142
rect 4847 36086 4903 36142
rect 4989 36086 5045 36142
rect 5131 36086 5187 36142
rect 5273 36086 5329 36142
rect 5415 36086 5471 36142
rect 5557 36086 5613 36142
rect 5699 36086 5755 36142
rect 5841 36086 5897 36142
rect 5983 36086 6039 36142
rect 6125 36086 6181 36142
rect 6267 36086 6323 36142
rect 6409 36086 6465 36142
rect 6551 36086 6607 36142
rect 6693 36086 6749 36142
rect 6835 36086 6891 36142
rect 6977 36086 7033 36142
rect 7119 36086 7175 36142
rect 7261 36086 7317 36142
rect 7403 36086 7459 36142
rect 7545 36086 7601 36142
rect 7687 36086 7743 36142
rect 7829 36086 7885 36142
rect 7971 36086 8027 36142
rect 8113 36086 8169 36142
rect 8255 36086 8311 36142
rect 8397 36086 8453 36142
rect 8539 36086 8595 36142
rect 8681 36086 8737 36142
rect 8823 36086 8879 36142
rect 8965 36086 9021 36142
rect 9107 36086 9163 36142
rect 9249 36086 9305 36142
rect 9391 36086 9447 36142
rect 9533 36086 9589 36142
rect 9675 36086 9731 36142
rect 9817 36086 9873 36142
rect 9959 36086 10015 36142
rect 10101 36086 10157 36142
rect 10243 36086 10299 36142
rect 10385 36086 10441 36142
rect 10527 36086 10583 36142
rect 10669 36086 10725 36142
rect 10811 36086 10867 36142
rect 10953 36086 11009 36142
rect 11095 36086 11151 36142
rect 11237 36086 11293 36142
rect 11379 36086 11435 36142
rect 11521 36086 11577 36142
rect 11663 36086 11719 36142
rect 11805 36086 11861 36142
rect 11947 36086 12003 36142
rect 12089 36086 12145 36142
rect 12231 36086 12287 36142
rect 12373 36086 12429 36142
rect 12515 36086 12571 36142
rect 12657 36086 12713 36142
rect 12799 36086 12855 36142
rect 12941 36086 12997 36142
rect 13083 36086 13139 36142
rect 13225 36086 13281 36142
rect 13367 36086 13423 36142
rect 13509 36086 13565 36142
rect 13651 36086 13707 36142
rect 13793 36086 13849 36142
rect 13935 36086 13991 36142
rect 14077 36086 14133 36142
rect 14219 36086 14275 36142
rect 14361 36086 14417 36142
rect 14503 36086 14559 36142
rect 14645 36086 14701 36142
rect 14787 36086 14843 36142
rect 161 35944 217 36000
rect 303 35944 359 36000
rect 445 35944 501 36000
rect 587 35944 643 36000
rect 729 35944 785 36000
rect 871 35944 927 36000
rect 1013 35944 1069 36000
rect 1155 35944 1211 36000
rect 1297 35944 1353 36000
rect 1439 35944 1495 36000
rect 1581 35944 1637 36000
rect 1723 35944 1779 36000
rect 1865 35944 1921 36000
rect 2007 35944 2063 36000
rect 2149 35944 2205 36000
rect 2291 35944 2347 36000
rect 2433 35944 2489 36000
rect 2575 35944 2631 36000
rect 2717 35944 2773 36000
rect 2859 35944 2915 36000
rect 3001 35944 3057 36000
rect 3143 35944 3199 36000
rect 3285 35944 3341 36000
rect 3427 35944 3483 36000
rect 3569 35944 3625 36000
rect 3711 35944 3767 36000
rect 3853 35944 3909 36000
rect 3995 35944 4051 36000
rect 4137 35944 4193 36000
rect 4279 35944 4335 36000
rect 4421 35944 4477 36000
rect 4563 35944 4619 36000
rect 4705 35944 4761 36000
rect 4847 35944 4903 36000
rect 4989 35944 5045 36000
rect 5131 35944 5187 36000
rect 5273 35944 5329 36000
rect 5415 35944 5471 36000
rect 5557 35944 5613 36000
rect 5699 35944 5755 36000
rect 5841 35944 5897 36000
rect 5983 35944 6039 36000
rect 6125 35944 6181 36000
rect 6267 35944 6323 36000
rect 6409 35944 6465 36000
rect 6551 35944 6607 36000
rect 6693 35944 6749 36000
rect 6835 35944 6891 36000
rect 6977 35944 7033 36000
rect 7119 35944 7175 36000
rect 7261 35944 7317 36000
rect 7403 35944 7459 36000
rect 7545 35944 7601 36000
rect 7687 35944 7743 36000
rect 7829 35944 7885 36000
rect 7971 35944 8027 36000
rect 8113 35944 8169 36000
rect 8255 35944 8311 36000
rect 8397 35944 8453 36000
rect 8539 35944 8595 36000
rect 8681 35944 8737 36000
rect 8823 35944 8879 36000
rect 8965 35944 9021 36000
rect 9107 35944 9163 36000
rect 9249 35944 9305 36000
rect 9391 35944 9447 36000
rect 9533 35944 9589 36000
rect 9675 35944 9731 36000
rect 9817 35944 9873 36000
rect 9959 35944 10015 36000
rect 10101 35944 10157 36000
rect 10243 35944 10299 36000
rect 10385 35944 10441 36000
rect 10527 35944 10583 36000
rect 10669 35944 10725 36000
rect 10811 35944 10867 36000
rect 10953 35944 11009 36000
rect 11095 35944 11151 36000
rect 11237 35944 11293 36000
rect 11379 35944 11435 36000
rect 11521 35944 11577 36000
rect 11663 35944 11719 36000
rect 11805 35944 11861 36000
rect 11947 35944 12003 36000
rect 12089 35944 12145 36000
rect 12231 35944 12287 36000
rect 12373 35944 12429 36000
rect 12515 35944 12571 36000
rect 12657 35944 12713 36000
rect 12799 35944 12855 36000
rect 12941 35944 12997 36000
rect 13083 35944 13139 36000
rect 13225 35944 13281 36000
rect 13367 35944 13423 36000
rect 13509 35944 13565 36000
rect 13651 35944 13707 36000
rect 13793 35944 13849 36000
rect 13935 35944 13991 36000
rect 14077 35944 14133 36000
rect 14219 35944 14275 36000
rect 14361 35944 14417 36000
rect 14503 35944 14559 36000
rect 14645 35944 14701 36000
rect 14787 35944 14843 36000
rect 161 35802 217 35858
rect 303 35802 359 35858
rect 445 35802 501 35858
rect 587 35802 643 35858
rect 729 35802 785 35858
rect 871 35802 927 35858
rect 1013 35802 1069 35858
rect 1155 35802 1211 35858
rect 1297 35802 1353 35858
rect 1439 35802 1495 35858
rect 1581 35802 1637 35858
rect 1723 35802 1779 35858
rect 1865 35802 1921 35858
rect 2007 35802 2063 35858
rect 2149 35802 2205 35858
rect 2291 35802 2347 35858
rect 2433 35802 2489 35858
rect 2575 35802 2631 35858
rect 2717 35802 2773 35858
rect 2859 35802 2915 35858
rect 3001 35802 3057 35858
rect 3143 35802 3199 35858
rect 3285 35802 3341 35858
rect 3427 35802 3483 35858
rect 3569 35802 3625 35858
rect 3711 35802 3767 35858
rect 3853 35802 3909 35858
rect 3995 35802 4051 35858
rect 4137 35802 4193 35858
rect 4279 35802 4335 35858
rect 4421 35802 4477 35858
rect 4563 35802 4619 35858
rect 4705 35802 4761 35858
rect 4847 35802 4903 35858
rect 4989 35802 5045 35858
rect 5131 35802 5187 35858
rect 5273 35802 5329 35858
rect 5415 35802 5471 35858
rect 5557 35802 5613 35858
rect 5699 35802 5755 35858
rect 5841 35802 5897 35858
rect 5983 35802 6039 35858
rect 6125 35802 6181 35858
rect 6267 35802 6323 35858
rect 6409 35802 6465 35858
rect 6551 35802 6607 35858
rect 6693 35802 6749 35858
rect 6835 35802 6891 35858
rect 6977 35802 7033 35858
rect 7119 35802 7175 35858
rect 7261 35802 7317 35858
rect 7403 35802 7459 35858
rect 7545 35802 7601 35858
rect 7687 35802 7743 35858
rect 7829 35802 7885 35858
rect 7971 35802 8027 35858
rect 8113 35802 8169 35858
rect 8255 35802 8311 35858
rect 8397 35802 8453 35858
rect 8539 35802 8595 35858
rect 8681 35802 8737 35858
rect 8823 35802 8879 35858
rect 8965 35802 9021 35858
rect 9107 35802 9163 35858
rect 9249 35802 9305 35858
rect 9391 35802 9447 35858
rect 9533 35802 9589 35858
rect 9675 35802 9731 35858
rect 9817 35802 9873 35858
rect 9959 35802 10015 35858
rect 10101 35802 10157 35858
rect 10243 35802 10299 35858
rect 10385 35802 10441 35858
rect 10527 35802 10583 35858
rect 10669 35802 10725 35858
rect 10811 35802 10867 35858
rect 10953 35802 11009 35858
rect 11095 35802 11151 35858
rect 11237 35802 11293 35858
rect 11379 35802 11435 35858
rect 11521 35802 11577 35858
rect 11663 35802 11719 35858
rect 11805 35802 11861 35858
rect 11947 35802 12003 35858
rect 12089 35802 12145 35858
rect 12231 35802 12287 35858
rect 12373 35802 12429 35858
rect 12515 35802 12571 35858
rect 12657 35802 12713 35858
rect 12799 35802 12855 35858
rect 12941 35802 12997 35858
rect 13083 35802 13139 35858
rect 13225 35802 13281 35858
rect 13367 35802 13423 35858
rect 13509 35802 13565 35858
rect 13651 35802 13707 35858
rect 13793 35802 13849 35858
rect 13935 35802 13991 35858
rect 14077 35802 14133 35858
rect 14219 35802 14275 35858
rect 14361 35802 14417 35858
rect 14503 35802 14559 35858
rect 14645 35802 14701 35858
rect 14787 35802 14843 35858
rect 161 35660 217 35716
rect 303 35660 359 35716
rect 445 35660 501 35716
rect 587 35660 643 35716
rect 729 35660 785 35716
rect 871 35660 927 35716
rect 1013 35660 1069 35716
rect 1155 35660 1211 35716
rect 1297 35660 1353 35716
rect 1439 35660 1495 35716
rect 1581 35660 1637 35716
rect 1723 35660 1779 35716
rect 1865 35660 1921 35716
rect 2007 35660 2063 35716
rect 2149 35660 2205 35716
rect 2291 35660 2347 35716
rect 2433 35660 2489 35716
rect 2575 35660 2631 35716
rect 2717 35660 2773 35716
rect 2859 35660 2915 35716
rect 3001 35660 3057 35716
rect 3143 35660 3199 35716
rect 3285 35660 3341 35716
rect 3427 35660 3483 35716
rect 3569 35660 3625 35716
rect 3711 35660 3767 35716
rect 3853 35660 3909 35716
rect 3995 35660 4051 35716
rect 4137 35660 4193 35716
rect 4279 35660 4335 35716
rect 4421 35660 4477 35716
rect 4563 35660 4619 35716
rect 4705 35660 4761 35716
rect 4847 35660 4903 35716
rect 4989 35660 5045 35716
rect 5131 35660 5187 35716
rect 5273 35660 5329 35716
rect 5415 35660 5471 35716
rect 5557 35660 5613 35716
rect 5699 35660 5755 35716
rect 5841 35660 5897 35716
rect 5983 35660 6039 35716
rect 6125 35660 6181 35716
rect 6267 35660 6323 35716
rect 6409 35660 6465 35716
rect 6551 35660 6607 35716
rect 6693 35660 6749 35716
rect 6835 35660 6891 35716
rect 6977 35660 7033 35716
rect 7119 35660 7175 35716
rect 7261 35660 7317 35716
rect 7403 35660 7459 35716
rect 7545 35660 7601 35716
rect 7687 35660 7743 35716
rect 7829 35660 7885 35716
rect 7971 35660 8027 35716
rect 8113 35660 8169 35716
rect 8255 35660 8311 35716
rect 8397 35660 8453 35716
rect 8539 35660 8595 35716
rect 8681 35660 8737 35716
rect 8823 35660 8879 35716
rect 8965 35660 9021 35716
rect 9107 35660 9163 35716
rect 9249 35660 9305 35716
rect 9391 35660 9447 35716
rect 9533 35660 9589 35716
rect 9675 35660 9731 35716
rect 9817 35660 9873 35716
rect 9959 35660 10015 35716
rect 10101 35660 10157 35716
rect 10243 35660 10299 35716
rect 10385 35660 10441 35716
rect 10527 35660 10583 35716
rect 10669 35660 10725 35716
rect 10811 35660 10867 35716
rect 10953 35660 11009 35716
rect 11095 35660 11151 35716
rect 11237 35660 11293 35716
rect 11379 35660 11435 35716
rect 11521 35660 11577 35716
rect 11663 35660 11719 35716
rect 11805 35660 11861 35716
rect 11947 35660 12003 35716
rect 12089 35660 12145 35716
rect 12231 35660 12287 35716
rect 12373 35660 12429 35716
rect 12515 35660 12571 35716
rect 12657 35660 12713 35716
rect 12799 35660 12855 35716
rect 12941 35660 12997 35716
rect 13083 35660 13139 35716
rect 13225 35660 13281 35716
rect 13367 35660 13423 35716
rect 13509 35660 13565 35716
rect 13651 35660 13707 35716
rect 13793 35660 13849 35716
rect 13935 35660 13991 35716
rect 14077 35660 14133 35716
rect 14219 35660 14275 35716
rect 14361 35660 14417 35716
rect 14503 35660 14559 35716
rect 14645 35660 14701 35716
rect 14787 35660 14843 35716
rect 161 35518 217 35574
rect 303 35518 359 35574
rect 445 35518 501 35574
rect 587 35518 643 35574
rect 729 35518 785 35574
rect 871 35518 927 35574
rect 1013 35518 1069 35574
rect 1155 35518 1211 35574
rect 1297 35518 1353 35574
rect 1439 35518 1495 35574
rect 1581 35518 1637 35574
rect 1723 35518 1779 35574
rect 1865 35518 1921 35574
rect 2007 35518 2063 35574
rect 2149 35518 2205 35574
rect 2291 35518 2347 35574
rect 2433 35518 2489 35574
rect 2575 35518 2631 35574
rect 2717 35518 2773 35574
rect 2859 35518 2915 35574
rect 3001 35518 3057 35574
rect 3143 35518 3199 35574
rect 3285 35518 3341 35574
rect 3427 35518 3483 35574
rect 3569 35518 3625 35574
rect 3711 35518 3767 35574
rect 3853 35518 3909 35574
rect 3995 35518 4051 35574
rect 4137 35518 4193 35574
rect 4279 35518 4335 35574
rect 4421 35518 4477 35574
rect 4563 35518 4619 35574
rect 4705 35518 4761 35574
rect 4847 35518 4903 35574
rect 4989 35518 5045 35574
rect 5131 35518 5187 35574
rect 5273 35518 5329 35574
rect 5415 35518 5471 35574
rect 5557 35518 5613 35574
rect 5699 35518 5755 35574
rect 5841 35518 5897 35574
rect 5983 35518 6039 35574
rect 6125 35518 6181 35574
rect 6267 35518 6323 35574
rect 6409 35518 6465 35574
rect 6551 35518 6607 35574
rect 6693 35518 6749 35574
rect 6835 35518 6891 35574
rect 6977 35518 7033 35574
rect 7119 35518 7175 35574
rect 7261 35518 7317 35574
rect 7403 35518 7459 35574
rect 7545 35518 7601 35574
rect 7687 35518 7743 35574
rect 7829 35518 7885 35574
rect 7971 35518 8027 35574
rect 8113 35518 8169 35574
rect 8255 35518 8311 35574
rect 8397 35518 8453 35574
rect 8539 35518 8595 35574
rect 8681 35518 8737 35574
rect 8823 35518 8879 35574
rect 8965 35518 9021 35574
rect 9107 35518 9163 35574
rect 9249 35518 9305 35574
rect 9391 35518 9447 35574
rect 9533 35518 9589 35574
rect 9675 35518 9731 35574
rect 9817 35518 9873 35574
rect 9959 35518 10015 35574
rect 10101 35518 10157 35574
rect 10243 35518 10299 35574
rect 10385 35518 10441 35574
rect 10527 35518 10583 35574
rect 10669 35518 10725 35574
rect 10811 35518 10867 35574
rect 10953 35518 11009 35574
rect 11095 35518 11151 35574
rect 11237 35518 11293 35574
rect 11379 35518 11435 35574
rect 11521 35518 11577 35574
rect 11663 35518 11719 35574
rect 11805 35518 11861 35574
rect 11947 35518 12003 35574
rect 12089 35518 12145 35574
rect 12231 35518 12287 35574
rect 12373 35518 12429 35574
rect 12515 35518 12571 35574
rect 12657 35518 12713 35574
rect 12799 35518 12855 35574
rect 12941 35518 12997 35574
rect 13083 35518 13139 35574
rect 13225 35518 13281 35574
rect 13367 35518 13423 35574
rect 13509 35518 13565 35574
rect 13651 35518 13707 35574
rect 13793 35518 13849 35574
rect 13935 35518 13991 35574
rect 14077 35518 14133 35574
rect 14219 35518 14275 35574
rect 14361 35518 14417 35574
rect 14503 35518 14559 35574
rect 14645 35518 14701 35574
rect 14787 35518 14843 35574
rect 161 35376 217 35432
rect 303 35376 359 35432
rect 445 35376 501 35432
rect 587 35376 643 35432
rect 729 35376 785 35432
rect 871 35376 927 35432
rect 1013 35376 1069 35432
rect 1155 35376 1211 35432
rect 1297 35376 1353 35432
rect 1439 35376 1495 35432
rect 1581 35376 1637 35432
rect 1723 35376 1779 35432
rect 1865 35376 1921 35432
rect 2007 35376 2063 35432
rect 2149 35376 2205 35432
rect 2291 35376 2347 35432
rect 2433 35376 2489 35432
rect 2575 35376 2631 35432
rect 2717 35376 2773 35432
rect 2859 35376 2915 35432
rect 3001 35376 3057 35432
rect 3143 35376 3199 35432
rect 3285 35376 3341 35432
rect 3427 35376 3483 35432
rect 3569 35376 3625 35432
rect 3711 35376 3767 35432
rect 3853 35376 3909 35432
rect 3995 35376 4051 35432
rect 4137 35376 4193 35432
rect 4279 35376 4335 35432
rect 4421 35376 4477 35432
rect 4563 35376 4619 35432
rect 4705 35376 4761 35432
rect 4847 35376 4903 35432
rect 4989 35376 5045 35432
rect 5131 35376 5187 35432
rect 5273 35376 5329 35432
rect 5415 35376 5471 35432
rect 5557 35376 5613 35432
rect 5699 35376 5755 35432
rect 5841 35376 5897 35432
rect 5983 35376 6039 35432
rect 6125 35376 6181 35432
rect 6267 35376 6323 35432
rect 6409 35376 6465 35432
rect 6551 35376 6607 35432
rect 6693 35376 6749 35432
rect 6835 35376 6891 35432
rect 6977 35376 7033 35432
rect 7119 35376 7175 35432
rect 7261 35376 7317 35432
rect 7403 35376 7459 35432
rect 7545 35376 7601 35432
rect 7687 35376 7743 35432
rect 7829 35376 7885 35432
rect 7971 35376 8027 35432
rect 8113 35376 8169 35432
rect 8255 35376 8311 35432
rect 8397 35376 8453 35432
rect 8539 35376 8595 35432
rect 8681 35376 8737 35432
rect 8823 35376 8879 35432
rect 8965 35376 9021 35432
rect 9107 35376 9163 35432
rect 9249 35376 9305 35432
rect 9391 35376 9447 35432
rect 9533 35376 9589 35432
rect 9675 35376 9731 35432
rect 9817 35376 9873 35432
rect 9959 35376 10015 35432
rect 10101 35376 10157 35432
rect 10243 35376 10299 35432
rect 10385 35376 10441 35432
rect 10527 35376 10583 35432
rect 10669 35376 10725 35432
rect 10811 35376 10867 35432
rect 10953 35376 11009 35432
rect 11095 35376 11151 35432
rect 11237 35376 11293 35432
rect 11379 35376 11435 35432
rect 11521 35376 11577 35432
rect 11663 35376 11719 35432
rect 11805 35376 11861 35432
rect 11947 35376 12003 35432
rect 12089 35376 12145 35432
rect 12231 35376 12287 35432
rect 12373 35376 12429 35432
rect 12515 35376 12571 35432
rect 12657 35376 12713 35432
rect 12799 35376 12855 35432
rect 12941 35376 12997 35432
rect 13083 35376 13139 35432
rect 13225 35376 13281 35432
rect 13367 35376 13423 35432
rect 13509 35376 13565 35432
rect 13651 35376 13707 35432
rect 13793 35376 13849 35432
rect 13935 35376 13991 35432
rect 14077 35376 14133 35432
rect 14219 35376 14275 35432
rect 14361 35376 14417 35432
rect 14503 35376 14559 35432
rect 14645 35376 14701 35432
rect 14787 35376 14843 35432
rect 161 35234 217 35290
rect 303 35234 359 35290
rect 445 35234 501 35290
rect 587 35234 643 35290
rect 729 35234 785 35290
rect 871 35234 927 35290
rect 1013 35234 1069 35290
rect 1155 35234 1211 35290
rect 1297 35234 1353 35290
rect 1439 35234 1495 35290
rect 1581 35234 1637 35290
rect 1723 35234 1779 35290
rect 1865 35234 1921 35290
rect 2007 35234 2063 35290
rect 2149 35234 2205 35290
rect 2291 35234 2347 35290
rect 2433 35234 2489 35290
rect 2575 35234 2631 35290
rect 2717 35234 2773 35290
rect 2859 35234 2915 35290
rect 3001 35234 3057 35290
rect 3143 35234 3199 35290
rect 3285 35234 3341 35290
rect 3427 35234 3483 35290
rect 3569 35234 3625 35290
rect 3711 35234 3767 35290
rect 3853 35234 3909 35290
rect 3995 35234 4051 35290
rect 4137 35234 4193 35290
rect 4279 35234 4335 35290
rect 4421 35234 4477 35290
rect 4563 35234 4619 35290
rect 4705 35234 4761 35290
rect 4847 35234 4903 35290
rect 4989 35234 5045 35290
rect 5131 35234 5187 35290
rect 5273 35234 5329 35290
rect 5415 35234 5471 35290
rect 5557 35234 5613 35290
rect 5699 35234 5755 35290
rect 5841 35234 5897 35290
rect 5983 35234 6039 35290
rect 6125 35234 6181 35290
rect 6267 35234 6323 35290
rect 6409 35234 6465 35290
rect 6551 35234 6607 35290
rect 6693 35234 6749 35290
rect 6835 35234 6891 35290
rect 6977 35234 7033 35290
rect 7119 35234 7175 35290
rect 7261 35234 7317 35290
rect 7403 35234 7459 35290
rect 7545 35234 7601 35290
rect 7687 35234 7743 35290
rect 7829 35234 7885 35290
rect 7971 35234 8027 35290
rect 8113 35234 8169 35290
rect 8255 35234 8311 35290
rect 8397 35234 8453 35290
rect 8539 35234 8595 35290
rect 8681 35234 8737 35290
rect 8823 35234 8879 35290
rect 8965 35234 9021 35290
rect 9107 35234 9163 35290
rect 9249 35234 9305 35290
rect 9391 35234 9447 35290
rect 9533 35234 9589 35290
rect 9675 35234 9731 35290
rect 9817 35234 9873 35290
rect 9959 35234 10015 35290
rect 10101 35234 10157 35290
rect 10243 35234 10299 35290
rect 10385 35234 10441 35290
rect 10527 35234 10583 35290
rect 10669 35234 10725 35290
rect 10811 35234 10867 35290
rect 10953 35234 11009 35290
rect 11095 35234 11151 35290
rect 11237 35234 11293 35290
rect 11379 35234 11435 35290
rect 11521 35234 11577 35290
rect 11663 35234 11719 35290
rect 11805 35234 11861 35290
rect 11947 35234 12003 35290
rect 12089 35234 12145 35290
rect 12231 35234 12287 35290
rect 12373 35234 12429 35290
rect 12515 35234 12571 35290
rect 12657 35234 12713 35290
rect 12799 35234 12855 35290
rect 12941 35234 12997 35290
rect 13083 35234 13139 35290
rect 13225 35234 13281 35290
rect 13367 35234 13423 35290
rect 13509 35234 13565 35290
rect 13651 35234 13707 35290
rect 13793 35234 13849 35290
rect 13935 35234 13991 35290
rect 14077 35234 14133 35290
rect 14219 35234 14275 35290
rect 14361 35234 14417 35290
rect 14503 35234 14559 35290
rect 14645 35234 14701 35290
rect 14787 35234 14843 35290
rect 161 35092 217 35148
rect 303 35092 359 35148
rect 445 35092 501 35148
rect 587 35092 643 35148
rect 729 35092 785 35148
rect 871 35092 927 35148
rect 1013 35092 1069 35148
rect 1155 35092 1211 35148
rect 1297 35092 1353 35148
rect 1439 35092 1495 35148
rect 1581 35092 1637 35148
rect 1723 35092 1779 35148
rect 1865 35092 1921 35148
rect 2007 35092 2063 35148
rect 2149 35092 2205 35148
rect 2291 35092 2347 35148
rect 2433 35092 2489 35148
rect 2575 35092 2631 35148
rect 2717 35092 2773 35148
rect 2859 35092 2915 35148
rect 3001 35092 3057 35148
rect 3143 35092 3199 35148
rect 3285 35092 3341 35148
rect 3427 35092 3483 35148
rect 3569 35092 3625 35148
rect 3711 35092 3767 35148
rect 3853 35092 3909 35148
rect 3995 35092 4051 35148
rect 4137 35092 4193 35148
rect 4279 35092 4335 35148
rect 4421 35092 4477 35148
rect 4563 35092 4619 35148
rect 4705 35092 4761 35148
rect 4847 35092 4903 35148
rect 4989 35092 5045 35148
rect 5131 35092 5187 35148
rect 5273 35092 5329 35148
rect 5415 35092 5471 35148
rect 5557 35092 5613 35148
rect 5699 35092 5755 35148
rect 5841 35092 5897 35148
rect 5983 35092 6039 35148
rect 6125 35092 6181 35148
rect 6267 35092 6323 35148
rect 6409 35092 6465 35148
rect 6551 35092 6607 35148
rect 6693 35092 6749 35148
rect 6835 35092 6891 35148
rect 6977 35092 7033 35148
rect 7119 35092 7175 35148
rect 7261 35092 7317 35148
rect 7403 35092 7459 35148
rect 7545 35092 7601 35148
rect 7687 35092 7743 35148
rect 7829 35092 7885 35148
rect 7971 35092 8027 35148
rect 8113 35092 8169 35148
rect 8255 35092 8311 35148
rect 8397 35092 8453 35148
rect 8539 35092 8595 35148
rect 8681 35092 8737 35148
rect 8823 35092 8879 35148
rect 8965 35092 9021 35148
rect 9107 35092 9163 35148
rect 9249 35092 9305 35148
rect 9391 35092 9447 35148
rect 9533 35092 9589 35148
rect 9675 35092 9731 35148
rect 9817 35092 9873 35148
rect 9959 35092 10015 35148
rect 10101 35092 10157 35148
rect 10243 35092 10299 35148
rect 10385 35092 10441 35148
rect 10527 35092 10583 35148
rect 10669 35092 10725 35148
rect 10811 35092 10867 35148
rect 10953 35092 11009 35148
rect 11095 35092 11151 35148
rect 11237 35092 11293 35148
rect 11379 35092 11435 35148
rect 11521 35092 11577 35148
rect 11663 35092 11719 35148
rect 11805 35092 11861 35148
rect 11947 35092 12003 35148
rect 12089 35092 12145 35148
rect 12231 35092 12287 35148
rect 12373 35092 12429 35148
rect 12515 35092 12571 35148
rect 12657 35092 12713 35148
rect 12799 35092 12855 35148
rect 12941 35092 12997 35148
rect 13083 35092 13139 35148
rect 13225 35092 13281 35148
rect 13367 35092 13423 35148
rect 13509 35092 13565 35148
rect 13651 35092 13707 35148
rect 13793 35092 13849 35148
rect 13935 35092 13991 35148
rect 14077 35092 14133 35148
rect 14219 35092 14275 35148
rect 14361 35092 14417 35148
rect 14503 35092 14559 35148
rect 14645 35092 14701 35148
rect 14787 35092 14843 35148
rect 161 34950 217 35006
rect 303 34950 359 35006
rect 445 34950 501 35006
rect 587 34950 643 35006
rect 729 34950 785 35006
rect 871 34950 927 35006
rect 1013 34950 1069 35006
rect 1155 34950 1211 35006
rect 1297 34950 1353 35006
rect 1439 34950 1495 35006
rect 1581 34950 1637 35006
rect 1723 34950 1779 35006
rect 1865 34950 1921 35006
rect 2007 34950 2063 35006
rect 2149 34950 2205 35006
rect 2291 34950 2347 35006
rect 2433 34950 2489 35006
rect 2575 34950 2631 35006
rect 2717 34950 2773 35006
rect 2859 34950 2915 35006
rect 3001 34950 3057 35006
rect 3143 34950 3199 35006
rect 3285 34950 3341 35006
rect 3427 34950 3483 35006
rect 3569 34950 3625 35006
rect 3711 34950 3767 35006
rect 3853 34950 3909 35006
rect 3995 34950 4051 35006
rect 4137 34950 4193 35006
rect 4279 34950 4335 35006
rect 4421 34950 4477 35006
rect 4563 34950 4619 35006
rect 4705 34950 4761 35006
rect 4847 34950 4903 35006
rect 4989 34950 5045 35006
rect 5131 34950 5187 35006
rect 5273 34950 5329 35006
rect 5415 34950 5471 35006
rect 5557 34950 5613 35006
rect 5699 34950 5755 35006
rect 5841 34950 5897 35006
rect 5983 34950 6039 35006
rect 6125 34950 6181 35006
rect 6267 34950 6323 35006
rect 6409 34950 6465 35006
rect 6551 34950 6607 35006
rect 6693 34950 6749 35006
rect 6835 34950 6891 35006
rect 6977 34950 7033 35006
rect 7119 34950 7175 35006
rect 7261 34950 7317 35006
rect 7403 34950 7459 35006
rect 7545 34950 7601 35006
rect 7687 34950 7743 35006
rect 7829 34950 7885 35006
rect 7971 34950 8027 35006
rect 8113 34950 8169 35006
rect 8255 34950 8311 35006
rect 8397 34950 8453 35006
rect 8539 34950 8595 35006
rect 8681 34950 8737 35006
rect 8823 34950 8879 35006
rect 8965 34950 9021 35006
rect 9107 34950 9163 35006
rect 9249 34950 9305 35006
rect 9391 34950 9447 35006
rect 9533 34950 9589 35006
rect 9675 34950 9731 35006
rect 9817 34950 9873 35006
rect 9959 34950 10015 35006
rect 10101 34950 10157 35006
rect 10243 34950 10299 35006
rect 10385 34950 10441 35006
rect 10527 34950 10583 35006
rect 10669 34950 10725 35006
rect 10811 34950 10867 35006
rect 10953 34950 11009 35006
rect 11095 34950 11151 35006
rect 11237 34950 11293 35006
rect 11379 34950 11435 35006
rect 11521 34950 11577 35006
rect 11663 34950 11719 35006
rect 11805 34950 11861 35006
rect 11947 34950 12003 35006
rect 12089 34950 12145 35006
rect 12231 34950 12287 35006
rect 12373 34950 12429 35006
rect 12515 34950 12571 35006
rect 12657 34950 12713 35006
rect 12799 34950 12855 35006
rect 12941 34950 12997 35006
rect 13083 34950 13139 35006
rect 13225 34950 13281 35006
rect 13367 34950 13423 35006
rect 13509 34950 13565 35006
rect 13651 34950 13707 35006
rect 13793 34950 13849 35006
rect 13935 34950 13991 35006
rect 14077 34950 14133 35006
rect 14219 34950 14275 35006
rect 14361 34950 14417 35006
rect 14503 34950 14559 35006
rect 14645 34950 14701 35006
rect 14787 34950 14843 35006
rect 161 34808 217 34864
rect 303 34808 359 34864
rect 445 34808 501 34864
rect 587 34808 643 34864
rect 729 34808 785 34864
rect 871 34808 927 34864
rect 1013 34808 1069 34864
rect 1155 34808 1211 34864
rect 1297 34808 1353 34864
rect 1439 34808 1495 34864
rect 1581 34808 1637 34864
rect 1723 34808 1779 34864
rect 1865 34808 1921 34864
rect 2007 34808 2063 34864
rect 2149 34808 2205 34864
rect 2291 34808 2347 34864
rect 2433 34808 2489 34864
rect 2575 34808 2631 34864
rect 2717 34808 2773 34864
rect 2859 34808 2915 34864
rect 3001 34808 3057 34864
rect 3143 34808 3199 34864
rect 3285 34808 3341 34864
rect 3427 34808 3483 34864
rect 3569 34808 3625 34864
rect 3711 34808 3767 34864
rect 3853 34808 3909 34864
rect 3995 34808 4051 34864
rect 4137 34808 4193 34864
rect 4279 34808 4335 34864
rect 4421 34808 4477 34864
rect 4563 34808 4619 34864
rect 4705 34808 4761 34864
rect 4847 34808 4903 34864
rect 4989 34808 5045 34864
rect 5131 34808 5187 34864
rect 5273 34808 5329 34864
rect 5415 34808 5471 34864
rect 5557 34808 5613 34864
rect 5699 34808 5755 34864
rect 5841 34808 5897 34864
rect 5983 34808 6039 34864
rect 6125 34808 6181 34864
rect 6267 34808 6323 34864
rect 6409 34808 6465 34864
rect 6551 34808 6607 34864
rect 6693 34808 6749 34864
rect 6835 34808 6891 34864
rect 6977 34808 7033 34864
rect 7119 34808 7175 34864
rect 7261 34808 7317 34864
rect 7403 34808 7459 34864
rect 7545 34808 7601 34864
rect 7687 34808 7743 34864
rect 7829 34808 7885 34864
rect 7971 34808 8027 34864
rect 8113 34808 8169 34864
rect 8255 34808 8311 34864
rect 8397 34808 8453 34864
rect 8539 34808 8595 34864
rect 8681 34808 8737 34864
rect 8823 34808 8879 34864
rect 8965 34808 9021 34864
rect 9107 34808 9163 34864
rect 9249 34808 9305 34864
rect 9391 34808 9447 34864
rect 9533 34808 9589 34864
rect 9675 34808 9731 34864
rect 9817 34808 9873 34864
rect 9959 34808 10015 34864
rect 10101 34808 10157 34864
rect 10243 34808 10299 34864
rect 10385 34808 10441 34864
rect 10527 34808 10583 34864
rect 10669 34808 10725 34864
rect 10811 34808 10867 34864
rect 10953 34808 11009 34864
rect 11095 34808 11151 34864
rect 11237 34808 11293 34864
rect 11379 34808 11435 34864
rect 11521 34808 11577 34864
rect 11663 34808 11719 34864
rect 11805 34808 11861 34864
rect 11947 34808 12003 34864
rect 12089 34808 12145 34864
rect 12231 34808 12287 34864
rect 12373 34808 12429 34864
rect 12515 34808 12571 34864
rect 12657 34808 12713 34864
rect 12799 34808 12855 34864
rect 12941 34808 12997 34864
rect 13083 34808 13139 34864
rect 13225 34808 13281 34864
rect 13367 34808 13423 34864
rect 13509 34808 13565 34864
rect 13651 34808 13707 34864
rect 13793 34808 13849 34864
rect 13935 34808 13991 34864
rect 14077 34808 14133 34864
rect 14219 34808 14275 34864
rect 14361 34808 14417 34864
rect 14503 34808 14559 34864
rect 14645 34808 14701 34864
rect 14787 34808 14843 34864
rect 161 34666 217 34722
rect 303 34666 359 34722
rect 445 34666 501 34722
rect 587 34666 643 34722
rect 729 34666 785 34722
rect 871 34666 927 34722
rect 1013 34666 1069 34722
rect 1155 34666 1211 34722
rect 1297 34666 1353 34722
rect 1439 34666 1495 34722
rect 1581 34666 1637 34722
rect 1723 34666 1779 34722
rect 1865 34666 1921 34722
rect 2007 34666 2063 34722
rect 2149 34666 2205 34722
rect 2291 34666 2347 34722
rect 2433 34666 2489 34722
rect 2575 34666 2631 34722
rect 2717 34666 2773 34722
rect 2859 34666 2915 34722
rect 3001 34666 3057 34722
rect 3143 34666 3199 34722
rect 3285 34666 3341 34722
rect 3427 34666 3483 34722
rect 3569 34666 3625 34722
rect 3711 34666 3767 34722
rect 3853 34666 3909 34722
rect 3995 34666 4051 34722
rect 4137 34666 4193 34722
rect 4279 34666 4335 34722
rect 4421 34666 4477 34722
rect 4563 34666 4619 34722
rect 4705 34666 4761 34722
rect 4847 34666 4903 34722
rect 4989 34666 5045 34722
rect 5131 34666 5187 34722
rect 5273 34666 5329 34722
rect 5415 34666 5471 34722
rect 5557 34666 5613 34722
rect 5699 34666 5755 34722
rect 5841 34666 5897 34722
rect 5983 34666 6039 34722
rect 6125 34666 6181 34722
rect 6267 34666 6323 34722
rect 6409 34666 6465 34722
rect 6551 34666 6607 34722
rect 6693 34666 6749 34722
rect 6835 34666 6891 34722
rect 6977 34666 7033 34722
rect 7119 34666 7175 34722
rect 7261 34666 7317 34722
rect 7403 34666 7459 34722
rect 7545 34666 7601 34722
rect 7687 34666 7743 34722
rect 7829 34666 7885 34722
rect 7971 34666 8027 34722
rect 8113 34666 8169 34722
rect 8255 34666 8311 34722
rect 8397 34666 8453 34722
rect 8539 34666 8595 34722
rect 8681 34666 8737 34722
rect 8823 34666 8879 34722
rect 8965 34666 9021 34722
rect 9107 34666 9163 34722
rect 9249 34666 9305 34722
rect 9391 34666 9447 34722
rect 9533 34666 9589 34722
rect 9675 34666 9731 34722
rect 9817 34666 9873 34722
rect 9959 34666 10015 34722
rect 10101 34666 10157 34722
rect 10243 34666 10299 34722
rect 10385 34666 10441 34722
rect 10527 34666 10583 34722
rect 10669 34666 10725 34722
rect 10811 34666 10867 34722
rect 10953 34666 11009 34722
rect 11095 34666 11151 34722
rect 11237 34666 11293 34722
rect 11379 34666 11435 34722
rect 11521 34666 11577 34722
rect 11663 34666 11719 34722
rect 11805 34666 11861 34722
rect 11947 34666 12003 34722
rect 12089 34666 12145 34722
rect 12231 34666 12287 34722
rect 12373 34666 12429 34722
rect 12515 34666 12571 34722
rect 12657 34666 12713 34722
rect 12799 34666 12855 34722
rect 12941 34666 12997 34722
rect 13083 34666 13139 34722
rect 13225 34666 13281 34722
rect 13367 34666 13423 34722
rect 13509 34666 13565 34722
rect 13651 34666 13707 34722
rect 13793 34666 13849 34722
rect 13935 34666 13991 34722
rect 14077 34666 14133 34722
rect 14219 34666 14275 34722
rect 14361 34666 14417 34722
rect 14503 34666 14559 34722
rect 14645 34666 14701 34722
rect 14787 34666 14843 34722
rect 161 34524 217 34580
rect 303 34524 359 34580
rect 445 34524 501 34580
rect 587 34524 643 34580
rect 729 34524 785 34580
rect 871 34524 927 34580
rect 1013 34524 1069 34580
rect 1155 34524 1211 34580
rect 1297 34524 1353 34580
rect 1439 34524 1495 34580
rect 1581 34524 1637 34580
rect 1723 34524 1779 34580
rect 1865 34524 1921 34580
rect 2007 34524 2063 34580
rect 2149 34524 2205 34580
rect 2291 34524 2347 34580
rect 2433 34524 2489 34580
rect 2575 34524 2631 34580
rect 2717 34524 2773 34580
rect 2859 34524 2915 34580
rect 3001 34524 3057 34580
rect 3143 34524 3199 34580
rect 3285 34524 3341 34580
rect 3427 34524 3483 34580
rect 3569 34524 3625 34580
rect 3711 34524 3767 34580
rect 3853 34524 3909 34580
rect 3995 34524 4051 34580
rect 4137 34524 4193 34580
rect 4279 34524 4335 34580
rect 4421 34524 4477 34580
rect 4563 34524 4619 34580
rect 4705 34524 4761 34580
rect 4847 34524 4903 34580
rect 4989 34524 5045 34580
rect 5131 34524 5187 34580
rect 5273 34524 5329 34580
rect 5415 34524 5471 34580
rect 5557 34524 5613 34580
rect 5699 34524 5755 34580
rect 5841 34524 5897 34580
rect 5983 34524 6039 34580
rect 6125 34524 6181 34580
rect 6267 34524 6323 34580
rect 6409 34524 6465 34580
rect 6551 34524 6607 34580
rect 6693 34524 6749 34580
rect 6835 34524 6891 34580
rect 6977 34524 7033 34580
rect 7119 34524 7175 34580
rect 7261 34524 7317 34580
rect 7403 34524 7459 34580
rect 7545 34524 7601 34580
rect 7687 34524 7743 34580
rect 7829 34524 7885 34580
rect 7971 34524 8027 34580
rect 8113 34524 8169 34580
rect 8255 34524 8311 34580
rect 8397 34524 8453 34580
rect 8539 34524 8595 34580
rect 8681 34524 8737 34580
rect 8823 34524 8879 34580
rect 8965 34524 9021 34580
rect 9107 34524 9163 34580
rect 9249 34524 9305 34580
rect 9391 34524 9447 34580
rect 9533 34524 9589 34580
rect 9675 34524 9731 34580
rect 9817 34524 9873 34580
rect 9959 34524 10015 34580
rect 10101 34524 10157 34580
rect 10243 34524 10299 34580
rect 10385 34524 10441 34580
rect 10527 34524 10583 34580
rect 10669 34524 10725 34580
rect 10811 34524 10867 34580
rect 10953 34524 11009 34580
rect 11095 34524 11151 34580
rect 11237 34524 11293 34580
rect 11379 34524 11435 34580
rect 11521 34524 11577 34580
rect 11663 34524 11719 34580
rect 11805 34524 11861 34580
rect 11947 34524 12003 34580
rect 12089 34524 12145 34580
rect 12231 34524 12287 34580
rect 12373 34524 12429 34580
rect 12515 34524 12571 34580
rect 12657 34524 12713 34580
rect 12799 34524 12855 34580
rect 12941 34524 12997 34580
rect 13083 34524 13139 34580
rect 13225 34524 13281 34580
rect 13367 34524 13423 34580
rect 13509 34524 13565 34580
rect 13651 34524 13707 34580
rect 13793 34524 13849 34580
rect 13935 34524 13991 34580
rect 14077 34524 14133 34580
rect 14219 34524 14275 34580
rect 14361 34524 14417 34580
rect 14503 34524 14559 34580
rect 14645 34524 14701 34580
rect 14787 34524 14843 34580
rect 161 34382 217 34438
rect 303 34382 359 34438
rect 445 34382 501 34438
rect 587 34382 643 34438
rect 729 34382 785 34438
rect 871 34382 927 34438
rect 1013 34382 1069 34438
rect 1155 34382 1211 34438
rect 1297 34382 1353 34438
rect 1439 34382 1495 34438
rect 1581 34382 1637 34438
rect 1723 34382 1779 34438
rect 1865 34382 1921 34438
rect 2007 34382 2063 34438
rect 2149 34382 2205 34438
rect 2291 34382 2347 34438
rect 2433 34382 2489 34438
rect 2575 34382 2631 34438
rect 2717 34382 2773 34438
rect 2859 34382 2915 34438
rect 3001 34382 3057 34438
rect 3143 34382 3199 34438
rect 3285 34382 3341 34438
rect 3427 34382 3483 34438
rect 3569 34382 3625 34438
rect 3711 34382 3767 34438
rect 3853 34382 3909 34438
rect 3995 34382 4051 34438
rect 4137 34382 4193 34438
rect 4279 34382 4335 34438
rect 4421 34382 4477 34438
rect 4563 34382 4619 34438
rect 4705 34382 4761 34438
rect 4847 34382 4903 34438
rect 4989 34382 5045 34438
rect 5131 34382 5187 34438
rect 5273 34382 5329 34438
rect 5415 34382 5471 34438
rect 5557 34382 5613 34438
rect 5699 34382 5755 34438
rect 5841 34382 5897 34438
rect 5983 34382 6039 34438
rect 6125 34382 6181 34438
rect 6267 34382 6323 34438
rect 6409 34382 6465 34438
rect 6551 34382 6607 34438
rect 6693 34382 6749 34438
rect 6835 34382 6891 34438
rect 6977 34382 7033 34438
rect 7119 34382 7175 34438
rect 7261 34382 7317 34438
rect 7403 34382 7459 34438
rect 7545 34382 7601 34438
rect 7687 34382 7743 34438
rect 7829 34382 7885 34438
rect 7971 34382 8027 34438
rect 8113 34382 8169 34438
rect 8255 34382 8311 34438
rect 8397 34382 8453 34438
rect 8539 34382 8595 34438
rect 8681 34382 8737 34438
rect 8823 34382 8879 34438
rect 8965 34382 9021 34438
rect 9107 34382 9163 34438
rect 9249 34382 9305 34438
rect 9391 34382 9447 34438
rect 9533 34382 9589 34438
rect 9675 34382 9731 34438
rect 9817 34382 9873 34438
rect 9959 34382 10015 34438
rect 10101 34382 10157 34438
rect 10243 34382 10299 34438
rect 10385 34382 10441 34438
rect 10527 34382 10583 34438
rect 10669 34382 10725 34438
rect 10811 34382 10867 34438
rect 10953 34382 11009 34438
rect 11095 34382 11151 34438
rect 11237 34382 11293 34438
rect 11379 34382 11435 34438
rect 11521 34382 11577 34438
rect 11663 34382 11719 34438
rect 11805 34382 11861 34438
rect 11947 34382 12003 34438
rect 12089 34382 12145 34438
rect 12231 34382 12287 34438
rect 12373 34382 12429 34438
rect 12515 34382 12571 34438
rect 12657 34382 12713 34438
rect 12799 34382 12855 34438
rect 12941 34382 12997 34438
rect 13083 34382 13139 34438
rect 13225 34382 13281 34438
rect 13367 34382 13423 34438
rect 13509 34382 13565 34438
rect 13651 34382 13707 34438
rect 13793 34382 13849 34438
rect 13935 34382 13991 34438
rect 14077 34382 14133 34438
rect 14219 34382 14275 34438
rect 14361 34382 14417 34438
rect 14503 34382 14559 34438
rect 14645 34382 14701 34438
rect 14787 34382 14843 34438
rect 161 34240 217 34296
rect 303 34240 359 34296
rect 445 34240 501 34296
rect 587 34240 643 34296
rect 729 34240 785 34296
rect 871 34240 927 34296
rect 1013 34240 1069 34296
rect 1155 34240 1211 34296
rect 1297 34240 1353 34296
rect 1439 34240 1495 34296
rect 1581 34240 1637 34296
rect 1723 34240 1779 34296
rect 1865 34240 1921 34296
rect 2007 34240 2063 34296
rect 2149 34240 2205 34296
rect 2291 34240 2347 34296
rect 2433 34240 2489 34296
rect 2575 34240 2631 34296
rect 2717 34240 2773 34296
rect 2859 34240 2915 34296
rect 3001 34240 3057 34296
rect 3143 34240 3199 34296
rect 3285 34240 3341 34296
rect 3427 34240 3483 34296
rect 3569 34240 3625 34296
rect 3711 34240 3767 34296
rect 3853 34240 3909 34296
rect 3995 34240 4051 34296
rect 4137 34240 4193 34296
rect 4279 34240 4335 34296
rect 4421 34240 4477 34296
rect 4563 34240 4619 34296
rect 4705 34240 4761 34296
rect 4847 34240 4903 34296
rect 4989 34240 5045 34296
rect 5131 34240 5187 34296
rect 5273 34240 5329 34296
rect 5415 34240 5471 34296
rect 5557 34240 5613 34296
rect 5699 34240 5755 34296
rect 5841 34240 5897 34296
rect 5983 34240 6039 34296
rect 6125 34240 6181 34296
rect 6267 34240 6323 34296
rect 6409 34240 6465 34296
rect 6551 34240 6607 34296
rect 6693 34240 6749 34296
rect 6835 34240 6891 34296
rect 6977 34240 7033 34296
rect 7119 34240 7175 34296
rect 7261 34240 7317 34296
rect 7403 34240 7459 34296
rect 7545 34240 7601 34296
rect 7687 34240 7743 34296
rect 7829 34240 7885 34296
rect 7971 34240 8027 34296
rect 8113 34240 8169 34296
rect 8255 34240 8311 34296
rect 8397 34240 8453 34296
rect 8539 34240 8595 34296
rect 8681 34240 8737 34296
rect 8823 34240 8879 34296
rect 8965 34240 9021 34296
rect 9107 34240 9163 34296
rect 9249 34240 9305 34296
rect 9391 34240 9447 34296
rect 9533 34240 9589 34296
rect 9675 34240 9731 34296
rect 9817 34240 9873 34296
rect 9959 34240 10015 34296
rect 10101 34240 10157 34296
rect 10243 34240 10299 34296
rect 10385 34240 10441 34296
rect 10527 34240 10583 34296
rect 10669 34240 10725 34296
rect 10811 34240 10867 34296
rect 10953 34240 11009 34296
rect 11095 34240 11151 34296
rect 11237 34240 11293 34296
rect 11379 34240 11435 34296
rect 11521 34240 11577 34296
rect 11663 34240 11719 34296
rect 11805 34240 11861 34296
rect 11947 34240 12003 34296
rect 12089 34240 12145 34296
rect 12231 34240 12287 34296
rect 12373 34240 12429 34296
rect 12515 34240 12571 34296
rect 12657 34240 12713 34296
rect 12799 34240 12855 34296
rect 12941 34240 12997 34296
rect 13083 34240 13139 34296
rect 13225 34240 13281 34296
rect 13367 34240 13423 34296
rect 13509 34240 13565 34296
rect 13651 34240 13707 34296
rect 13793 34240 13849 34296
rect 13935 34240 13991 34296
rect 14077 34240 14133 34296
rect 14219 34240 14275 34296
rect 14361 34240 14417 34296
rect 14503 34240 14559 34296
rect 14645 34240 14701 34296
rect 14787 34240 14843 34296
rect 161 34098 217 34154
rect 303 34098 359 34154
rect 445 34098 501 34154
rect 587 34098 643 34154
rect 729 34098 785 34154
rect 871 34098 927 34154
rect 1013 34098 1069 34154
rect 1155 34098 1211 34154
rect 1297 34098 1353 34154
rect 1439 34098 1495 34154
rect 1581 34098 1637 34154
rect 1723 34098 1779 34154
rect 1865 34098 1921 34154
rect 2007 34098 2063 34154
rect 2149 34098 2205 34154
rect 2291 34098 2347 34154
rect 2433 34098 2489 34154
rect 2575 34098 2631 34154
rect 2717 34098 2773 34154
rect 2859 34098 2915 34154
rect 3001 34098 3057 34154
rect 3143 34098 3199 34154
rect 3285 34098 3341 34154
rect 3427 34098 3483 34154
rect 3569 34098 3625 34154
rect 3711 34098 3767 34154
rect 3853 34098 3909 34154
rect 3995 34098 4051 34154
rect 4137 34098 4193 34154
rect 4279 34098 4335 34154
rect 4421 34098 4477 34154
rect 4563 34098 4619 34154
rect 4705 34098 4761 34154
rect 4847 34098 4903 34154
rect 4989 34098 5045 34154
rect 5131 34098 5187 34154
rect 5273 34098 5329 34154
rect 5415 34098 5471 34154
rect 5557 34098 5613 34154
rect 5699 34098 5755 34154
rect 5841 34098 5897 34154
rect 5983 34098 6039 34154
rect 6125 34098 6181 34154
rect 6267 34098 6323 34154
rect 6409 34098 6465 34154
rect 6551 34098 6607 34154
rect 6693 34098 6749 34154
rect 6835 34098 6891 34154
rect 6977 34098 7033 34154
rect 7119 34098 7175 34154
rect 7261 34098 7317 34154
rect 7403 34098 7459 34154
rect 7545 34098 7601 34154
rect 7687 34098 7743 34154
rect 7829 34098 7885 34154
rect 7971 34098 8027 34154
rect 8113 34098 8169 34154
rect 8255 34098 8311 34154
rect 8397 34098 8453 34154
rect 8539 34098 8595 34154
rect 8681 34098 8737 34154
rect 8823 34098 8879 34154
rect 8965 34098 9021 34154
rect 9107 34098 9163 34154
rect 9249 34098 9305 34154
rect 9391 34098 9447 34154
rect 9533 34098 9589 34154
rect 9675 34098 9731 34154
rect 9817 34098 9873 34154
rect 9959 34098 10015 34154
rect 10101 34098 10157 34154
rect 10243 34098 10299 34154
rect 10385 34098 10441 34154
rect 10527 34098 10583 34154
rect 10669 34098 10725 34154
rect 10811 34098 10867 34154
rect 10953 34098 11009 34154
rect 11095 34098 11151 34154
rect 11237 34098 11293 34154
rect 11379 34098 11435 34154
rect 11521 34098 11577 34154
rect 11663 34098 11719 34154
rect 11805 34098 11861 34154
rect 11947 34098 12003 34154
rect 12089 34098 12145 34154
rect 12231 34098 12287 34154
rect 12373 34098 12429 34154
rect 12515 34098 12571 34154
rect 12657 34098 12713 34154
rect 12799 34098 12855 34154
rect 12941 34098 12997 34154
rect 13083 34098 13139 34154
rect 13225 34098 13281 34154
rect 13367 34098 13423 34154
rect 13509 34098 13565 34154
rect 13651 34098 13707 34154
rect 13793 34098 13849 34154
rect 13935 34098 13991 34154
rect 14077 34098 14133 34154
rect 14219 34098 14275 34154
rect 14361 34098 14417 34154
rect 14503 34098 14559 34154
rect 14645 34098 14701 34154
rect 14787 34098 14843 34154
rect 161 33956 217 34012
rect 303 33956 359 34012
rect 445 33956 501 34012
rect 587 33956 643 34012
rect 729 33956 785 34012
rect 871 33956 927 34012
rect 1013 33956 1069 34012
rect 1155 33956 1211 34012
rect 1297 33956 1353 34012
rect 1439 33956 1495 34012
rect 1581 33956 1637 34012
rect 1723 33956 1779 34012
rect 1865 33956 1921 34012
rect 2007 33956 2063 34012
rect 2149 33956 2205 34012
rect 2291 33956 2347 34012
rect 2433 33956 2489 34012
rect 2575 33956 2631 34012
rect 2717 33956 2773 34012
rect 2859 33956 2915 34012
rect 3001 33956 3057 34012
rect 3143 33956 3199 34012
rect 3285 33956 3341 34012
rect 3427 33956 3483 34012
rect 3569 33956 3625 34012
rect 3711 33956 3767 34012
rect 3853 33956 3909 34012
rect 3995 33956 4051 34012
rect 4137 33956 4193 34012
rect 4279 33956 4335 34012
rect 4421 33956 4477 34012
rect 4563 33956 4619 34012
rect 4705 33956 4761 34012
rect 4847 33956 4903 34012
rect 4989 33956 5045 34012
rect 5131 33956 5187 34012
rect 5273 33956 5329 34012
rect 5415 33956 5471 34012
rect 5557 33956 5613 34012
rect 5699 33956 5755 34012
rect 5841 33956 5897 34012
rect 5983 33956 6039 34012
rect 6125 33956 6181 34012
rect 6267 33956 6323 34012
rect 6409 33956 6465 34012
rect 6551 33956 6607 34012
rect 6693 33956 6749 34012
rect 6835 33956 6891 34012
rect 6977 33956 7033 34012
rect 7119 33956 7175 34012
rect 7261 33956 7317 34012
rect 7403 33956 7459 34012
rect 7545 33956 7601 34012
rect 7687 33956 7743 34012
rect 7829 33956 7885 34012
rect 7971 33956 8027 34012
rect 8113 33956 8169 34012
rect 8255 33956 8311 34012
rect 8397 33956 8453 34012
rect 8539 33956 8595 34012
rect 8681 33956 8737 34012
rect 8823 33956 8879 34012
rect 8965 33956 9021 34012
rect 9107 33956 9163 34012
rect 9249 33956 9305 34012
rect 9391 33956 9447 34012
rect 9533 33956 9589 34012
rect 9675 33956 9731 34012
rect 9817 33956 9873 34012
rect 9959 33956 10015 34012
rect 10101 33956 10157 34012
rect 10243 33956 10299 34012
rect 10385 33956 10441 34012
rect 10527 33956 10583 34012
rect 10669 33956 10725 34012
rect 10811 33956 10867 34012
rect 10953 33956 11009 34012
rect 11095 33956 11151 34012
rect 11237 33956 11293 34012
rect 11379 33956 11435 34012
rect 11521 33956 11577 34012
rect 11663 33956 11719 34012
rect 11805 33956 11861 34012
rect 11947 33956 12003 34012
rect 12089 33956 12145 34012
rect 12231 33956 12287 34012
rect 12373 33956 12429 34012
rect 12515 33956 12571 34012
rect 12657 33956 12713 34012
rect 12799 33956 12855 34012
rect 12941 33956 12997 34012
rect 13083 33956 13139 34012
rect 13225 33956 13281 34012
rect 13367 33956 13423 34012
rect 13509 33956 13565 34012
rect 13651 33956 13707 34012
rect 13793 33956 13849 34012
rect 13935 33956 13991 34012
rect 14077 33956 14133 34012
rect 14219 33956 14275 34012
rect 14361 33956 14417 34012
rect 14503 33956 14559 34012
rect 14645 33956 14701 34012
rect 14787 33956 14843 34012
rect 161 33814 217 33870
rect 303 33814 359 33870
rect 445 33814 501 33870
rect 587 33814 643 33870
rect 729 33814 785 33870
rect 871 33814 927 33870
rect 1013 33814 1069 33870
rect 1155 33814 1211 33870
rect 1297 33814 1353 33870
rect 1439 33814 1495 33870
rect 1581 33814 1637 33870
rect 1723 33814 1779 33870
rect 1865 33814 1921 33870
rect 2007 33814 2063 33870
rect 2149 33814 2205 33870
rect 2291 33814 2347 33870
rect 2433 33814 2489 33870
rect 2575 33814 2631 33870
rect 2717 33814 2773 33870
rect 2859 33814 2915 33870
rect 3001 33814 3057 33870
rect 3143 33814 3199 33870
rect 3285 33814 3341 33870
rect 3427 33814 3483 33870
rect 3569 33814 3625 33870
rect 3711 33814 3767 33870
rect 3853 33814 3909 33870
rect 3995 33814 4051 33870
rect 4137 33814 4193 33870
rect 4279 33814 4335 33870
rect 4421 33814 4477 33870
rect 4563 33814 4619 33870
rect 4705 33814 4761 33870
rect 4847 33814 4903 33870
rect 4989 33814 5045 33870
rect 5131 33814 5187 33870
rect 5273 33814 5329 33870
rect 5415 33814 5471 33870
rect 5557 33814 5613 33870
rect 5699 33814 5755 33870
rect 5841 33814 5897 33870
rect 5983 33814 6039 33870
rect 6125 33814 6181 33870
rect 6267 33814 6323 33870
rect 6409 33814 6465 33870
rect 6551 33814 6607 33870
rect 6693 33814 6749 33870
rect 6835 33814 6891 33870
rect 6977 33814 7033 33870
rect 7119 33814 7175 33870
rect 7261 33814 7317 33870
rect 7403 33814 7459 33870
rect 7545 33814 7601 33870
rect 7687 33814 7743 33870
rect 7829 33814 7885 33870
rect 7971 33814 8027 33870
rect 8113 33814 8169 33870
rect 8255 33814 8311 33870
rect 8397 33814 8453 33870
rect 8539 33814 8595 33870
rect 8681 33814 8737 33870
rect 8823 33814 8879 33870
rect 8965 33814 9021 33870
rect 9107 33814 9163 33870
rect 9249 33814 9305 33870
rect 9391 33814 9447 33870
rect 9533 33814 9589 33870
rect 9675 33814 9731 33870
rect 9817 33814 9873 33870
rect 9959 33814 10015 33870
rect 10101 33814 10157 33870
rect 10243 33814 10299 33870
rect 10385 33814 10441 33870
rect 10527 33814 10583 33870
rect 10669 33814 10725 33870
rect 10811 33814 10867 33870
rect 10953 33814 11009 33870
rect 11095 33814 11151 33870
rect 11237 33814 11293 33870
rect 11379 33814 11435 33870
rect 11521 33814 11577 33870
rect 11663 33814 11719 33870
rect 11805 33814 11861 33870
rect 11947 33814 12003 33870
rect 12089 33814 12145 33870
rect 12231 33814 12287 33870
rect 12373 33814 12429 33870
rect 12515 33814 12571 33870
rect 12657 33814 12713 33870
rect 12799 33814 12855 33870
rect 12941 33814 12997 33870
rect 13083 33814 13139 33870
rect 13225 33814 13281 33870
rect 13367 33814 13423 33870
rect 13509 33814 13565 33870
rect 13651 33814 13707 33870
rect 13793 33814 13849 33870
rect 13935 33814 13991 33870
rect 14077 33814 14133 33870
rect 14219 33814 14275 33870
rect 14361 33814 14417 33870
rect 14503 33814 14559 33870
rect 14645 33814 14701 33870
rect 14787 33814 14843 33870
rect 161 33672 217 33728
rect 303 33672 359 33728
rect 445 33672 501 33728
rect 587 33672 643 33728
rect 729 33672 785 33728
rect 871 33672 927 33728
rect 1013 33672 1069 33728
rect 1155 33672 1211 33728
rect 1297 33672 1353 33728
rect 1439 33672 1495 33728
rect 1581 33672 1637 33728
rect 1723 33672 1779 33728
rect 1865 33672 1921 33728
rect 2007 33672 2063 33728
rect 2149 33672 2205 33728
rect 2291 33672 2347 33728
rect 2433 33672 2489 33728
rect 2575 33672 2631 33728
rect 2717 33672 2773 33728
rect 2859 33672 2915 33728
rect 3001 33672 3057 33728
rect 3143 33672 3199 33728
rect 3285 33672 3341 33728
rect 3427 33672 3483 33728
rect 3569 33672 3625 33728
rect 3711 33672 3767 33728
rect 3853 33672 3909 33728
rect 3995 33672 4051 33728
rect 4137 33672 4193 33728
rect 4279 33672 4335 33728
rect 4421 33672 4477 33728
rect 4563 33672 4619 33728
rect 4705 33672 4761 33728
rect 4847 33672 4903 33728
rect 4989 33672 5045 33728
rect 5131 33672 5187 33728
rect 5273 33672 5329 33728
rect 5415 33672 5471 33728
rect 5557 33672 5613 33728
rect 5699 33672 5755 33728
rect 5841 33672 5897 33728
rect 5983 33672 6039 33728
rect 6125 33672 6181 33728
rect 6267 33672 6323 33728
rect 6409 33672 6465 33728
rect 6551 33672 6607 33728
rect 6693 33672 6749 33728
rect 6835 33672 6891 33728
rect 6977 33672 7033 33728
rect 7119 33672 7175 33728
rect 7261 33672 7317 33728
rect 7403 33672 7459 33728
rect 7545 33672 7601 33728
rect 7687 33672 7743 33728
rect 7829 33672 7885 33728
rect 7971 33672 8027 33728
rect 8113 33672 8169 33728
rect 8255 33672 8311 33728
rect 8397 33672 8453 33728
rect 8539 33672 8595 33728
rect 8681 33672 8737 33728
rect 8823 33672 8879 33728
rect 8965 33672 9021 33728
rect 9107 33672 9163 33728
rect 9249 33672 9305 33728
rect 9391 33672 9447 33728
rect 9533 33672 9589 33728
rect 9675 33672 9731 33728
rect 9817 33672 9873 33728
rect 9959 33672 10015 33728
rect 10101 33672 10157 33728
rect 10243 33672 10299 33728
rect 10385 33672 10441 33728
rect 10527 33672 10583 33728
rect 10669 33672 10725 33728
rect 10811 33672 10867 33728
rect 10953 33672 11009 33728
rect 11095 33672 11151 33728
rect 11237 33672 11293 33728
rect 11379 33672 11435 33728
rect 11521 33672 11577 33728
rect 11663 33672 11719 33728
rect 11805 33672 11861 33728
rect 11947 33672 12003 33728
rect 12089 33672 12145 33728
rect 12231 33672 12287 33728
rect 12373 33672 12429 33728
rect 12515 33672 12571 33728
rect 12657 33672 12713 33728
rect 12799 33672 12855 33728
rect 12941 33672 12997 33728
rect 13083 33672 13139 33728
rect 13225 33672 13281 33728
rect 13367 33672 13423 33728
rect 13509 33672 13565 33728
rect 13651 33672 13707 33728
rect 13793 33672 13849 33728
rect 13935 33672 13991 33728
rect 14077 33672 14133 33728
rect 14219 33672 14275 33728
rect 14361 33672 14417 33728
rect 14503 33672 14559 33728
rect 14645 33672 14701 33728
rect 14787 33672 14843 33728
rect 161 33530 217 33586
rect 303 33530 359 33586
rect 445 33530 501 33586
rect 587 33530 643 33586
rect 729 33530 785 33586
rect 871 33530 927 33586
rect 1013 33530 1069 33586
rect 1155 33530 1211 33586
rect 1297 33530 1353 33586
rect 1439 33530 1495 33586
rect 1581 33530 1637 33586
rect 1723 33530 1779 33586
rect 1865 33530 1921 33586
rect 2007 33530 2063 33586
rect 2149 33530 2205 33586
rect 2291 33530 2347 33586
rect 2433 33530 2489 33586
rect 2575 33530 2631 33586
rect 2717 33530 2773 33586
rect 2859 33530 2915 33586
rect 3001 33530 3057 33586
rect 3143 33530 3199 33586
rect 3285 33530 3341 33586
rect 3427 33530 3483 33586
rect 3569 33530 3625 33586
rect 3711 33530 3767 33586
rect 3853 33530 3909 33586
rect 3995 33530 4051 33586
rect 4137 33530 4193 33586
rect 4279 33530 4335 33586
rect 4421 33530 4477 33586
rect 4563 33530 4619 33586
rect 4705 33530 4761 33586
rect 4847 33530 4903 33586
rect 4989 33530 5045 33586
rect 5131 33530 5187 33586
rect 5273 33530 5329 33586
rect 5415 33530 5471 33586
rect 5557 33530 5613 33586
rect 5699 33530 5755 33586
rect 5841 33530 5897 33586
rect 5983 33530 6039 33586
rect 6125 33530 6181 33586
rect 6267 33530 6323 33586
rect 6409 33530 6465 33586
rect 6551 33530 6607 33586
rect 6693 33530 6749 33586
rect 6835 33530 6891 33586
rect 6977 33530 7033 33586
rect 7119 33530 7175 33586
rect 7261 33530 7317 33586
rect 7403 33530 7459 33586
rect 7545 33530 7601 33586
rect 7687 33530 7743 33586
rect 7829 33530 7885 33586
rect 7971 33530 8027 33586
rect 8113 33530 8169 33586
rect 8255 33530 8311 33586
rect 8397 33530 8453 33586
rect 8539 33530 8595 33586
rect 8681 33530 8737 33586
rect 8823 33530 8879 33586
rect 8965 33530 9021 33586
rect 9107 33530 9163 33586
rect 9249 33530 9305 33586
rect 9391 33530 9447 33586
rect 9533 33530 9589 33586
rect 9675 33530 9731 33586
rect 9817 33530 9873 33586
rect 9959 33530 10015 33586
rect 10101 33530 10157 33586
rect 10243 33530 10299 33586
rect 10385 33530 10441 33586
rect 10527 33530 10583 33586
rect 10669 33530 10725 33586
rect 10811 33530 10867 33586
rect 10953 33530 11009 33586
rect 11095 33530 11151 33586
rect 11237 33530 11293 33586
rect 11379 33530 11435 33586
rect 11521 33530 11577 33586
rect 11663 33530 11719 33586
rect 11805 33530 11861 33586
rect 11947 33530 12003 33586
rect 12089 33530 12145 33586
rect 12231 33530 12287 33586
rect 12373 33530 12429 33586
rect 12515 33530 12571 33586
rect 12657 33530 12713 33586
rect 12799 33530 12855 33586
rect 12941 33530 12997 33586
rect 13083 33530 13139 33586
rect 13225 33530 13281 33586
rect 13367 33530 13423 33586
rect 13509 33530 13565 33586
rect 13651 33530 13707 33586
rect 13793 33530 13849 33586
rect 13935 33530 13991 33586
rect 14077 33530 14133 33586
rect 14219 33530 14275 33586
rect 14361 33530 14417 33586
rect 14503 33530 14559 33586
rect 14645 33530 14701 33586
rect 14787 33530 14843 33586
rect 161 33388 217 33444
rect 303 33388 359 33444
rect 445 33388 501 33444
rect 587 33388 643 33444
rect 729 33388 785 33444
rect 871 33388 927 33444
rect 1013 33388 1069 33444
rect 1155 33388 1211 33444
rect 1297 33388 1353 33444
rect 1439 33388 1495 33444
rect 1581 33388 1637 33444
rect 1723 33388 1779 33444
rect 1865 33388 1921 33444
rect 2007 33388 2063 33444
rect 2149 33388 2205 33444
rect 2291 33388 2347 33444
rect 2433 33388 2489 33444
rect 2575 33388 2631 33444
rect 2717 33388 2773 33444
rect 2859 33388 2915 33444
rect 3001 33388 3057 33444
rect 3143 33388 3199 33444
rect 3285 33388 3341 33444
rect 3427 33388 3483 33444
rect 3569 33388 3625 33444
rect 3711 33388 3767 33444
rect 3853 33388 3909 33444
rect 3995 33388 4051 33444
rect 4137 33388 4193 33444
rect 4279 33388 4335 33444
rect 4421 33388 4477 33444
rect 4563 33388 4619 33444
rect 4705 33388 4761 33444
rect 4847 33388 4903 33444
rect 4989 33388 5045 33444
rect 5131 33388 5187 33444
rect 5273 33388 5329 33444
rect 5415 33388 5471 33444
rect 5557 33388 5613 33444
rect 5699 33388 5755 33444
rect 5841 33388 5897 33444
rect 5983 33388 6039 33444
rect 6125 33388 6181 33444
rect 6267 33388 6323 33444
rect 6409 33388 6465 33444
rect 6551 33388 6607 33444
rect 6693 33388 6749 33444
rect 6835 33388 6891 33444
rect 6977 33388 7033 33444
rect 7119 33388 7175 33444
rect 7261 33388 7317 33444
rect 7403 33388 7459 33444
rect 7545 33388 7601 33444
rect 7687 33388 7743 33444
rect 7829 33388 7885 33444
rect 7971 33388 8027 33444
rect 8113 33388 8169 33444
rect 8255 33388 8311 33444
rect 8397 33388 8453 33444
rect 8539 33388 8595 33444
rect 8681 33388 8737 33444
rect 8823 33388 8879 33444
rect 8965 33388 9021 33444
rect 9107 33388 9163 33444
rect 9249 33388 9305 33444
rect 9391 33388 9447 33444
rect 9533 33388 9589 33444
rect 9675 33388 9731 33444
rect 9817 33388 9873 33444
rect 9959 33388 10015 33444
rect 10101 33388 10157 33444
rect 10243 33388 10299 33444
rect 10385 33388 10441 33444
rect 10527 33388 10583 33444
rect 10669 33388 10725 33444
rect 10811 33388 10867 33444
rect 10953 33388 11009 33444
rect 11095 33388 11151 33444
rect 11237 33388 11293 33444
rect 11379 33388 11435 33444
rect 11521 33388 11577 33444
rect 11663 33388 11719 33444
rect 11805 33388 11861 33444
rect 11947 33388 12003 33444
rect 12089 33388 12145 33444
rect 12231 33388 12287 33444
rect 12373 33388 12429 33444
rect 12515 33388 12571 33444
rect 12657 33388 12713 33444
rect 12799 33388 12855 33444
rect 12941 33388 12997 33444
rect 13083 33388 13139 33444
rect 13225 33388 13281 33444
rect 13367 33388 13423 33444
rect 13509 33388 13565 33444
rect 13651 33388 13707 33444
rect 13793 33388 13849 33444
rect 13935 33388 13991 33444
rect 14077 33388 14133 33444
rect 14219 33388 14275 33444
rect 14361 33388 14417 33444
rect 14503 33388 14559 33444
rect 14645 33388 14701 33444
rect 14787 33388 14843 33444
rect 161 33246 217 33302
rect 303 33246 359 33302
rect 445 33246 501 33302
rect 587 33246 643 33302
rect 729 33246 785 33302
rect 871 33246 927 33302
rect 1013 33246 1069 33302
rect 1155 33246 1211 33302
rect 1297 33246 1353 33302
rect 1439 33246 1495 33302
rect 1581 33246 1637 33302
rect 1723 33246 1779 33302
rect 1865 33246 1921 33302
rect 2007 33246 2063 33302
rect 2149 33246 2205 33302
rect 2291 33246 2347 33302
rect 2433 33246 2489 33302
rect 2575 33246 2631 33302
rect 2717 33246 2773 33302
rect 2859 33246 2915 33302
rect 3001 33246 3057 33302
rect 3143 33246 3199 33302
rect 3285 33246 3341 33302
rect 3427 33246 3483 33302
rect 3569 33246 3625 33302
rect 3711 33246 3767 33302
rect 3853 33246 3909 33302
rect 3995 33246 4051 33302
rect 4137 33246 4193 33302
rect 4279 33246 4335 33302
rect 4421 33246 4477 33302
rect 4563 33246 4619 33302
rect 4705 33246 4761 33302
rect 4847 33246 4903 33302
rect 4989 33246 5045 33302
rect 5131 33246 5187 33302
rect 5273 33246 5329 33302
rect 5415 33246 5471 33302
rect 5557 33246 5613 33302
rect 5699 33246 5755 33302
rect 5841 33246 5897 33302
rect 5983 33246 6039 33302
rect 6125 33246 6181 33302
rect 6267 33246 6323 33302
rect 6409 33246 6465 33302
rect 6551 33246 6607 33302
rect 6693 33246 6749 33302
rect 6835 33246 6891 33302
rect 6977 33246 7033 33302
rect 7119 33246 7175 33302
rect 7261 33246 7317 33302
rect 7403 33246 7459 33302
rect 7545 33246 7601 33302
rect 7687 33246 7743 33302
rect 7829 33246 7885 33302
rect 7971 33246 8027 33302
rect 8113 33246 8169 33302
rect 8255 33246 8311 33302
rect 8397 33246 8453 33302
rect 8539 33246 8595 33302
rect 8681 33246 8737 33302
rect 8823 33246 8879 33302
rect 8965 33246 9021 33302
rect 9107 33246 9163 33302
rect 9249 33246 9305 33302
rect 9391 33246 9447 33302
rect 9533 33246 9589 33302
rect 9675 33246 9731 33302
rect 9817 33246 9873 33302
rect 9959 33246 10015 33302
rect 10101 33246 10157 33302
rect 10243 33246 10299 33302
rect 10385 33246 10441 33302
rect 10527 33246 10583 33302
rect 10669 33246 10725 33302
rect 10811 33246 10867 33302
rect 10953 33246 11009 33302
rect 11095 33246 11151 33302
rect 11237 33246 11293 33302
rect 11379 33246 11435 33302
rect 11521 33246 11577 33302
rect 11663 33246 11719 33302
rect 11805 33246 11861 33302
rect 11947 33246 12003 33302
rect 12089 33246 12145 33302
rect 12231 33246 12287 33302
rect 12373 33246 12429 33302
rect 12515 33246 12571 33302
rect 12657 33246 12713 33302
rect 12799 33246 12855 33302
rect 12941 33246 12997 33302
rect 13083 33246 13139 33302
rect 13225 33246 13281 33302
rect 13367 33246 13423 33302
rect 13509 33246 13565 33302
rect 13651 33246 13707 33302
rect 13793 33246 13849 33302
rect 13935 33246 13991 33302
rect 14077 33246 14133 33302
rect 14219 33246 14275 33302
rect 14361 33246 14417 33302
rect 14503 33246 14559 33302
rect 14645 33246 14701 33302
rect 14787 33246 14843 33302
rect 161 32885 217 32941
rect 303 32885 359 32941
rect 445 32885 501 32941
rect 587 32885 643 32941
rect 729 32885 785 32941
rect 871 32885 927 32941
rect 1013 32885 1069 32941
rect 1155 32885 1211 32941
rect 1297 32885 1353 32941
rect 1439 32885 1495 32941
rect 1581 32885 1637 32941
rect 1723 32885 1779 32941
rect 1865 32885 1921 32941
rect 2007 32885 2063 32941
rect 2149 32885 2205 32941
rect 2291 32885 2347 32941
rect 2433 32885 2489 32941
rect 2575 32885 2631 32941
rect 2717 32885 2773 32941
rect 2859 32885 2915 32941
rect 3001 32885 3057 32941
rect 3143 32885 3199 32941
rect 3285 32885 3341 32941
rect 3427 32885 3483 32941
rect 3569 32885 3625 32941
rect 3711 32885 3767 32941
rect 3853 32885 3909 32941
rect 3995 32885 4051 32941
rect 4137 32885 4193 32941
rect 4279 32885 4335 32941
rect 4421 32885 4477 32941
rect 4563 32885 4619 32941
rect 4705 32885 4761 32941
rect 4847 32885 4903 32941
rect 4989 32885 5045 32941
rect 5131 32885 5187 32941
rect 5273 32885 5329 32941
rect 5415 32885 5471 32941
rect 5557 32885 5613 32941
rect 5699 32885 5755 32941
rect 5841 32885 5897 32941
rect 5983 32885 6039 32941
rect 6125 32885 6181 32941
rect 6267 32885 6323 32941
rect 6409 32885 6465 32941
rect 6551 32885 6607 32941
rect 6693 32885 6749 32941
rect 6835 32885 6891 32941
rect 6977 32885 7033 32941
rect 7119 32885 7175 32941
rect 7261 32885 7317 32941
rect 7403 32885 7459 32941
rect 7545 32885 7601 32941
rect 7687 32885 7743 32941
rect 7829 32885 7885 32941
rect 7971 32885 8027 32941
rect 8113 32885 8169 32941
rect 8255 32885 8311 32941
rect 8397 32885 8453 32941
rect 8539 32885 8595 32941
rect 8681 32885 8737 32941
rect 8823 32885 8879 32941
rect 8965 32885 9021 32941
rect 9107 32885 9163 32941
rect 9249 32885 9305 32941
rect 9391 32885 9447 32941
rect 9533 32885 9589 32941
rect 9675 32885 9731 32941
rect 9817 32885 9873 32941
rect 9959 32885 10015 32941
rect 10101 32885 10157 32941
rect 10243 32885 10299 32941
rect 10385 32885 10441 32941
rect 10527 32885 10583 32941
rect 10669 32885 10725 32941
rect 10811 32885 10867 32941
rect 10953 32885 11009 32941
rect 11095 32885 11151 32941
rect 11237 32885 11293 32941
rect 11379 32885 11435 32941
rect 11521 32885 11577 32941
rect 11663 32885 11719 32941
rect 11805 32885 11861 32941
rect 11947 32885 12003 32941
rect 12089 32885 12145 32941
rect 12231 32885 12287 32941
rect 12373 32885 12429 32941
rect 12515 32885 12571 32941
rect 12657 32885 12713 32941
rect 12799 32885 12855 32941
rect 12941 32885 12997 32941
rect 13083 32885 13139 32941
rect 13225 32885 13281 32941
rect 13367 32885 13423 32941
rect 13509 32885 13565 32941
rect 13651 32885 13707 32941
rect 13793 32885 13849 32941
rect 13935 32885 13991 32941
rect 14077 32885 14133 32941
rect 14219 32885 14275 32941
rect 14361 32885 14417 32941
rect 14503 32885 14559 32941
rect 14645 32885 14701 32941
rect 14787 32885 14843 32941
rect 161 32743 217 32799
rect 303 32743 359 32799
rect 445 32743 501 32799
rect 587 32743 643 32799
rect 729 32743 785 32799
rect 871 32743 927 32799
rect 1013 32743 1069 32799
rect 1155 32743 1211 32799
rect 1297 32743 1353 32799
rect 1439 32743 1495 32799
rect 1581 32743 1637 32799
rect 1723 32743 1779 32799
rect 1865 32743 1921 32799
rect 2007 32743 2063 32799
rect 2149 32743 2205 32799
rect 2291 32743 2347 32799
rect 2433 32743 2489 32799
rect 2575 32743 2631 32799
rect 2717 32743 2773 32799
rect 2859 32743 2915 32799
rect 3001 32743 3057 32799
rect 3143 32743 3199 32799
rect 3285 32743 3341 32799
rect 3427 32743 3483 32799
rect 3569 32743 3625 32799
rect 3711 32743 3767 32799
rect 3853 32743 3909 32799
rect 3995 32743 4051 32799
rect 4137 32743 4193 32799
rect 4279 32743 4335 32799
rect 4421 32743 4477 32799
rect 4563 32743 4619 32799
rect 4705 32743 4761 32799
rect 4847 32743 4903 32799
rect 4989 32743 5045 32799
rect 5131 32743 5187 32799
rect 5273 32743 5329 32799
rect 5415 32743 5471 32799
rect 5557 32743 5613 32799
rect 5699 32743 5755 32799
rect 5841 32743 5897 32799
rect 5983 32743 6039 32799
rect 6125 32743 6181 32799
rect 6267 32743 6323 32799
rect 6409 32743 6465 32799
rect 6551 32743 6607 32799
rect 6693 32743 6749 32799
rect 6835 32743 6891 32799
rect 6977 32743 7033 32799
rect 7119 32743 7175 32799
rect 7261 32743 7317 32799
rect 7403 32743 7459 32799
rect 7545 32743 7601 32799
rect 7687 32743 7743 32799
rect 7829 32743 7885 32799
rect 7971 32743 8027 32799
rect 8113 32743 8169 32799
rect 8255 32743 8311 32799
rect 8397 32743 8453 32799
rect 8539 32743 8595 32799
rect 8681 32743 8737 32799
rect 8823 32743 8879 32799
rect 8965 32743 9021 32799
rect 9107 32743 9163 32799
rect 9249 32743 9305 32799
rect 9391 32743 9447 32799
rect 9533 32743 9589 32799
rect 9675 32743 9731 32799
rect 9817 32743 9873 32799
rect 9959 32743 10015 32799
rect 10101 32743 10157 32799
rect 10243 32743 10299 32799
rect 10385 32743 10441 32799
rect 10527 32743 10583 32799
rect 10669 32743 10725 32799
rect 10811 32743 10867 32799
rect 10953 32743 11009 32799
rect 11095 32743 11151 32799
rect 11237 32743 11293 32799
rect 11379 32743 11435 32799
rect 11521 32743 11577 32799
rect 11663 32743 11719 32799
rect 11805 32743 11861 32799
rect 11947 32743 12003 32799
rect 12089 32743 12145 32799
rect 12231 32743 12287 32799
rect 12373 32743 12429 32799
rect 12515 32743 12571 32799
rect 12657 32743 12713 32799
rect 12799 32743 12855 32799
rect 12941 32743 12997 32799
rect 13083 32743 13139 32799
rect 13225 32743 13281 32799
rect 13367 32743 13423 32799
rect 13509 32743 13565 32799
rect 13651 32743 13707 32799
rect 13793 32743 13849 32799
rect 13935 32743 13991 32799
rect 14077 32743 14133 32799
rect 14219 32743 14275 32799
rect 14361 32743 14417 32799
rect 14503 32743 14559 32799
rect 14645 32743 14701 32799
rect 14787 32743 14843 32799
rect 161 32601 217 32657
rect 303 32601 359 32657
rect 445 32601 501 32657
rect 587 32601 643 32657
rect 729 32601 785 32657
rect 871 32601 927 32657
rect 1013 32601 1069 32657
rect 1155 32601 1211 32657
rect 1297 32601 1353 32657
rect 1439 32601 1495 32657
rect 1581 32601 1637 32657
rect 1723 32601 1779 32657
rect 1865 32601 1921 32657
rect 2007 32601 2063 32657
rect 2149 32601 2205 32657
rect 2291 32601 2347 32657
rect 2433 32601 2489 32657
rect 2575 32601 2631 32657
rect 2717 32601 2773 32657
rect 2859 32601 2915 32657
rect 3001 32601 3057 32657
rect 3143 32601 3199 32657
rect 3285 32601 3341 32657
rect 3427 32601 3483 32657
rect 3569 32601 3625 32657
rect 3711 32601 3767 32657
rect 3853 32601 3909 32657
rect 3995 32601 4051 32657
rect 4137 32601 4193 32657
rect 4279 32601 4335 32657
rect 4421 32601 4477 32657
rect 4563 32601 4619 32657
rect 4705 32601 4761 32657
rect 4847 32601 4903 32657
rect 4989 32601 5045 32657
rect 5131 32601 5187 32657
rect 5273 32601 5329 32657
rect 5415 32601 5471 32657
rect 5557 32601 5613 32657
rect 5699 32601 5755 32657
rect 5841 32601 5897 32657
rect 5983 32601 6039 32657
rect 6125 32601 6181 32657
rect 6267 32601 6323 32657
rect 6409 32601 6465 32657
rect 6551 32601 6607 32657
rect 6693 32601 6749 32657
rect 6835 32601 6891 32657
rect 6977 32601 7033 32657
rect 7119 32601 7175 32657
rect 7261 32601 7317 32657
rect 7403 32601 7459 32657
rect 7545 32601 7601 32657
rect 7687 32601 7743 32657
rect 7829 32601 7885 32657
rect 7971 32601 8027 32657
rect 8113 32601 8169 32657
rect 8255 32601 8311 32657
rect 8397 32601 8453 32657
rect 8539 32601 8595 32657
rect 8681 32601 8737 32657
rect 8823 32601 8879 32657
rect 8965 32601 9021 32657
rect 9107 32601 9163 32657
rect 9249 32601 9305 32657
rect 9391 32601 9447 32657
rect 9533 32601 9589 32657
rect 9675 32601 9731 32657
rect 9817 32601 9873 32657
rect 9959 32601 10015 32657
rect 10101 32601 10157 32657
rect 10243 32601 10299 32657
rect 10385 32601 10441 32657
rect 10527 32601 10583 32657
rect 10669 32601 10725 32657
rect 10811 32601 10867 32657
rect 10953 32601 11009 32657
rect 11095 32601 11151 32657
rect 11237 32601 11293 32657
rect 11379 32601 11435 32657
rect 11521 32601 11577 32657
rect 11663 32601 11719 32657
rect 11805 32601 11861 32657
rect 11947 32601 12003 32657
rect 12089 32601 12145 32657
rect 12231 32601 12287 32657
rect 12373 32601 12429 32657
rect 12515 32601 12571 32657
rect 12657 32601 12713 32657
rect 12799 32601 12855 32657
rect 12941 32601 12997 32657
rect 13083 32601 13139 32657
rect 13225 32601 13281 32657
rect 13367 32601 13423 32657
rect 13509 32601 13565 32657
rect 13651 32601 13707 32657
rect 13793 32601 13849 32657
rect 13935 32601 13991 32657
rect 14077 32601 14133 32657
rect 14219 32601 14275 32657
rect 14361 32601 14417 32657
rect 14503 32601 14559 32657
rect 14645 32601 14701 32657
rect 14787 32601 14843 32657
rect 161 32459 217 32515
rect 303 32459 359 32515
rect 445 32459 501 32515
rect 587 32459 643 32515
rect 729 32459 785 32515
rect 871 32459 927 32515
rect 1013 32459 1069 32515
rect 1155 32459 1211 32515
rect 1297 32459 1353 32515
rect 1439 32459 1495 32515
rect 1581 32459 1637 32515
rect 1723 32459 1779 32515
rect 1865 32459 1921 32515
rect 2007 32459 2063 32515
rect 2149 32459 2205 32515
rect 2291 32459 2347 32515
rect 2433 32459 2489 32515
rect 2575 32459 2631 32515
rect 2717 32459 2773 32515
rect 2859 32459 2915 32515
rect 3001 32459 3057 32515
rect 3143 32459 3199 32515
rect 3285 32459 3341 32515
rect 3427 32459 3483 32515
rect 3569 32459 3625 32515
rect 3711 32459 3767 32515
rect 3853 32459 3909 32515
rect 3995 32459 4051 32515
rect 4137 32459 4193 32515
rect 4279 32459 4335 32515
rect 4421 32459 4477 32515
rect 4563 32459 4619 32515
rect 4705 32459 4761 32515
rect 4847 32459 4903 32515
rect 4989 32459 5045 32515
rect 5131 32459 5187 32515
rect 5273 32459 5329 32515
rect 5415 32459 5471 32515
rect 5557 32459 5613 32515
rect 5699 32459 5755 32515
rect 5841 32459 5897 32515
rect 5983 32459 6039 32515
rect 6125 32459 6181 32515
rect 6267 32459 6323 32515
rect 6409 32459 6465 32515
rect 6551 32459 6607 32515
rect 6693 32459 6749 32515
rect 6835 32459 6891 32515
rect 6977 32459 7033 32515
rect 7119 32459 7175 32515
rect 7261 32459 7317 32515
rect 7403 32459 7459 32515
rect 7545 32459 7601 32515
rect 7687 32459 7743 32515
rect 7829 32459 7885 32515
rect 7971 32459 8027 32515
rect 8113 32459 8169 32515
rect 8255 32459 8311 32515
rect 8397 32459 8453 32515
rect 8539 32459 8595 32515
rect 8681 32459 8737 32515
rect 8823 32459 8879 32515
rect 8965 32459 9021 32515
rect 9107 32459 9163 32515
rect 9249 32459 9305 32515
rect 9391 32459 9447 32515
rect 9533 32459 9589 32515
rect 9675 32459 9731 32515
rect 9817 32459 9873 32515
rect 9959 32459 10015 32515
rect 10101 32459 10157 32515
rect 10243 32459 10299 32515
rect 10385 32459 10441 32515
rect 10527 32459 10583 32515
rect 10669 32459 10725 32515
rect 10811 32459 10867 32515
rect 10953 32459 11009 32515
rect 11095 32459 11151 32515
rect 11237 32459 11293 32515
rect 11379 32459 11435 32515
rect 11521 32459 11577 32515
rect 11663 32459 11719 32515
rect 11805 32459 11861 32515
rect 11947 32459 12003 32515
rect 12089 32459 12145 32515
rect 12231 32459 12287 32515
rect 12373 32459 12429 32515
rect 12515 32459 12571 32515
rect 12657 32459 12713 32515
rect 12799 32459 12855 32515
rect 12941 32459 12997 32515
rect 13083 32459 13139 32515
rect 13225 32459 13281 32515
rect 13367 32459 13423 32515
rect 13509 32459 13565 32515
rect 13651 32459 13707 32515
rect 13793 32459 13849 32515
rect 13935 32459 13991 32515
rect 14077 32459 14133 32515
rect 14219 32459 14275 32515
rect 14361 32459 14417 32515
rect 14503 32459 14559 32515
rect 14645 32459 14701 32515
rect 14787 32459 14843 32515
rect 161 32317 217 32373
rect 303 32317 359 32373
rect 445 32317 501 32373
rect 587 32317 643 32373
rect 729 32317 785 32373
rect 871 32317 927 32373
rect 1013 32317 1069 32373
rect 1155 32317 1211 32373
rect 1297 32317 1353 32373
rect 1439 32317 1495 32373
rect 1581 32317 1637 32373
rect 1723 32317 1779 32373
rect 1865 32317 1921 32373
rect 2007 32317 2063 32373
rect 2149 32317 2205 32373
rect 2291 32317 2347 32373
rect 2433 32317 2489 32373
rect 2575 32317 2631 32373
rect 2717 32317 2773 32373
rect 2859 32317 2915 32373
rect 3001 32317 3057 32373
rect 3143 32317 3199 32373
rect 3285 32317 3341 32373
rect 3427 32317 3483 32373
rect 3569 32317 3625 32373
rect 3711 32317 3767 32373
rect 3853 32317 3909 32373
rect 3995 32317 4051 32373
rect 4137 32317 4193 32373
rect 4279 32317 4335 32373
rect 4421 32317 4477 32373
rect 4563 32317 4619 32373
rect 4705 32317 4761 32373
rect 4847 32317 4903 32373
rect 4989 32317 5045 32373
rect 5131 32317 5187 32373
rect 5273 32317 5329 32373
rect 5415 32317 5471 32373
rect 5557 32317 5613 32373
rect 5699 32317 5755 32373
rect 5841 32317 5897 32373
rect 5983 32317 6039 32373
rect 6125 32317 6181 32373
rect 6267 32317 6323 32373
rect 6409 32317 6465 32373
rect 6551 32317 6607 32373
rect 6693 32317 6749 32373
rect 6835 32317 6891 32373
rect 6977 32317 7033 32373
rect 7119 32317 7175 32373
rect 7261 32317 7317 32373
rect 7403 32317 7459 32373
rect 7545 32317 7601 32373
rect 7687 32317 7743 32373
rect 7829 32317 7885 32373
rect 7971 32317 8027 32373
rect 8113 32317 8169 32373
rect 8255 32317 8311 32373
rect 8397 32317 8453 32373
rect 8539 32317 8595 32373
rect 8681 32317 8737 32373
rect 8823 32317 8879 32373
rect 8965 32317 9021 32373
rect 9107 32317 9163 32373
rect 9249 32317 9305 32373
rect 9391 32317 9447 32373
rect 9533 32317 9589 32373
rect 9675 32317 9731 32373
rect 9817 32317 9873 32373
rect 9959 32317 10015 32373
rect 10101 32317 10157 32373
rect 10243 32317 10299 32373
rect 10385 32317 10441 32373
rect 10527 32317 10583 32373
rect 10669 32317 10725 32373
rect 10811 32317 10867 32373
rect 10953 32317 11009 32373
rect 11095 32317 11151 32373
rect 11237 32317 11293 32373
rect 11379 32317 11435 32373
rect 11521 32317 11577 32373
rect 11663 32317 11719 32373
rect 11805 32317 11861 32373
rect 11947 32317 12003 32373
rect 12089 32317 12145 32373
rect 12231 32317 12287 32373
rect 12373 32317 12429 32373
rect 12515 32317 12571 32373
rect 12657 32317 12713 32373
rect 12799 32317 12855 32373
rect 12941 32317 12997 32373
rect 13083 32317 13139 32373
rect 13225 32317 13281 32373
rect 13367 32317 13423 32373
rect 13509 32317 13565 32373
rect 13651 32317 13707 32373
rect 13793 32317 13849 32373
rect 13935 32317 13991 32373
rect 14077 32317 14133 32373
rect 14219 32317 14275 32373
rect 14361 32317 14417 32373
rect 14503 32317 14559 32373
rect 14645 32317 14701 32373
rect 14787 32317 14843 32373
rect 161 32175 217 32231
rect 303 32175 359 32231
rect 445 32175 501 32231
rect 587 32175 643 32231
rect 729 32175 785 32231
rect 871 32175 927 32231
rect 1013 32175 1069 32231
rect 1155 32175 1211 32231
rect 1297 32175 1353 32231
rect 1439 32175 1495 32231
rect 1581 32175 1637 32231
rect 1723 32175 1779 32231
rect 1865 32175 1921 32231
rect 2007 32175 2063 32231
rect 2149 32175 2205 32231
rect 2291 32175 2347 32231
rect 2433 32175 2489 32231
rect 2575 32175 2631 32231
rect 2717 32175 2773 32231
rect 2859 32175 2915 32231
rect 3001 32175 3057 32231
rect 3143 32175 3199 32231
rect 3285 32175 3341 32231
rect 3427 32175 3483 32231
rect 3569 32175 3625 32231
rect 3711 32175 3767 32231
rect 3853 32175 3909 32231
rect 3995 32175 4051 32231
rect 4137 32175 4193 32231
rect 4279 32175 4335 32231
rect 4421 32175 4477 32231
rect 4563 32175 4619 32231
rect 4705 32175 4761 32231
rect 4847 32175 4903 32231
rect 4989 32175 5045 32231
rect 5131 32175 5187 32231
rect 5273 32175 5329 32231
rect 5415 32175 5471 32231
rect 5557 32175 5613 32231
rect 5699 32175 5755 32231
rect 5841 32175 5897 32231
rect 5983 32175 6039 32231
rect 6125 32175 6181 32231
rect 6267 32175 6323 32231
rect 6409 32175 6465 32231
rect 6551 32175 6607 32231
rect 6693 32175 6749 32231
rect 6835 32175 6891 32231
rect 6977 32175 7033 32231
rect 7119 32175 7175 32231
rect 7261 32175 7317 32231
rect 7403 32175 7459 32231
rect 7545 32175 7601 32231
rect 7687 32175 7743 32231
rect 7829 32175 7885 32231
rect 7971 32175 8027 32231
rect 8113 32175 8169 32231
rect 8255 32175 8311 32231
rect 8397 32175 8453 32231
rect 8539 32175 8595 32231
rect 8681 32175 8737 32231
rect 8823 32175 8879 32231
rect 8965 32175 9021 32231
rect 9107 32175 9163 32231
rect 9249 32175 9305 32231
rect 9391 32175 9447 32231
rect 9533 32175 9589 32231
rect 9675 32175 9731 32231
rect 9817 32175 9873 32231
rect 9959 32175 10015 32231
rect 10101 32175 10157 32231
rect 10243 32175 10299 32231
rect 10385 32175 10441 32231
rect 10527 32175 10583 32231
rect 10669 32175 10725 32231
rect 10811 32175 10867 32231
rect 10953 32175 11009 32231
rect 11095 32175 11151 32231
rect 11237 32175 11293 32231
rect 11379 32175 11435 32231
rect 11521 32175 11577 32231
rect 11663 32175 11719 32231
rect 11805 32175 11861 32231
rect 11947 32175 12003 32231
rect 12089 32175 12145 32231
rect 12231 32175 12287 32231
rect 12373 32175 12429 32231
rect 12515 32175 12571 32231
rect 12657 32175 12713 32231
rect 12799 32175 12855 32231
rect 12941 32175 12997 32231
rect 13083 32175 13139 32231
rect 13225 32175 13281 32231
rect 13367 32175 13423 32231
rect 13509 32175 13565 32231
rect 13651 32175 13707 32231
rect 13793 32175 13849 32231
rect 13935 32175 13991 32231
rect 14077 32175 14133 32231
rect 14219 32175 14275 32231
rect 14361 32175 14417 32231
rect 14503 32175 14559 32231
rect 14645 32175 14701 32231
rect 14787 32175 14843 32231
rect 161 32033 217 32089
rect 303 32033 359 32089
rect 445 32033 501 32089
rect 587 32033 643 32089
rect 729 32033 785 32089
rect 871 32033 927 32089
rect 1013 32033 1069 32089
rect 1155 32033 1211 32089
rect 1297 32033 1353 32089
rect 1439 32033 1495 32089
rect 1581 32033 1637 32089
rect 1723 32033 1779 32089
rect 1865 32033 1921 32089
rect 2007 32033 2063 32089
rect 2149 32033 2205 32089
rect 2291 32033 2347 32089
rect 2433 32033 2489 32089
rect 2575 32033 2631 32089
rect 2717 32033 2773 32089
rect 2859 32033 2915 32089
rect 3001 32033 3057 32089
rect 3143 32033 3199 32089
rect 3285 32033 3341 32089
rect 3427 32033 3483 32089
rect 3569 32033 3625 32089
rect 3711 32033 3767 32089
rect 3853 32033 3909 32089
rect 3995 32033 4051 32089
rect 4137 32033 4193 32089
rect 4279 32033 4335 32089
rect 4421 32033 4477 32089
rect 4563 32033 4619 32089
rect 4705 32033 4761 32089
rect 4847 32033 4903 32089
rect 4989 32033 5045 32089
rect 5131 32033 5187 32089
rect 5273 32033 5329 32089
rect 5415 32033 5471 32089
rect 5557 32033 5613 32089
rect 5699 32033 5755 32089
rect 5841 32033 5897 32089
rect 5983 32033 6039 32089
rect 6125 32033 6181 32089
rect 6267 32033 6323 32089
rect 6409 32033 6465 32089
rect 6551 32033 6607 32089
rect 6693 32033 6749 32089
rect 6835 32033 6891 32089
rect 6977 32033 7033 32089
rect 7119 32033 7175 32089
rect 7261 32033 7317 32089
rect 7403 32033 7459 32089
rect 7545 32033 7601 32089
rect 7687 32033 7743 32089
rect 7829 32033 7885 32089
rect 7971 32033 8027 32089
rect 8113 32033 8169 32089
rect 8255 32033 8311 32089
rect 8397 32033 8453 32089
rect 8539 32033 8595 32089
rect 8681 32033 8737 32089
rect 8823 32033 8879 32089
rect 8965 32033 9021 32089
rect 9107 32033 9163 32089
rect 9249 32033 9305 32089
rect 9391 32033 9447 32089
rect 9533 32033 9589 32089
rect 9675 32033 9731 32089
rect 9817 32033 9873 32089
rect 9959 32033 10015 32089
rect 10101 32033 10157 32089
rect 10243 32033 10299 32089
rect 10385 32033 10441 32089
rect 10527 32033 10583 32089
rect 10669 32033 10725 32089
rect 10811 32033 10867 32089
rect 10953 32033 11009 32089
rect 11095 32033 11151 32089
rect 11237 32033 11293 32089
rect 11379 32033 11435 32089
rect 11521 32033 11577 32089
rect 11663 32033 11719 32089
rect 11805 32033 11861 32089
rect 11947 32033 12003 32089
rect 12089 32033 12145 32089
rect 12231 32033 12287 32089
rect 12373 32033 12429 32089
rect 12515 32033 12571 32089
rect 12657 32033 12713 32089
rect 12799 32033 12855 32089
rect 12941 32033 12997 32089
rect 13083 32033 13139 32089
rect 13225 32033 13281 32089
rect 13367 32033 13423 32089
rect 13509 32033 13565 32089
rect 13651 32033 13707 32089
rect 13793 32033 13849 32089
rect 13935 32033 13991 32089
rect 14077 32033 14133 32089
rect 14219 32033 14275 32089
rect 14361 32033 14417 32089
rect 14503 32033 14559 32089
rect 14645 32033 14701 32089
rect 14787 32033 14843 32089
rect 161 31891 217 31947
rect 303 31891 359 31947
rect 445 31891 501 31947
rect 587 31891 643 31947
rect 729 31891 785 31947
rect 871 31891 927 31947
rect 1013 31891 1069 31947
rect 1155 31891 1211 31947
rect 1297 31891 1353 31947
rect 1439 31891 1495 31947
rect 1581 31891 1637 31947
rect 1723 31891 1779 31947
rect 1865 31891 1921 31947
rect 2007 31891 2063 31947
rect 2149 31891 2205 31947
rect 2291 31891 2347 31947
rect 2433 31891 2489 31947
rect 2575 31891 2631 31947
rect 2717 31891 2773 31947
rect 2859 31891 2915 31947
rect 3001 31891 3057 31947
rect 3143 31891 3199 31947
rect 3285 31891 3341 31947
rect 3427 31891 3483 31947
rect 3569 31891 3625 31947
rect 3711 31891 3767 31947
rect 3853 31891 3909 31947
rect 3995 31891 4051 31947
rect 4137 31891 4193 31947
rect 4279 31891 4335 31947
rect 4421 31891 4477 31947
rect 4563 31891 4619 31947
rect 4705 31891 4761 31947
rect 4847 31891 4903 31947
rect 4989 31891 5045 31947
rect 5131 31891 5187 31947
rect 5273 31891 5329 31947
rect 5415 31891 5471 31947
rect 5557 31891 5613 31947
rect 5699 31891 5755 31947
rect 5841 31891 5897 31947
rect 5983 31891 6039 31947
rect 6125 31891 6181 31947
rect 6267 31891 6323 31947
rect 6409 31891 6465 31947
rect 6551 31891 6607 31947
rect 6693 31891 6749 31947
rect 6835 31891 6891 31947
rect 6977 31891 7033 31947
rect 7119 31891 7175 31947
rect 7261 31891 7317 31947
rect 7403 31891 7459 31947
rect 7545 31891 7601 31947
rect 7687 31891 7743 31947
rect 7829 31891 7885 31947
rect 7971 31891 8027 31947
rect 8113 31891 8169 31947
rect 8255 31891 8311 31947
rect 8397 31891 8453 31947
rect 8539 31891 8595 31947
rect 8681 31891 8737 31947
rect 8823 31891 8879 31947
rect 8965 31891 9021 31947
rect 9107 31891 9163 31947
rect 9249 31891 9305 31947
rect 9391 31891 9447 31947
rect 9533 31891 9589 31947
rect 9675 31891 9731 31947
rect 9817 31891 9873 31947
rect 9959 31891 10015 31947
rect 10101 31891 10157 31947
rect 10243 31891 10299 31947
rect 10385 31891 10441 31947
rect 10527 31891 10583 31947
rect 10669 31891 10725 31947
rect 10811 31891 10867 31947
rect 10953 31891 11009 31947
rect 11095 31891 11151 31947
rect 11237 31891 11293 31947
rect 11379 31891 11435 31947
rect 11521 31891 11577 31947
rect 11663 31891 11719 31947
rect 11805 31891 11861 31947
rect 11947 31891 12003 31947
rect 12089 31891 12145 31947
rect 12231 31891 12287 31947
rect 12373 31891 12429 31947
rect 12515 31891 12571 31947
rect 12657 31891 12713 31947
rect 12799 31891 12855 31947
rect 12941 31891 12997 31947
rect 13083 31891 13139 31947
rect 13225 31891 13281 31947
rect 13367 31891 13423 31947
rect 13509 31891 13565 31947
rect 13651 31891 13707 31947
rect 13793 31891 13849 31947
rect 13935 31891 13991 31947
rect 14077 31891 14133 31947
rect 14219 31891 14275 31947
rect 14361 31891 14417 31947
rect 14503 31891 14559 31947
rect 14645 31891 14701 31947
rect 14787 31891 14843 31947
rect 161 31749 217 31805
rect 303 31749 359 31805
rect 445 31749 501 31805
rect 587 31749 643 31805
rect 729 31749 785 31805
rect 871 31749 927 31805
rect 1013 31749 1069 31805
rect 1155 31749 1211 31805
rect 1297 31749 1353 31805
rect 1439 31749 1495 31805
rect 1581 31749 1637 31805
rect 1723 31749 1779 31805
rect 1865 31749 1921 31805
rect 2007 31749 2063 31805
rect 2149 31749 2205 31805
rect 2291 31749 2347 31805
rect 2433 31749 2489 31805
rect 2575 31749 2631 31805
rect 2717 31749 2773 31805
rect 2859 31749 2915 31805
rect 3001 31749 3057 31805
rect 3143 31749 3199 31805
rect 3285 31749 3341 31805
rect 3427 31749 3483 31805
rect 3569 31749 3625 31805
rect 3711 31749 3767 31805
rect 3853 31749 3909 31805
rect 3995 31749 4051 31805
rect 4137 31749 4193 31805
rect 4279 31749 4335 31805
rect 4421 31749 4477 31805
rect 4563 31749 4619 31805
rect 4705 31749 4761 31805
rect 4847 31749 4903 31805
rect 4989 31749 5045 31805
rect 5131 31749 5187 31805
rect 5273 31749 5329 31805
rect 5415 31749 5471 31805
rect 5557 31749 5613 31805
rect 5699 31749 5755 31805
rect 5841 31749 5897 31805
rect 5983 31749 6039 31805
rect 6125 31749 6181 31805
rect 6267 31749 6323 31805
rect 6409 31749 6465 31805
rect 6551 31749 6607 31805
rect 6693 31749 6749 31805
rect 6835 31749 6891 31805
rect 6977 31749 7033 31805
rect 7119 31749 7175 31805
rect 7261 31749 7317 31805
rect 7403 31749 7459 31805
rect 7545 31749 7601 31805
rect 7687 31749 7743 31805
rect 7829 31749 7885 31805
rect 7971 31749 8027 31805
rect 8113 31749 8169 31805
rect 8255 31749 8311 31805
rect 8397 31749 8453 31805
rect 8539 31749 8595 31805
rect 8681 31749 8737 31805
rect 8823 31749 8879 31805
rect 8965 31749 9021 31805
rect 9107 31749 9163 31805
rect 9249 31749 9305 31805
rect 9391 31749 9447 31805
rect 9533 31749 9589 31805
rect 9675 31749 9731 31805
rect 9817 31749 9873 31805
rect 9959 31749 10015 31805
rect 10101 31749 10157 31805
rect 10243 31749 10299 31805
rect 10385 31749 10441 31805
rect 10527 31749 10583 31805
rect 10669 31749 10725 31805
rect 10811 31749 10867 31805
rect 10953 31749 11009 31805
rect 11095 31749 11151 31805
rect 11237 31749 11293 31805
rect 11379 31749 11435 31805
rect 11521 31749 11577 31805
rect 11663 31749 11719 31805
rect 11805 31749 11861 31805
rect 11947 31749 12003 31805
rect 12089 31749 12145 31805
rect 12231 31749 12287 31805
rect 12373 31749 12429 31805
rect 12515 31749 12571 31805
rect 12657 31749 12713 31805
rect 12799 31749 12855 31805
rect 12941 31749 12997 31805
rect 13083 31749 13139 31805
rect 13225 31749 13281 31805
rect 13367 31749 13423 31805
rect 13509 31749 13565 31805
rect 13651 31749 13707 31805
rect 13793 31749 13849 31805
rect 13935 31749 13991 31805
rect 14077 31749 14133 31805
rect 14219 31749 14275 31805
rect 14361 31749 14417 31805
rect 14503 31749 14559 31805
rect 14645 31749 14701 31805
rect 14787 31749 14843 31805
rect 161 31607 217 31663
rect 303 31607 359 31663
rect 445 31607 501 31663
rect 587 31607 643 31663
rect 729 31607 785 31663
rect 871 31607 927 31663
rect 1013 31607 1069 31663
rect 1155 31607 1211 31663
rect 1297 31607 1353 31663
rect 1439 31607 1495 31663
rect 1581 31607 1637 31663
rect 1723 31607 1779 31663
rect 1865 31607 1921 31663
rect 2007 31607 2063 31663
rect 2149 31607 2205 31663
rect 2291 31607 2347 31663
rect 2433 31607 2489 31663
rect 2575 31607 2631 31663
rect 2717 31607 2773 31663
rect 2859 31607 2915 31663
rect 3001 31607 3057 31663
rect 3143 31607 3199 31663
rect 3285 31607 3341 31663
rect 3427 31607 3483 31663
rect 3569 31607 3625 31663
rect 3711 31607 3767 31663
rect 3853 31607 3909 31663
rect 3995 31607 4051 31663
rect 4137 31607 4193 31663
rect 4279 31607 4335 31663
rect 4421 31607 4477 31663
rect 4563 31607 4619 31663
rect 4705 31607 4761 31663
rect 4847 31607 4903 31663
rect 4989 31607 5045 31663
rect 5131 31607 5187 31663
rect 5273 31607 5329 31663
rect 5415 31607 5471 31663
rect 5557 31607 5613 31663
rect 5699 31607 5755 31663
rect 5841 31607 5897 31663
rect 5983 31607 6039 31663
rect 6125 31607 6181 31663
rect 6267 31607 6323 31663
rect 6409 31607 6465 31663
rect 6551 31607 6607 31663
rect 6693 31607 6749 31663
rect 6835 31607 6891 31663
rect 6977 31607 7033 31663
rect 7119 31607 7175 31663
rect 7261 31607 7317 31663
rect 7403 31607 7459 31663
rect 7545 31607 7601 31663
rect 7687 31607 7743 31663
rect 7829 31607 7885 31663
rect 7971 31607 8027 31663
rect 8113 31607 8169 31663
rect 8255 31607 8311 31663
rect 8397 31607 8453 31663
rect 8539 31607 8595 31663
rect 8681 31607 8737 31663
rect 8823 31607 8879 31663
rect 8965 31607 9021 31663
rect 9107 31607 9163 31663
rect 9249 31607 9305 31663
rect 9391 31607 9447 31663
rect 9533 31607 9589 31663
rect 9675 31607 9731 31663
rect 9817 31607 9873 31663
rect 9959 31607 10015 31663
rect 10101 31607 10157 31663
rect 10243 31607 10299 31663
rect 10385 31607 10441 31663
rect 10527 31607 10583 31663
rect 10669 31607 10725 31663
rect 10811 31607 10867 31663
rect 10953 31607 11009 31663
rect 11095 31607 11151 31663
rect 11237 31607 11293 31663
rect 11379 31607 11435 31663
rect 11521 31607 11577 31663
rect 11663 31607 11719 31663
rect 11805 31607 11861 31663
rect 11947 31607 12003 31663
rect 12089 31607 12145 31663
rect 12231 31607 12287 31663
rect 12373 31607 12429 31663
rect 12515 31607 12571 31663
rect 12657 31607 12713 31663
rect 12799 31607 12855 31663
rect 12941 31607 12997 31663
rect 13083 31607 13139 31663
rect 13225 31607 13281 31663
rect 13367 31607 13423 31663
rect 13509 31607 13565 31663
rect 13651 31607 13707 31663
rect 13793 31607 13849 31663
rect 13935 31607 13991 31663
rect 14077 31607 14133 31663
rect 14219 31607 14275 31663
rect 14361 31607 14417 31663
rect 14503 31607 14559 31663
rect 14645 31607 14701 31663
rect 14787 31607 14843 31663
rect 161 31465 217 31521
rect 303 31465 359 31521
rect 445 31465 501 31521
rect 587 31465 643 31521
rect 729 31465 785 31521
rect 871 31465 927 31521
rect 1013 31465 1069 31521
rect 1155 31465 1211 31521
rect 1297 31465 1353 31521
rect 1439 31465 1495 31521
rect 1581 31465 1637 31521
rect 1723 31465 1779 31521
rect 1865 31465 1921 31521
rect 2007 31465 2063 31521
rect 2149 31465 2205 31521
rect 2291 31465 2347 31521
rect 2433 31465 2489 31521
rect 2575 31465 2631 31521
rect 2717 31465 2773 31521
rect 2859 31465 2915 31521
rect 3001 31465 3057 31521
rect 3143 31465 3199 31521
rect 3285 31465 3341 31521
rect 3427 31465 3483 31521
rect 3569 31465 3625 31521
rect 3711 31465 3767 31521
rect 3853 31465 3909 31521
rect 3995 31465 4051 31521
rect 4137 31465 4193 31521
rect 4279 31465 4335 31521
rect 4421 31465 4477 31521
rect 4563 31465 4619 31521
rect 4705 31465 4761 31521
rect 4847 31465 4903 31521
rect 4989 31465 5045 31521
rect 5131 31465 5187 31521
rect 5273 31465 5329 31521
rect 5415 31465 5471 31521
rect 5557 31465 5613 31521
rect 5699 31465 5755 31521
rect 5841 31465 5897 31521
rect 5983 31465 6039 31521
rect 6125 31465 6181 31521
rect 6267 31465 6323 31521
rect 6409 31465 6465 31521
rect 6551 31465 6607 31521
rect 6693 31465 6749 31521
rect 6835 31465 6891 31521
rect 6977 31465 7033 31521
rect 7119 31465 7175 31521
rect 7261 31465 7317 31521
rect 7403 31465 7459 31521
rect 7545 31465 7601 31521
rect 7687 31465 7743 31521
rect 7829 31465 7885 31521
rect 7971 31465 8027 31521
rect 8113 31465 8169 31521
rect 8255 31465 8311 31521
rect 8397 31465 8453 31521
rect 8539 31465 8595 31521
rect 8681 31465 8737 31521
rect 8823 31465 8879 31521
rect 8965 31465 9021 31521
rect 9107 31465 9163 31521
rect 9249 31465 9305 31521
rect 9391 31465 9447 31521
rect 9533 31465 9589 31521
rect 9675 31465 9731 31521
rect 9817 31465 9873 31521
rect 9959 31465 10015 31521
rect 10101 31465 10157 31521
rect 10243 31465 10299 31521
rect 10385 31465 10441 31521
rect 10527 31465 10583 31521
rect 10669 31465 10725 31521
rect 10811 31465 10867 31521
rect 10953 31465 11009 31521
rect 11095 31465 11151 31521
rect 11237 31465 11293 31521
rect 11379 31465 11435 31521
rect 11521 31465 11577 31521
rect 11663 31465 11719 31521
rect 11805 31465 11861 31521
rect 11947 31465 12003 31521
rect 12089 31465 12145 31521
rect 12231 31465 12287 31521
rect 12373 31465 12429 31521
rect 12515 31465 12571 31521
rect 12657 31465 12713 31521
rect 12799 31465 12855 31521
rect 12941 31465 12997 31521
rect 13083 31465 13139 31521
rect 13225 31465 13281 31521
rect 13367 31465 13423 31521
rect 13509 31465 13565 31521
rect 13651 31465 13707 31521
rect 13793 31465 13849 31521
rect 13935 31465 13991 31521
rect 14077 31465 14133 31521
rect 14219 31465 14275 31521
rect 14361 31465 14417 31521
rect 14503 31465 14559 31521
rect 14645 31465 14701 31521
rect 14787 31465 14843 31521
rect 161 31323 217 31379
rect 303 31323 359 31379
rect 445 31323 501 31379
rect 587 31323 643 31379
rect 729 31323 785 31379
rect 871 31323 927 31379
rect 1013 31323 1069 31379
rect 1155 31323 1211 31379
rect 1297 31323 1353 31379
rect 1439 31323 1495 31379
rect 1581 31323 1637 31379
rect 1723 31323 1779 31379
rect 1865 31323 1921 31379
rect 2007 31323 2063 31379
rect 2149 31323 2205 31379
rect 2291 31323 2347 31379
rect 2433 31323 2489 31379
rect 2575 31323 2631 31379
rect 2717 31323 2773 31379
rect 2859 31323 2915 31379
rect 3001 31323 3057 31379
rect 3143 31323 3199 31379
rect 3285 31323 3341 31379
rect 3427 31323 3483 31379
rect 3569 31323 3625 31379
rect 3711 31323 3767 31379
rect 3853 31323 3909 31379
rect 3995 31323 4051 31379
rect 4137 31323 4193 31379
rect 4279 31323 4335 31379
rect 4421 31323 4477 31379
rect 4563 31323 4619 31379
rect 4705 31323 4761 31379
rect 4847 31323 4903 31379
rect 4989 31323 5045 31379
rect 5131 31323 5187 31379
rect 5273 31323 5329 31379
rect 5415 31323 5471 31379
rect 5557 31323 5613 31379
rect 5699 31323 5755 31379
rect 5841 31323 5897 31379
rect 5983 31323 6039 31379
rect 6125 31323 6181 31379
rect 6267 31323 6323 31379
rect 6409 31323 6465 31379
rect 6551 31323 6607 31379
rect 6693 31323 6749 31379
rect 6835 31323 6891 31379
rect 6977 31323 7033 31379
rect 7119 31323 7175 31379
rect 7261 31323 7317 31379
rect 7403 31323 7459 31379
rect 7545 31323 7601 31379
rect 7687 31323 7743 31379
rect 7829 31323 7885 31379
rect 7971 31323 8027 31379
rect 8113 31323 8169 31379
rect 8255 31323 8311 31379
rect 8397 31323 8453 31379
rect 8539 31323 8595 31379
rect 8681 31323 8737 31379
rect 8823 31323 8879 31379
rect 8965 31323 9021 31379
rect 9107 31323 9163 31379
rect 9249 31323 9305 31379
rect 9391 31323 9447 31379
rect 9533 31323 9589 31379
rect 9675 31323 9731 31379
rect 9817 31323 9873 31379
rect 9959 31323 10015 31379
rect 10101 31323 10157 31379
rect 10243 31323 10299 31379
rect 10385 31323 10441 31379
rect 10527 31323 10583 31379
rect 10669 31323 10725 31379
rect 10811 31323 10867 31379
rect 10953 31323 11009 31379
rect 11095 31323 11151 31379
rect 11237 31323 11293 31379
rect 11379 31323 11435 31379
rect 11521 31323 11577 31379
rect 11663 31323 11719 31379
rect 11805 31323 11861 31379
rect 11947 31323 12003 31379
rect 12089 31323 12145 31379
rect 12231 31323 12287 31379
rect 12373 31323 12429 31379
rect 12515 31323 12571 31379
rect 12657 31323 12713 31379
rect 12799 31323 12855 31379
rect 12941 31323 12997 31379
rect 13083 31323 13139 31379
rect 13225 31323 13281 31379
rect 13367 31323 13423 31379
rect 13509 31323 13565 31379
rect 13651 31323 13707 31379
rect 13793 31323 13849 31379
rect 13935 31323 13991 31379
rect 14077 31323 14133 31379
rect 14219 31323 14275 31379
rect 14361 31323 14417 31379
rect 14503 31323 14559 31379
rect 14645 31323 14701 31379
rect 14787 31323 14843 31379
rect 161 31181 217 31237
rect 303 31181 359 31237
rect 445 31181 501 31237
rect 587 31181 643 31237
rect 729 31181 785 31237
rect 871 31181 927 31237
rect 1013 31181 1069 31237
rect 1155 31181 1211 31237
rect 1297 31181 1353 31237
rect 1439 31181 1495 31237
rect 1581 31181 1637 31237
rect 1723 31181 1779 31237
rect 1865 31181 1921 31237
rect 2007 31181 2063 31237
rect 2149 31181 2205 31237
rect 2291 31181 2347 31237
rect 2433 31181 2489 31237
rect 2575 31181 2631 31237
rect 2717 31181 2773 31237
rect 2859 31181 2915 31237
rect 3001 31181 3057 31237
rect 3143 31181 3199 31237
rect 3285 31181 3341 31237
rect 3427 31181 3483 31237
rect 3569 31181 3625 31237
rect 3711 31181 3767 31237
rect 3853 31181 3909 31237
rect 3995 31181 4051 31237
rect 4137 31181 4193 31237
rect 4279 31181 4335 31237
rect 4421 31181 4477 31237
rect 4563 31181 4619 31237
rect 4705 31181 4761 31237
rect 4847 31181 4903 31237
rect 4989 31181 5045 31237
rect 5131 31181 5187 31237
rect 5273 31181 5329 31237
rect 5415 31181 5471 31237
rect 5557 31181 5613 31237
rect 5699 31181 5755 31237
rect 5841 31181 5897 31237
rect 5983 31181 6039 31237
rect 6125 31181 6181 31237
rect 6267 31181 6323 31237
rect 6409 31181 6465 31237
rect 6551 31181 6607 31237
rect 6693 31181 6749 31237
rect 6835 31181 6891 31237
rect 6977 31181 7033 31237
rect 7119 31181 7175 31237
rect 7261 31181 7317 31237
rect 7403 31181 7459 31237
rect 7545 31181 7601 31237
rect 7687 31181 7743 31237
rect 7829 31181 7885 31237
rect 7971 31181 8027 31237
rect 8113 31181 8169 31237
rect 8255 31181 8311 31237
rect 8397 31181 8453 31237
rect 8539 31181 8595 31237
rect 8681 31181 8737 31237
rect 8823 31181 8879 31237
rect 8965 31181 9021 31237
rect 9107 31181 9163 31237
rect 9249 31181 9305 31237
rect 9391 31181 9447 31237
rect 9533 31181 9589 31237
rect 9675 31181 9731 31237
rect 9817 31181 9873 31237
rect 9959 31181 10015 31237
rect 10101 31181 10157 31237
rect 10243 31181 10299 31237
rect 10385 31181 10441 31237
rect 10527 31181 10583 31237
rect 10669 31181 10725 31237
rect 10811 31181 10867 31237
rect 10953 31181 11009 31237
rect 11095 31181 11151 31237
rect 11237 31181 11293 31237
rect 11379 31181 11435 31237
rect 11521 31181 11577 31237
rect 11663 31181 11719 31237
rect 11805 31181 11861 31237
rect 11947 31181 12003 31237
rect 12089 31181 12145 31237
rect 12231 31181 12287 31237
rect 12373 31181 12429 31237
rect 12515 31181 12571 31237
rect 12657 31181 12713 31237
rect 12799 31181 12855 31237
rect 12941 31181 12997 31237
rect 13083 31181 13139 31237
rect 13225 31181 13281 31237
rect 13367 31181 13423 31237
rect 13509 31181 13565 31237
rect 13651 31181 13707 31237
rect 13793 31181 13849 31237
rect 13935 31181 13991 31237
rect 14077 31181 14133 31237
rect 14219 31181 14275 31237
rect 14361 31181 14417 31237
rect 14503 31181 14559 31237
rect 14645 31181 14701 31237
rect 14787 31181 14843 31237
rect 161 31039 217 31095
rect 303 31039 359 31095
rect 445 31039 501 31095
rect 587 31039 643 31095
rect 729 31039 785 31095
rect 871 31039 927 31095
rect 1013 31039 1069 31095
rect 1155 31039 1211 31095
rect 1297 31039 1353 31095
rect 1439 31039 1495 31095
rect 1581 31039 1637 31095
rect 1723 31039 1779 31095
rect 1865 31039 1921 31095
rect 2007 31039 2063 31095
rect 2149 31039 2205 31095
rect 2291 31039 2347 31095
rect 2433 31039 2489 31095
rect 2575 31039 2631 31095
rect 2717 31039 2773 31095
rect 2859 31039 2915 31095
rect 3001 31039 3057 31095
rect 3143 31039 3199 31095
rect 3285 31039 3341 31095
rect 3427 31039 3483 31095
rect 3569 31039 3625 31095
rect 3711 31039 3767 31095
rect 3853 31039 3909 31095
rect 3995 31039 4051 31095
rect 4137 31039 4193 31095
rect 4279 31039 4335 31095
rect 4421 31039 4477 31095
rect 4563 31039 4619 31095
rect 4705 31039 4761 31095
rect 4847 31039 4903 31095
rect 4989 31039 5045 31095
rect 5131 31039 5187 31095
rect 5273 31039 5329 31095
rect 5415 31039 5471 31095
rect 5557 31039 5613 31095
rect 5699 31039 5755 31095
rect 5841 31039 5897 31095
rect 5983 31039 6039 31095
rect 6125 31039 6181 31095
rect 6267 31039 6323 31095
rect 6409 31039 6465 31095
rect 6551 31039 6607 31095
rect 6693 31039 6749 31095
rect 6835 31039 6891 31095
rect 6977 31039 7033 31095
rect 7119 31039 7175 31095
rect 7261 31039 7317 31095
rect 7403 31039 7459 31095
rect 7545 31039 7601 31095
rect 7687 31039 7743 31095
rect 7829 31039 7885 31095
rect 7971 31039 8027 31095
rect 8113 31039 8169 31095
rect 8255 31039 8311 31095
rect 8397 31039 8453 31095
rect 8539 31039 8595 31095
rect 8681 31039 8737 31095
rect 8823 31039 8879 31095
rect 8965 31039 9021 31095
rect 9107 31039 9163 31095
rect 9249 31039 9305 31095
rect 9391 31039 9447 31095
rect 9533 31039 9589 31095
rect 9675 31039 9731 31095
rect 9817 31039 9873 31095
rect 9959 31039 10015 31095
rect 10101 31039 10157 31095
rect 10243 31039 10299 31095
rect 10385 31039 10441 31095
rect 10527 31039 10583 31095
rect 10669 31039 10725 31095
rect 10811 31039 10867 31095
rect 10953 31039 11009 31095
rect 11095 31039 11151 31095
rect 11237 31039 11293 31095
rect 11379 31039 11435 31095
rect 11521 31039 11577 31095
rect 11663 31039 11719 31095
rect 11805 31039 11861 31095
rect 11947 31039 12003 31095
rect 12089 31039 12145 31095
rect 12231 31039 12287 31095
rect 12373 31039 12429 31095
rect 12515 31039 12571 31095
rect 12657 31039 12713 31095
rect 12799 31039 12855 31095
rect 12941 31039 12997 31095
rect 13083 31039 13139 31095
rect 13225 31039 13281 31095
rect 13367 31039 13423 31095
rect 13509 31039 13565 31095
rect 13651 31039 13707 31095
rect 13793 31039 13849 31095
rect 13935 31039 13991 31095
rect 14077 31039 14133 31095
rect 14219 31039 14275 31095
rect 14361 31039 14417 31095
rect 14503 31039 14559 31095
rect 14645 31039 14701 31095
rect 14787 31039 14843 31095
rect 161 30897 217 30953
rect 303 30897 359 30953
rect 445 30897 501 30953
rect 587 30897 643 30953
rect 729 30897 785 30953
rect 871 30897 927 30953
rect 1013 30897 1069 30953
rect 1155 30897 1211 30953
rect 1297 30897 1353 30953
rect 1439 30897 1495 30953
rect 1581 30897 1637 30953
rect 1723 30897 1779 30953
rect 1865 30897 1921 30953
rect 2007 30897 2063 30953
rect 2149 30897 2205 30953
rect 2291 30897 2347 30953
rect 2433 30897 2489 30953
rect 2575 30897 2631 30953
rect 2717 30897 2773 30953
rect 2859 30897 2915 30953
rect 3001 30897 3057 30953
rect 3143 30897 3199 30953
rect 3285 30897 3341 30953
rect 3427 30897 3483 30953
rect 3569 30897 3625 30953
rect 3711 30897 3767 30953
rect 3853 30897 3909 30953
rect 3995 30897 4051 30953
rect 4137 30897 4193 30953
rect 4279 30897 4335 30953
rect 4421 30897 4477 30953
rect 4563 30897 4619 30953
rect 4705 30897 4761 30953
rect 4847 30897 4903 30953
rect 4989 30897 5045 30953
rect 5131 30897 5187 30953
rect 5273 30897 5329 30953
rect 5415 30897 5471 30953
rect 5557 30897 5613 30953
rect 5699 30897 5755 30953
rect 5841 30897 5897 30953
rect 5983 30897 6039 30953
rect 6125 30897 6181 30953
rect 6267 30897 6323 30953
rect 6409 30897 6465 30953
rect 6551 30897 6607 30953
rect 6693 30897 6749 30953
rect 6835 30897 6891 30953
rect 6977 30897 7033 30953
rect 7119 30897 7175 30953
rect 7261 30897 7317 30953
rect 7403 30897 7459 30953
rect 7545 30897 7601 30953
rect 7687 30897 7743 30953
rect 7829 30897 7885 30953
rect 7971 30897 8027 30953
rect 8113 30897 8169 30953
rect 8255 30897 8311 30953
rect 8397 30897 8453 30953
rect 8539 30897 8595 30953
rect 8681 30897 8737 30953
rect 8823 30897 8879 30953
rect 8965 30897 9021 30953
rect 9107 30897 9163 30953
rect 9249 30897 9305 30953
rect 9391 30897 9447 30953
rect 9533 30897 9589 30953
rect 9675 30897 9731 30953
rect 9817 30897 9873 30953
rect 9959 30897 10015 30953
rect 10101 30897 10157 30953
rect 10243 30897 10299 30953
rect 10385 30897 10441 30953
rect 10527 30897 10583 30953
rect 10669 30897 10725 30953
rect 10811 30897 10867 30953
rect 10953 30897 11009 30953
rect 11095 30897 11151 30953
rect 11237 30897 11293 30953
rect 11379 30897 11435 30953
rect 11521 30897 11577 30953
rect 11663 30897 11719 30953
rect 11805 30897 11861 30953
rect 11947 30897 12003 30953
rect 12089 30897 12145 30953
rect 12231 30897 12287 30953
rect 12373 30897 12429 30953
rect 12515 30897 12571 30953
rect 12657 30897 12713 30953
rect 12799 30897 12855 30953
rect 12941 30897 12997 30953
rect 13083 30897 13139 30953
rect 13225 30897 13281 30953
rect 13367 30897 13423 30953
rect 13509 30897 13565 30953
rect 13651 30897 13707 30953
rect 13793 30897 13849 30953
rect 13935 30897 13991 30953
rect 14077 30897 14133 30953
rect 14219 30897 14275 30953
rect 14361 30897 14417 30953
rect 14503 30897 14559 30953
rect 14645 30897 14701 30953
rect 14787 30897 14843 30953
rect 161 30755 217 30811
rect 303 30755 359 30811
rect 445 30755 501 30811
rect 587 30755 643 30811
rect 729 30755 785 30811
rect 871 30755 927 30811
rect 1013 30755 1069 30811
rect 1155 30755 1211 30811
rect 1297 30755 1353 30811
rect 1439 30755 1495 30811
rect 1581 30755 1637 30811
rect 1723 30755 1779 30811
rect 1865 30755 1921 30811
rect 2007 30755 2063 30811
rect 2149 30755 2205 30811
rect 2291 30755 2347 30811
rect 2433 30755 2489 30811
rect 2575 30755 2631 30811
rect 2717 30755 2773 30811
rect 2859 30755 2915 30811
rect 3001 30755 3057 30811
rect 3143 30755 3199 30811
rect 3285 30755 3341 30811
rect 3427 30755 3483 30811
rect 3569 30755 3625 30811
rect 3711 30755 3767 30811
rect 3853 30755 3909 30811
rect 3995 30755 4051 30811
rect 4137 30755 4193 30811
rect 4279 30755 4335 30811
rect 4421 30755 4477 30811
rect 4563 30755 4619 30811
rect 4705 30755 4761 30811
rect 4847 30755 4903 30811
rect 4989 30755 5045 30811
rect 5131 30755 5187 30811
rect 5273 30755 5329 30811
rect 5415 30755 5471 30811
rect 5557 30755 5613 30811
rect 5699 30755 5755 30811
rect 5841 30755 5897 30811
rect 5983 30755 6039 30811
rect 6125 30755 6181 30811
rect 6267 30755 6323 30811
rect 6409 30755 6465 30811
rect 6551 30755 6607 30811
rect 6693 30755 6749 30811
rect 6835 30755 6891 30811
rect 6977 30755 7033 30811
rect 7119 30755 7175 30811
rect 7261 30755 7317 30811
rect 7403 30755 7459 30811
rect 7545 30755 7601 30811
rect 7687 30755 7743 30811
rect 7829 30755 7885 30811
rect 7971 30755 8027 30811
rect 8113 30755 8169 30811
rect 8255 30755 8311 30811
rect 8397 30755 8453 30811
rect 8539 30755 8595 30811
rect 8681 30755 8737 30811
rect 8823 30755 8879 30811
rect 8965 30755 9021 30811
rect 9107 30755 9163 30811
rect 9249 30755 9305 30811
rect 9391 30755 9447 30811
rect 9533 30755 9589 30811
rect 9675 30755 9731 30811
rect 9817 30755 9873 30811
rect 9959 30755 10015 30811
rect 10101 30755 10157 30811
rect 10243 30755 10299 30811
rect 10385 30755 10441 30811
rect 10527 30755 10583 30811
rect 10669 30755 10725 30811
rect 10811 30755 10867 30811
rect 10953 30755 11009 30811
rect 11095 30755 11151 30811
rect 11237 30755 11293 30811
rect 11379 30755 11435 30811
rect 11521 30755 11577 30811
rect 11663 30755 11719 30811
rect 11805 30755 11861 30811
rect 11947 30755 12003 30811
rect 12089 30755 12145 30811
rect 12231 30755 12287 30811
rect 12373 30755 12429 30811
rect 12515 30755 12571 30811
rect 12657 30755 12713 30811
rect 12799 30755 12855 30811
rect 12941 30755 12997 30811
rect 13083 30755 13139 30811
rect 13225 30755 13281 30811
rect 13367 30755 13423 30811
rect 13509 30755 13565 30811
rect 13651 30755 13707 30811
rect 13793 30755 13849 30811
rect 13935 30755 13991 30811
rect 14077 30755 14133 30811
rect 14219 30755 14275 30811
rect 14361 30755 14417 30811
rect 14503 30755 14559 30811
rect 14645 30755 14701 30811
rect 14787 30755 14843 30811
rect 161 30613 217 30669
rect 303 30613 359 30669
rect 445 30613 501 30669
rect 587 30613 643 30669
rect 729 30613 785 30669
rect 871 30613 927 30669
rect 1013 30613 1069 30669
rect 1155 30613 1211 30669
rect 1297 30613 1353 30669
rect 1439 30613 1495 30669
rect 1581 30613 1637 30669
rect 1723 30613 1779 30669
rect 1865 30613 1921 30669
rect 2007 30613 2063 30669
rect 2149 30613 2205 30669
rect 2291 30613 2347 30669
rect 2433 30613 2489 30669
rect 2575 30613 2631 30669
rect 2717 30613 2773 30669
rect 2859 30613 2915 30669
rect 3001 30613 3057 30669
rect 3143 30613 3199 30669
rect 3285 30613 3341 30669
rect 3427 30613 3483 30669
rect 3569 30613 3625 30669
rect 3711 30613 3767 30669
rect 3853 30613 3909 30669
rect 3995 30613 4051 30669
rect 4137 30613 4193 30669
rect 4279 30613 4335 30669
rect 4421 30613 4477 30669
rect 4563 30613 4619 30669
rect 4705 30613 4761 30669
rect 4847 30613 4903 30669
rect 4989 30613 5045 30669
rect 5131 30613 5187 30669
rect 5273 30613 5329 30669
rect 5415 30613 5471 30669
rect 5557 30613 5613 30669
rect 5699 30613 5755 30669
rect 5841 30613 5897 30669
rect 5983 30613 6039 30669
rect 6125 30613 6181 30669
rect 6267 30613 6323 30669
rect 6409 30613 6465 30669
rect 6551 30613 6607 30669
rect 6693 30613 6749 30669
rect 6835 30613 6891 30669
rect 6977 30613 7033 30669
rect 7119 30613 7175 30669
rect 7261 30613 7317 30669
rect 7403 30613 7459 30669
rect 7545 30613 7601 30669
rect 7687 30613 7743 30669
rect 7829 30613 7885 30669
rect 7971 30613 8027 30669
rect 8113 30613 8169 30669
rect 8255 30613 8311 30669
rect 8397 30613 8453 30669
rect 8539 30613 8595 30669
rect 8681 30613 8737 30669
rect 8823 30613 8879 30669
rect 8965 30613 9021 30669
rect 9107 30613 9163 30669
rect 9249 30613 9305 30669
rect 9391 30613 9447 30669
rect 9533 30613 9589 30669
rect 9675 30613 9731 30669
rect 9817 30613 9873 30669
rect 9959 30613 10015 30669
rect 10101 30613 10157 30669
rect 10243 30613 10299 30669
rect 10385 30613 10441 30669
rect 10527 30613 10583 30669
rect 10669 30613 10725 30669
rect 10811 30613 10867 30669
rect 10953 30613 11009 30669
rect 11095 30613 11151 30669
rect 11237 30613 11293 30669
rect 11379 30613 11435 30669
rect 11521 30613 11577 30669
rect 11663 30613 11719 30669
rect 11805 30613 11861 30669
rect 11947 30613 12003 30669
rect 12089 30613 12145 30669
rect 12231 30613 12287 30669
rect 12373 30613 12429 30669
rect 12515 30613 12571 30669
rect 12657 30613 12713 30669
rect 12799 30613 12855 30669
rect 12941 30613 12997 30669
rect 13083 30613 13139 30669
rect 13225 30613 13281 30669
rect 13367 30613 13423 30669
rect 13509 30613 13565 30669
rect 13651 30613 13707 30669
rect 13793 30613 13849 30669
rect 13935 30613 13991 30669
rect 14077 30613 14133 30669
rect 14219 30613 14275 30669
rect 14361 30613 14417 30669
rect 14503 30613 14559 30669
rect 14645 30613 14701 30669
rect 14787 30613 14843 30669
rect 161 30471 217 30527
rect 303 30471 359 30527
rect 445 30471 501 30527
rect 587 30471 643 30527
rect 729 30471 785 30527
rect 871 30471 927 30527
rect 1013 30471 1069 30527
rect 1155 30471 1211 30527
rect 1297 30471 1353 30527
rect 1439 30471 1495 30527
rect 1581 30471 1637 30527
rect 1723 30471 1779 30527
rect 1865 30471 1921 30527
rect 2007 30471 2063 30527
rect 2149 30471 2205 30527
rect 2291 30471 2347 30527
rect 2433 30471 2489 30527
rect 2575 30471 2631 30527
rect 2717 30471 2773 30527
rect 2859 30471 2915 30527
rect 3001 30471 3057 30527
rect 3143 30471 3199 30527
rect 3285 30471 3341 30527
rect 3427 30471 3483 30527
rect 3569 30471 3625 30527
rect 3711 30471 3767 30527
rect 3853 30471 3909 30527
rect 3995 30471 4051 30527
rect 4137 30471 4193 30527
rect 4279 30471 4335 30527
rect 4421 30471 4477 30527
rect 4563 30471 4619 30527
rect 4705 30471 4761 30527
rect 4847 30471 4903 30527
rect 4989 30471 5045 30527
rect 5131 30471 5187 30527
rect 5273 30471 5329 30527
rect 5415 30471 5471 30527
rect 5557 30471 5613 30527
rect 5699 30471 5755 30527
rect 5841 30471 5897 30527
rect 5983 30471 6039 30527
rect 6125 30471 6181 30527
rect 6267 30471 6323 30527
rect 6409 30471 6465 30527
rect 6551 30471 6607 30527
rect 6693 30471 6749 30527
rect 6835 30471 6891 30527
rect 6977 30471 7033 30527
rect 7119 30471 7175 30527
rect 7261 30471 7317 30527
rect 7403 30471 7459 30527
rect 7545 30471 7601 30527
rect 7687 30471 7743 30527
rect 7829 30471 7885 30527
rect 7971 30471 8027 30527
rect 8113 30471 8169 30527
rect 8255 30471 8311 30527
rect 8397 30471 8453 30527
rect 8539 30471 8595 30527
rect 8681 30471 8737 30527
rect 8823 30471 8879 30527
rect 8965 30471 9021 30527
rect 9107 30471 9163 30527
rect 9249 30471 9305 30527
rect 9391 30471 9447 30527
rect 9533 30471 9589 30527
rect 9675 30471 9731 30527
rect 9817 30471 9873 30527
rect 9959 30471 10015 30527
rect 10101 30471 10157 30527
rect 10243 30471 10299 30527
rect 10385 30471 10441 30527
rect 10527 30471 10583 30527
rect 10669 30471 10725 30527
rect 10811 30471 10867 30527
rect 10953 30471 11009 30527
rect 11095 30471 11151 30527
rect 11237 30471 11293 30527
rect 11379 30471 11435 30527
rect 11521 30471 11577 30527
rect 11663 30471 11719 30527
rect 11805 30471 11861 30527
rect 11947 30471 12003 30527
rect 12089 30471 12145 30527
rect 12231 30471 12287 30527
rect 12373 30471 12429 30527
rect 12515 30471 12571 30527
rect 12657 30471 12713 30527
rect 12799 30471 12855 30527
rect 12941 30471 12997 30527
rect 13083 30471 13139 30527
rect 13225 30471 13281 30527
rect 13367 30471 13423 30527
rect 13509 30471 13565 30527
rect 13651 30471 13707 30527
rect 13793 30471 13849 30527
rect 13935 30471 13991 30527
rect 14077 30471 14133 30527
rect 14219 30471 14275 30527
rect 14361 30471 14417 30527
rect 14503 30471 14559 30527
rect 14645 30471 14701 30527
rect 14787 30471 14843 30527
rect 161 30329 217 30385
rect 303 30329 359 30385
rect 445 30329 501 30385
rect 587 30329 643 30385
rect 729 30329 785 30385
rect 871 30329 927 30385
rect 1013 30329 1069 30385
rect 1155 30329 1211 30385
rect 1297 30329 1353 30385
rect 1439 30329 1495 30385
rect 1581 30329 1637 30385
rect 1723 30329 1779 30385
rect 1865 30329 1921 30385
rect 2007 30329 2063 30385
rect 2149 30329 2205 30385
rect 2291 30329 2347 30385
rect 2433 30329 2489 30385
rect 2575 30329 2631 30385
rect 2717 30329 2773 30385
rect 2859 30329 2915 30385
rect 3001 30329 3057 30385
rect 3143 30329 3199 30385
rect 3285 30329 3341 30385
rect 3427 30329 3483 30385
rect 3569 30329 3625 30385
rect 3711 30329 3767 30385
rect 3853 30329 3909 30385
rect 3995 30329 4051 30385
rect 4137 30329 4193 30385
rect 4279 30329 4335 30385
rect 4421 30329 4477 30385
rect 4563 30329 4619 30385
rect 4705 30329 4761 30385
rect 4847 30329 4903 30385
rect 4989 30329 5045 30385
rect 5131 30329 5187 30385
rect 5273 30329 5329 30385
rect 5415 30329 5471 30385
rect 5557 30329 5613 30385
rect 5699 30329 5755 30385
rect 5841 30329 5897 30385
rect 5983 30329 6039 30385
rect 6125 30329 6181 30385
rect 6267 30329 6323 30385
rect 6409 30329 6465 30385
rect 6551 30329 6607 30385
rect 6693 30329 6749 30385
rect 6835 30329 6891 30385
rect 6977 30329 7033 30385
rect 7119 30329 7175 30385
rect 7261 30329 7317 30385
rect 7403 30329 7459 30385
rect 7545 30329 7601 30385
rect 7687 30329 7743 30385
rect 7829 30329 7885 30385
rect 7971 30329 8027 30385
rect 8113 30329 8169 30385
rect 8255 30329 8311 30385
rect 8397 30329 8453 30385
rect 8539 30329 8595 30385
rect 8681 30329 8737 30385
rect 8823 30329 8879 30385
rect 8965 30329 9021 30385
rect 9107 30329 9163 30385
rect 9249 30329 9305 30385
rect 9391 30329 9447 30385
rect 9533 30329 9589 30385
rect 9675 30329 9731 30385
rect 9817 30329 9873 30385
rect 9959 30329 10015 30385
rect 10101 30329 10157 30385
rect 10243 30329 10299 30385
rect 10385 30329 10441 30385
rect 10527 30329 10583 30385
rect 10669 30329 10725 30385
rect 10811 30329 10867 30385
rect 10953 30329 11009 30385
rect 11095 30329 11151 30385
rect 11237 30329 11293 30385
rect 11379 30329 11435 30385
rect 11521 30329 11577 30385
rect 11663 30329 11719 30385
rect 11805 30329 11861 30385
rect 11947 30329 12003 30385
rect 12089 30329 12145 30385
rect 12231 30329 12287 30385
rect 12373 30329 12429 30385
rect 12515 30329 12571 30385
rect 12657 30329 12713 30385
rect 12799 30329 12855 30385
rect 12941 30329 12997 30385
rect 13083 30329 13139 30385
rect 13225 30329 13281 30385
rect 13367 30329 13423 30385
rect 13509 30329 13565 30385
rect 13651 30329 13707 30385
rect 13793 30329 13849 30385
rect 13935 30329 13991 30385
rect 14077 30329 14133 30385
rect 14219 30329 14275 30385
rect 14361 30329 14417 30385
rect 14503 30329 14559 30385
rect 14645 30329 14701 30385
rect 14787 30329 14843 30385
rect 161 30187 217 30243
rect 303 30187 359 30243
rect 445 30187 501 30243
rect 587 30187 643 30243
rect 729 30187 785 30243
rect 871 30187 927 30243
rect 1013 30187 1069 30243
rect 1155 30187 1211 30243
rect 1297 30187 1353 30243
rect 1439 30187 1495 30243
rect 1581 30187 1637 30243
rect 1723 30187 1779 30243
rect 1865 30187 1921 30243
rect 2007 30187 2063 30243
rect 2149 30187 2205 30243
rect 2291 30187 2347 30243
rect 2433 30187 2489 30243
rect 2575 30187 2631 30243
rect 2717 30187 2773 30243
rect 2859 30187 2915 30243
rect 3001 30187 3057 30243
rect 3143 30187 3199 30243
rect 3285 30187 3341 30243
rect 3427 30187 3483 30243
rect 3569 30187 3625 30243
rect 3711 30187 3767 30243
rect 3853 30187 3909 30243
rect 3995 30187 4051 30243
rect 4137 30187 4193 30243
rect 4279 30187 4335 30243
rect 4421 30187 4477 30243
rect 4563 30187 4619 30243
rect 4705 30187 4761 30243
rect 4847 30187 4903 30243
rect 4989 30187 5045 30243
rect 5131 30187 5187 30243
rect 5273 30187 5329 30243
rect 5415 30187 5471 30243
rect 5557 30187 5613 30243
rect 5699 30187 5755 30243
rect 5841 30187 5897 30243
rect 5983 30187 6039 30243
rect 6125 30187 6181 30243
rect 6267 30187 6323 30243
rect 6409 30187 6465 30243
rect 6551 30187 6607 30243
rect 6693 30187 6749 30243
rect 6835 30187 6891 30243
rect 6977 30187 7033 30243
rect 7119 30187 7175 30243
rect 7261 30187 7317 30243
rect 7403 30187 7459 30243
rect 7545 30187 7601 30243
rect 7687 30187 7743 30243
rect 7829 30187 7885 30243
rect 7971 30187 8027 30243
rect 8113 30187 8169 30243
rect 8255 30187 8311 30243
rect 8397 30187 8453 30243
rect 8539 30187 8595 30243
rect 8681 30187 8737 30243
rect 8823 30187 8879 30243
rect 8965 30187 9021 30243
rect 9107 30187 9163 30243
rect 9249 30187 9305 30243
rect 9391 30187 9447 30243
rect 9533 30187 9589 30243
rect 9675 30187 9731 30243
rect 9817 30187 9873 30243
rect 9959 30187 10015 30243
rect 10101 30187 10157 30243
rect 10243 30187 10299 30243
rect 10385 30187 10441 30243
rect 10527 30187 10583 30243
rect 10669 30187 10725 30243
rect 10811 30187 10867 30243
rect 10953 30187 11009 30243
rect 11095 30187 11151 30243
rect 11237 30187 11293 30243
rect 11379 30187 11435 30243
rect 11521 30187 11577 30243
rect 11663 30187 11719 30243
rect 11805 30187 11861 30243
rect 11947 30187 12003 30243
rect 12089 30187 12145 30243
rect 12231 30187 12287 30243
rect 12373 30187 12429 30243
rect 12515 30187 12571 30243
rect 12657 30187 12713 30243
rect 12799 30187 12855 30243
rect 12941 30187 12997 30243
rect 13083 30187 13139 30243
rect 13225 30187 13281 30243
rect 13367 30187 13423 30243
rect 13509 30187 13565 30243
rect 13651 30187 13707 30243
rect 13793 30187 13849 30243
rect 13935 30187 13991 30243
rect 14077 30187 14133 30243
rect 14219 30187 14275 30243
rect 14361 30187 14417 30243
rect 14503 30187 14559 30243
rect 14645 30187 14701 30243
rect 14787 30187 14843 30243
rect 161 30045 217 30101
rect 303 30045 359 30101
rect 445 30045 501 30101
rect 587 30045 643 30101
rect 729 30045 785 30101
rect 871 30045 927 30101
rect 1013 30045 1069 30101
rect 1155 30045 1211 30101
rect 1297 30045 1353 30101
rect 1439 30045 1495 30101
rect 1581 30045 1637 30101
rect 1723 30045 1779 30101
rect 1865 30045 1921 30101
rect 2007 30045 2063 30101
rect 2149 30045 2205 30101
rect 2291 30045 2347 30101
rect 2433 30045 2489 30101
rect 2575 30045 2631 30101
rect 2717 30045 2773 30101
rect 2859 30045 2915 30101
rect 3001 30045 3057 30101
rect 3143 30045 3199 30101
rect 3285 30045 3341 30101
rect 3427 30045 3483 30101
rect 3569 30045 3625 30101
rect 3711 30045 3767 30101
rect 3853 30045 3909 30101
rect 3995 30045 4051 30101
rect 4137 30045 4193 30101
rect 4279 30045 4335 30101
rect 4421 30045 4477 30101
rect 4563 30045 4619 30101
rect 4705 30045 4761 30101
rect 4847 30045 4903 30101
rect 4989 30045 5045 30101
rect 5131 30045 5187 30101
rect 5273 30045 5329 30101
rect 5415 30045 5471 30101
rect 5557 30045 5613 30101
rect 5699 30045 5755 30101
rect 5841 30045 5897 30101
rect 5983 30045 6039 30101
rect 6125 30045 6181 30101
rect 6267 30045 6323 30101
rect 6409 30045 6465 30101
rect 6551 30045 6607 30101
rect 6693 30045 6749 30101
rect 6835 30045 6891 30101
rect 6977 30045 7033 30101
rect 7119 30045 7175 30101
rect 7261 30045 7317 30101
rect 7403 30045 7459 30101
rect 7545 30045 7601 30101
rect 7687 30045 7743 30101
rect 7829 30045 7885 30101
rect 7971 30045 8027 30101
rect 8113 30045 8169 30101
rect 8255 30045 8311 30101
rect 8397 30045 8453 30101
rect 8539 30045 8595 30101
rect 8681 30045 8737 30101
rect 8823 30045 8879 30101
rect 8965 30045 9021 30101
rect 9107 30045 9163 30101
rect 9249 30045 9305 30101
rect 9391 30045 9447 30101
rect 9533 30045 9589 30101
rect 9675 30045 9731 30101
rect 9817 30045 9873 30101
rect 9959 30045 10015 30101
rect 10101 30045 10157 30101
rect 10243 30045 10299 30101
rect 10385 30045 10441 30101
rect 10527 30045 10583 30101
rect 10669 30045 10725 30101
rect 10811 30045 10867 30101
rect 10953 30045 11009 30101
rect 11095 30045 11151 30101
rect 11237 30045 11293 30101
rect 11379 30045 11435 30101
rect 11521 30045 11577 30101
rect 11663 30045 11719 30101
rect 11805 30045 11861 30101
rect 11947 30045 12003 30101
rect 12089 30045 12145 30101
rect 12231 30045 12287 30101
rect 12373 30045 12429 30101
rect 12515 30045 12571 30101
rect 12657 30045 12713 30101
rect 12799 30045 12855 30101
rect 12941 30045 12997 30101
rect 13083 30045 13139 30101
rect 13225 30045 13281 30101
rect 13367 30045 13423 30101
rect 13509 30045 13565 30101
rect 13651 30045 13707 30101
rect 13793 30045 13849 30101
rect 13935 30045 13991 30101
rect 14077 30045 14133 30101
rect 14219 30045 14275 30101
rect 14361 30045 14417 30101
rect 14503 30045 14559 30101
rect 14645 30045 14701 30101
rect 14787 30045 14843 30101
rect 161 29685 217 29741
rect 303 29685 359 29741
rect 445 29685 501 29741
rect 587 29685 643 29741
rect 729 29685 785 29741
rect 871 29685 927 29741
rect 1013 29685 1069 29741
rect 1155 29685 1211 29741
rect 1297 29685 1353 29741
rect 1439 29685 1495 29741
rect 1581 29685 1637 29741
rect 1723 29685 1779 29741
rect 1865 29685 1921 29741
rect 2007 29685 2063 29741
rect 2149 29685 2205 29741
rect 2291 29685 2347 29741
rect 2433 29685 2489 29741
rect 2575 29685 2631 29741
rect 2717 29685 2773 29741
rect 2859 29685 2915 29741
rect 3001 29685 3057 29741
rect 3143 29685 3199 29741
rect 3285 29685 3341 29741
rect 3427 29685 3483 29741
rect 3569 29685 3625 29741
rect 3711 29685 3767 29741
rect 3853 29685 3909 29741
rect 3995 29685 4051 29741
rect 4137 29685 4193 29741
rect 4279 29685 4335 29741
rect 4421 29685 4477 29741
rect 4563 29685 4619 29741
rect 4705 29685 4761 29741
rect 4847 29685 4903 29741
rect 4989 29685 5045 29741
rect 5131 29685 5187 29741
rect 5273 29685 5329 29741
rect 5415 29685 5471 29741
rect 5557 29685 5613 29741
rect 5699 29685 5755 29741
rect 5841 29685 5897 29741
rect 5983 29685 6039 29741
rect 6125 29685 6181 29741
rect 6267 29685 6323 29741
rect 6409 29685 6465 29741
rect 6551 29685 6607 29741
rect 6693 29685 6749 29741
rect 6835 29685 6891 29741
rect 6977 29685 7033 29741
rect 7119 29685 7175 29741
rect 7261 29685 7317 29741
rect 7403 29685 7459 29741
rect 7545 29685 7601 29741
rect 7687 29685 7743 29741
rect 7829 29685 7885 29741
rect 7971 29685 8027 29741
rect 8113 29685 8169 29741
rect 8255 29685 8311 29741
rect 8397 29685 8453 29741
rect 8539 29685 8595 29741
rect 8681 29685 8737 29741
rect 8823 29685 8879 29741
rect 8965 29685 9021 29741
rect 9107 29685 9163 29741
rect 9249 29685 9305 29741
rect 9391 29685 9447 29741
rect 9533 29685 9589 29741
rect 9675 29685 9731 29741
rect 9817 29685 9873 29741
rect 9959 29685 10015 29741
rect 10101 29685 10157 29741
rect 10243 29685 10299 29741
rect 10385 29685 10441 29741
rect 10527 29685 10583 29741
rect 10669 29685 10725 29741
rect 10811 29685 10867 29741
rect 10953 29685 11009 29741
rect 11095 29685 11151 29741
rect 11237 29685 11293 29741
rect 11379 29685 11435 29741
rect 11521 29685 11577 29741
rect 11663 29685 11719 29741
rect 11805 29685 11861 29741
rect 11947 29685 12003 29741
rect 12089 29685 12145 29741
rect 12231 29685 12287 29741
rect 12373 29685 12429 29741
rect 12515 29685 12571 29741
rect 12657 29685 12713 29741
rect 12799 29685 12855 29741
rect 12941 29685 12997 29741
rect 13083 29685 13139 29741
rect 13225 29685 13281 29741
rect 13367 29685 13423 29741
rect 13509 29685 13565 29741
rect 13651 29685 13707 29741
rect 13793 29685 13849 29741
rect 13935 29685 13991 29741
rect 14077 29685 14133 29741
rect 14219 29685 14275 29741
rect 14361 29685 14417 29741
rect 14503 29685 14559 29741
rect 14645 29685 14701 29741
rect 14787 29685 14843 29741
rect 161 29543 217 29599
rect 303 29543 359 29599
rect 445 29543 501 29599
rect 587 29543 643 29599
rect 729 29543 785 29599
rect 871 29543 927 29599
rect 1013 29543 1069 29599
rect 1155 29543 1211 29599
rect 1297 29543 1353 29599
rect 1439 29543 1495 29599
rect 1581 29543 1637 29599
rect 1723 29543 1779 29599
rect 1865 29543 1921 29599
rect 2007 29543 2063 29599
rect 2149 29543 2205 29599
rect 2291 29543 2347 29599
rect 2433 29543 2489 29599
rect 2575 29543 2631 29599
rect 2717 29543 2773 29599
rect 2859 29543 2915 29599
rect 3001 29543 3057 29599
rect 3143 29543 3199 29599
rect 3285 29543 3341 29599
rect 3427 29543 3483 29599
rect 3569 29543 3625 29599
rect 3711 29543 3767 29599
rect 3853 29543 3909 29599
rect 3995 29543 4051 29599
rect 4137 29543 4193 29599
rect 4279 29543 4335 29599
rect 4421 29543 4477 29599
rect 4563 29543 4619 29599
rect 4705 29543 4761 29599
rect 4847 29543 4903 29599
rect 4989 29543 5045 29599
rect 5131 29543 5187 29599
rect 5273 29543 5329 29599
rect 5415 29543 5471 29599
rect 5557 29543 5613 29599
rect 5699 29543 5755 29599
rect 5841 29543 5897 29599
rect 5983 29543 6039 29599
rect 6125 29543 6181 29599
rect 6267 29543 6323 29599
rect 6409 29543 6465 29599
rect 6551 29543 6607 29599
rect 6693 29543 6749 29599
rect 6835 29543 6891 29599
rect 6977 29543 7033 29599
rect 7119 29543 7175 29599
rect 7261 29543 7317 29599
rect 7403 29543 7459 29599
rect 7545 29543 7601 29599
rect 7687 29543 7743 29599
rect 7829 29543 7885 29599
rect 7971 29543 8027 29599
rect 8113 29543 8169 29599
rect 8255 29543 8311 29599
rect 8397 29543 8453 29599
rect 8539 29543 8595 29599
rect 8681 29543 8737 29599
rect 8823 29543 8879 29599
rect 8965 29543 9021 29599
rect 9107 29543 9163 29599
rect 9249 29543 9305 29599
rect 9391 29543 9447 29599
rect 9533 29543 9589 29599
rect 9675 29543 9731 29599
rect 9817 29543 9873 29599
rect 9959 29543 10015 29599
rect 10101 29543 10157 29599
rect 10243 29543 10299 29599
rect 10385 29543 10441 29599
rect 10527 29543 10583 29599
rect 10669 29543 10725 29599
rect 10811 29543 10867 29599
rect 10953 29543 11009 29599
rect 11095 29543 11151 29599
rect 11237 29543 11293 29599
rect 11379 29543 11435 29599
rect 11521 29543 11577 29599
rect 11663 29543 11719 29599
rect 11805 29543 11861 29599
rect 11947 29543 12003 29599
rect 12089 29543 12145 29599
rect 12231 29543 12287 29599
rect 12373 29543 12429 29599
rect 12515 29543 12571 29599
rect 12657 29543 12713 29599
rect 12799 29543 12855 29599
rect 12941 29543 12997 29599
rect 13083 29543 13139 29599
rect 13225 29543 13281 29599
rect 13367 29543 13423 29599
rect 13509 29543 13565 29599
rect 13651 29543 13707 29599
rect 13793 29543 13849 29599
rect 13935 29543 13991 29599
rect 14077 29543 14133 29599
rect 14219 29543 14275 29599
rect 14361 29543 14417 29599
rect 14503 29543 14559 29599
rect 14645 29543 14701 29599
rect 14787 29543 14843 29599
rect 161 29401 217 29457
rect 303 29401 359 29457
rect 445 29401 501 29457
rect 587 29401 643 29457
rect 729 29401 785 29457
rect 871 29401 927 29457
rect 1013 29401 1069 29457
rect 1155 29401 1211 29457
rect 1297 29401 1353 29457
rect 1439 29401 1495 29457
rect 1581 29401 1637 29457
rect 1723 29401 1779 29457
rect 1865 29401 1921 29457
rect 2007 29401 2063 29457
rect 2149 29401 2205 29457
rect 2291 29401 2347 29457
rect 2433 29401 2489 29457
rect 2575 29401 2631 29457
rect 2717 29401 2773 29457
rect 2859 29401 2915 29457
rect 3001 29401 3057 29457
rect 3143 29401 3199 29457
rect 3285 29401 3341 29457
rect 3427 29401 3483 29457
rect 3569 29401 3625 29457
rect 3711 29401 3767 29457
rect 3853 29401 3909 29457
rect 3995 29401 4051 29457
rect 4137 29401 4193 29457
rect 4279 29401 4335 29457
rect 4421 29401 4477 29457
rect 4563 29401 4619 29457
rect 4705 29401 4761 29457
rect 4847 29401 4903 29457
rect 4989 29401 5045 29457
rect 5131 29401 5187 29457
rect 5273 29401 5329 29457
rect 5415 29401 5471 29457
rect 5557 29401 5613 29457
rect 5699 29401 5755 29457
rect 5841 29401 5897 29457
rect 5983 29401 6039 29457
rect 6125 29401 6181 29457
rect 6267 29401 6323 29457
rect 6409 29401 6465 29457
rect 6551 29401 6607 29457
rect 6693 29401 6749 29457
rect 6835 29401 6891 29457
rect 6977 29401 7033 29457
rect 7119 29401 7175 29457
rect 7261 29401 7317 29457
rect 7403 29401 7459 29457
rect 7545 29401 7601 29457
rect 7687 29401 7743 29457
rect 7829 29401 7885 29457
rect 7971 29401 8027 29457
rect 8113 29401 8169 29457
rect 8255 29401 8311 29457
rect 8397 29401 8453 29457
rect 8539 29401 8595 29457
rect 8681 29401 8737 29457
rect 8823 29401 8879 29457
rect 8965 29401 9021 29457
rect 9107 29401 9163 29457
rect 9249 29401 9305 29457
rect 9391 29401 9447 29457
rect 9533 29401 9589 29457
rect 9675 29401 9731 29457
rect 9817 29401 9873 29457
rect 9959 29401 10015 29457
rect 10101 29401 10157 29457
rect 10243 29401 10299 29457
rect 10385 29401 10441 29457
rect 10527 29401 10583 29457
rect 10669 29401 10725 29457
rect 10811 29401 10867 29457
rect 10953 29401 11009 29457
rect 11095 29401 11151 29457
rect 11237 29401 11293 29457
rect 11379 29401 11435 29457
rect 11521 29401 11577 29457
rect 11663 29401 11719 29457
rect 11805 29401 11861 29457
rect 11947 29401 12003 29457
rect 12089 29401 12145 29457
rect 12231 29401 12287 29457
rect 12373 29401 12429 29457
rect 12515 29401 12571 29457
rect 12657 29401 12713 29457
rect 12799 29401 12855 29457
rect 12941 29401 12997 29457
rect 13083 29401 13139 29457
rect 13225 29401 13281 29457
rect 13367 29401 13423 29457
rect 13509 29401 13565 29457
rect 13651 29401 13707 29457
rect 13793 29401 13849 29457
rect 13935 29401 13991 29457
rect 14077 29401 14133 29457
rect 14219 29401 14275 29457
rect 14361 29401 14417 29457
rect 14503 29401 14559 29457
rect 14645 29401 14701 29457
rect 14787 29401 14843 29457
rect 161 29259 217 29315
rect 303 29259 359 29315
rect 445 29259 501 29315
rect 587 29259 643 29315
rect 729 29259 785 29315
rect 871 29259 927 29315
rect 1013 29259 1069 29315
rect 1155 29259 1211 29315
rect 1297 29259 1353 29315
rect 1439 29259 1495 29315
rect 1581 29259 1637 29315
rect 1723 29259 1779 29315
rect 1865 29259 1921 29315
rect 2007 29259 2063 29315
rect 2149 29259 2205 29315
rect 2291 29259 2347 29315
rect 2433 29259 2489 29315
rect 2575 29259 2631 29315
rect 2717 29259 2773 29315
rect 2859 29259 2915 29315
rect 3001 29259 3057 29315
rect 3143 29259 3199 29315
rect 3285 29259 3341 29315
rect 3427 29259 3483 29315
rect 3569 29259 3625 29315
rect 3711 29259 3767 29315
rect 3853 29259 3909 29315
rect 3995 29259 4051 29315
rect 4137 29259 4193 29315
rect 4279 29259 4335 29315
rect 4421 29259 4477 29315
rect 4563 29259 4619 29315
rect 4705 29259 4761 29315
rect 4847 29259 4903 29315
rect 4989 29259 5045 29315
rect 5131 29259 5187 29315
rect 5273 29259 5329 29315
rect 5415 29259 5471 29315
rect 5557 29259 5613 29315
rect 5699 29259 5755 29315
rect 5841 29259 5897 29315
rect 5983 29259 6039 29315
rect 6125 29259 6181 29315
rect 6267 29259 6323 29315
rect 6409 29259 6465 29315
rect 6551 29259 6607 29315
rect 6693 29259 6749 29315
rect 6835 29259 6891 29315
rect 6977 29259 7033 29315
rect 7119 29259 7175 29315
rect 7261 29259 7317 29315
rect 7403 29259 7459 29315
rect 7545 29259 7601 29315
rect 7687 29259 7743 29315
rect 7829 29259 7885 29315
rect 7971 29259 8027 29315
rect 8113 29259 8169 29315
rect 8255 29259 8311 29315
rect 8397 29259 8453 29315
rect 8539 29259 8595 29315
rect 8681 29259 8737 29315
rect 8823 29259 8879 29315
rect 8965 29259 9021 29315
rect 9107 29259 9163 29315
rect 9249 29259 9305 29315
rect 9391 29259 9447 29315
rect 9533 29259 9589 29315
rect 9675 29259 9731 29315
rect 9817 29259 9873 29315
rect 9959 29259 10015 29315
rect 10101 29259 10157 29315
rect 10243 29259 10299 29315
rect 10385 29259 10441 29315
rect 10527 29259 10583 29315
rect 10669 29259 10725 29315
rect 10811 29259 10867 29315
rect 10953 29259 11009 29315
rect 11095 29259 11151 29315
rect 11237 29259 11293 29315
rect 11379 29259 11435 29315
rect 11521 29259 11577 29315
rect 11663 29259 11719 29315
rect 11805 29259 11861 29315
rect 11947 29259 12003 29315
rect 12089 29259 12145 29315
rect 12231 29259 12287 29315
rect 12373 29259 12429 29315
rect 12515 29259 12571 29315
rect 12657 29259 12713 29315
rect 12799 29259 12855 29315
rect 12941 29259 12997 29315
rect 13083 29259 13139 29315
rect 13225 29259 13281 29315
rect 13367 29259 13423 29315
rect 13509 29259 13565 29315
rect 13651 29259 13707 29315
rect 13793 29259 13849 29315
rect 13935 29259 13991 29315
rect 14077 29259 14133 29315
rect 14219 29259 14275 29315
rect 14361 29259 14417 29315
rect 14503 29259 14559 29315
rect 14645 29259 14701 29315
rect 14787 29259 14843 29315
rect 161 29117 217 29173
rect 303 29117 359 29173
rect 445 29117 501 29173
rect 587 29117 643 29173
rect 729 29117 785 29173
rect 871 29117 927 29173
rect 1013 29117 1069 29173
rect 1155 29117 1211 29173
rect 1297 29117 1353 29173
rect 1439 29117 1495 29173
rect 1581 29117 1637 29173
rect 1723 29117 1779 29173
rect 1865 29117 1921 29173
rect 2007 29117 2063 29173
rect 2149 29117 2205 29173
rect 2291 29117 2347 29173
rect 2433 29117 2489 29173
rect 2575 29117 2631 29173
rect 2717 29117 2773 29173
rect 2859 29117 2915 29173
rect 3001 29117 3057 29173
rect 3143 29117 3199 29173
rect 3285 29117 3341 29173
rect 3427 29117 3483 29173
rect 3569 29117 3625 29173
rect 3711 29117 3767 29173
rect 3853 29117 3909 29173
rect 3995 29117 4051 29173
rect 4137 29117 4193 29173
rect 4279 29117 4335 29173
rect 4421 29117 4477 29173
rect 4563 29117 4619 29173
rect 4705 29117 4761 29173
rect 4847 29117 4903 29173
rect 4989 29117 5045 29173
rect 5131 29117 5187 29173
rect 5273 29117 5329 29173
rect 5415 29117 5471 29173
rect 5557 29117 5613 29173
rect 5699 29117 5755 29173
rect 5841 29117 5897 29173
rect 5983 29117 6039 29173
rect 6125 29117 6181 29173
rect 6267 29117 6323 29173
rect 6409 29117 6465 29173
rect 6551 29117 6607 29173
rect 6693 29117 6749 29173
rect 6835 29117 6891 29173
rect 6977 29117 7033 29173
rect 7119 29117 7175 29173
rect 7261 29117 7317 29173
rect 7403 29117 7459 29173
rect 7545 29117 7601 29173
rect 7687 29117 7743 29173
rect 7829 29117 7885 29173
rect 7971 29117 8027 29173
rect 8113 29117 8169 29173
rect 8255 29117 8311 29173
rect 8397 29117 8453 29173
rect 8539 29117 8595 29173
rect 8681 29117 8737 29173
rect 8823 29117 8879 29173
rect 8965 29117 9021 29173
rect 9107 29117 9163 29173
rect 9249 29117 9305 29173
rect 9391 29117 9447 29173
rect 9533 29117 9589 29173
rect 9675 29117 9731 29173
rect 9817 29117 9873 29173
rect 9959 29117 10015 29173
rect 10101 29117 10157 29173
rect 10243 29117 10299 29173
rect 10385 29117 10441 29173
rect 10527 29117 10583 29173
rect 10669 29117 10725 29173
rect 10811 29117 10867 29173
rect 10953 29117 11009 29173
rect 11095 29117 11151 29173
rect 11237 29117 11293 29173
rect 11379 29117 11435 29173
rect 11521 29117 11577 29173
rect 11663 29117 11719 29173
rect 11805 29117 11861 29173
rect 11947 29117 12003 29173
rect 12089 29117 12145 29173
rect 12231 29117 12287 29173
rect 12373 29117 12429 29173
rect 12515 29117 12571 29173
rect 12657 29117 12713 29173
rect 12799 29117 12855 29173
rect 12941 29117 12997 29173
rect 13083 29117 13139 29173
rect 13225 29117 13281 29173
rect 13367 29117 13423 29173
rect 13509 29117 13565 29173
rect 13651 29117 13707 29173
rect 13793 29117 13849 29173
rect 13935 29117 13991 29173
rect 14077 29117 14133 29173
rect 14219 29117 14275 29173
rect 14361 29117 14417 29173
rect 14503 29117 14559 29173
rect 14645 29117 14701 29173
rect 14787 29117 14843 29173
rect 161 28975 217 29031
rect 303 28975 359 29031
rect 445 28975 501 29031
rect 587 28975 643 29031
rect 729 28975 785 29031
rect 871 28975 927 29031
rect 1013 28975 1069 29031
rect 1155 28975 1211 29031
rect 1297 28975 1353 29031
rect 1439 28975 1495 29031
rect 1581 28975 1637 29031
rect 1723 28975 1779 29031
rect 1865 28975 1921 29031
rect 2007 28975 2063 29031
rect 2149 28975 2205 29031
rect 2291 28975 2347 29031
rect 2433 28975 2489 29031
rect 2575 28975 2631 29031
rect 2717 28975 2773 29031
rect 2859 28975 2915 29031
rect 3001 28975 3057 29031
rect 3143 28975 3199 29031
rect 3285 28975 3341 29031
rect 3427 28975 3483 29031
rect 3569 28975 3625 29031
rect 3711 28975 3767 29031
rect 3853 28975 3909 29031
rect 3995 28975 4051 29031
rect 4137 28975 4193 29031
rect 4279 28975 4335 29031
rect 4421 28975 4477 29031
rect 4563 28975 4619 29031
rect 4705 28975 4761 29031
rect 4847 28975 4903 29031
rect 4989 28975 5045 29031
rect 5131 28975 5187 29031
rect 5273 28975 5329 29031
rect 5415 28975 5471 29031
rect 5557 28975 5613 29031
rect 5699 28975 5755 29031
rect 5841 28975 5897 29031
rect 5983 28975 6039 29031
rect 6125 28975 6181 29031
rect 6267 28975 6323 29031
rect 6409 28975 6465 29031
rect 6551 28975 6607 29031
rect 6693 28975 6749 29031
rect 6835 28975 6891 29031
rect 6977 28975 7033 29031
rect 7119 28975 7175 29031
rect 7261 28975 7317 29031
rect 7403 28975 7459 29031
rect 7545 28975 7601 29031
rect 7687 28975 7743 29031
rect 7829 28975 7885 29031
rect 7971 28975 8027 29031
rect 8113 28975 8169 29031
rect 8255 28975 8311 29031
rect 8397 28975 8453 29031
rect 8539 28975 8595 29031
rect 8681 28975 8737 29031
rect 8823 28975 8879 29031
rect 8965 28975 9021 29031
rect 9107 28975 9163 29031
rect 9249 28975 9305 29031
rect 9391 28975 9447 29031
rect 9533 28975 9589 29031
rect 9675 28975 9731 29031
rect 9817 28975 9873 29031
rect 9959 28975 10015 29031
rect 10101 28975 10157 29031
rect 10243 28975 10299 29031
rect 10385 28975 10441 29031
rect 10527 28975 10583 29031
rect 10669 28975 10725 29031
rect 10811 28975 10867 29031
rect 10953 28975 11009 29031
rect 11095 28975 11151 29031
rect 11237 28975 11293 29031
rect 11379 28975 11435 29031
rect 11521 28975 11577 29031
rect 11663 28975 11719 29031
rect 11805 28975 11861 29031
rect 11947 28975 12003 29031
rect 12089 28975 12145 29031
rect 12231 28975 12287 29031
rect 12373 28975 12429 29031
rect 12515 28975 12571 29031
rect 12657 28975 12713 29031
rect 12799 28975 12855 29031
rect 12941 28975 12997 29031
rect 13083 28975 13139 29031
rect 13225 28975 13281 29031
rect 13367 28975 13423 29031
rect 13509 28975 13565 29031
rect 13651 28975 13707 29031
rect 13793 28975 13849 29031
rect 13935 28975 13991 29031
rect 14077 28975 14133 29031
rect 14219 28975 14275 29031
rect 14361 28975 14417 29031
rect 14503 28975 14559 29031
rect 14645 28975 14701 29031
rect 14787 28975 14843 29031
rect 161 28833 217 28889
rect 303 28833 359 28889
rect 445 28833 501 28889
rect 587 28833 643 28889
rect 729 28833 785 28889
rect 871 28833 927 28889
rect 1013 28833 1069 28889
rect 1155 28833 1211 28889
rect 1297 28833 1353 28889
rect 1439 28833 1495 28889
rect 1581 28833 1637 28889
rect 1723 28833 1779 28889
rect 1865 28833 1921 28889
rect 2007 28833 2063 28889
rect 2149 28833 2205 28889
rect 2291 28833 2347 28889
rect 2433 28833 2489 28889
rect 2575 28833 2631 28889
rect 2717 28833 2773 28889
rect 2859 28833 2915 28889
rect 3001 28833 3057 28889
rect 3143 28833 3199 28889
rect 3285 28833 3341 28889
rect 3427 28833 3483 28889
rect 3569 28833 3625 28889
rect 3711 28833 3767 28889
rect 3853 28833 3909 28889
rect 3995 28833 4051 28889
rect 4137 28833 4193 28889
rect 4279 28833 4335 28889
rect 4421 28833 4477 28889
rect 4563 28833 4619 28889
rect 4705 28833 4761 28889
rect 4847 28833 4903 28889
rect 4989 28833 5045 28889
rect 5131 28833 5187 28889
rect 5273 28833 5329 28889
rect 5415 28833 5471 28889
rect 5557 28833 5613 28889
rect 5699 28833 5755 28889
rect 5841 28833 5897 28889
rect 5983 28833 6039 28889
rect 6125 28833 6181 28889
rect 6267 28833 6323 28889
rect 6409 28833 6465 28889
rect 6551 28833 6607 28889
rect 6693 28833 6749 28889
rect 6835 28833 6891 28889
rect 6977 28833 7033 28889
rect 7119 28833 7175 28889
rect 7261 28833 7317 28889
rect 7403 28833 7459 28889
rect 7545 28833 7601 28889
rect 7687 28833 7743 28889
rect 7829 28833 7885 28889
rect 7971 28833 8027 28889
rect 8113 28833 8169 28889
rect 8255 28833 8311 28889
rect 8397 28833 8453 28889
rect 8539 28833 8595 28889
rect 8681 28833 8737 28889
rect 8823 28833 8879 28889
rect 8965 28833 9021 28889
rect 9107 28833 9163 28889
rect 9249 28833 9305 28889
rect 9391 28833 9447 28889
rect 9533 28833 9589 28889
rect 9675 28833 9731 28889
rect 9817 28833 9873 28889
rect 9959 28833 10015 28889
rect 10101 28833 10157 28889
rect 10243 28833 10299 28889
rect 10385 28833 10441 28889
rect 10527 28833 10583 28889
rect 10669 28833 10725 28889
rect 10811 28833 10867 28889
rect 10953 28833 11009 28889
rect 11095 28833 11151 28889
rect 11237 28833 11293 28889
rect 11379 28833 11435 28889
rect 11521 28833 11577 28889
rect 11663 28833 11719 28889
rect 11805 28833 11861 28889
rect 11947 28833 12003 28889
rect 12089 28833 12145 28889
rect 12231 28833 12287 28889
rect 12373 28833 12429 28889
rect 12515 28833 12571 28889
rect 12657 28833 12713 28889
rect 12799 28833 12855 28889
rect 12941 28833 12997 28889
rect 13083 28833 13139 28889
rect 13225 28833 13281 28889
rect 13367 28833 13423 28889
rect 13509 28833 13565 28889
rect 13651 28833 13707 28889
rect 13793 28833 13849 28889
rect 13935 28833 13991 28889
rect 14077 28833 14133 28889
rect 14219 28833 14275 28889
rect 14361 28833 14417 28889
rect 14503 28833 14559 28889
rect 14645 28833 14701 28889
rect 14787 28833 14843 28889
rect 161 28691 217 28747
rect 303 28691 359 28747
rect 445 28691 501 28747
rect 587 28691 643 28747
rect 729 28691 785 28747
rect 871 28691 927 28747
rect 1013 28691 1069 28747
rect 1155 28691 1211 28747
rect 1297 28691 1353 28747
rect 1439 28691 1495 28747
rect 1581 28691 1637 28747
rect 1723 28691 1779 28747
rect 1865 28691 1921 28747
rect 2007 28691 2063 28747
rect 2149 28691 2205 28747
rect 2291 28691 2347 28747
rect 2433 28691 2489 28747
rect 2575 28691 2631 28747
rect 2717 28691 2773 28747
rect 2859 28691 2915 28747
rect 3001 28691 3057 28747
rect 3143 28691 3199 28747
rect 3285 28691 3341 28747
rect 3427 28691 3483 28747
rect 3569 28691 3625 28747
rect 3711 28691 3767 28747
rect 3853 28691 3909 28747
rect 3995 28691 4051 28747
rect 4137 28691 4193 28747
rect 4279 28691 4335 28747
rect 4421 28691 4477 28747
rect 4563 28691 4619 28747
rect 4705 28691 4761 28747
rect 4847 28691 4903 28747
rect 4989 28691 5045 28747
rect 5131 28691 5187 28747
rect 5273 28691 5329 28747
rect 5415 28691 5471 28747
rect 5557 28691 5613 28747
rect 5699 28691 5755 28747
rect 5841 28691 5897 28747
rect 5983 28691 6039 28747
rect 6125 28691 6181 28747
rect 6267 28691 6323 28747
rect 6409 28691 6465 28747
rect 6551 28691 6607 28747
rect 6693 28691 6749 28747
rect 6835 28691 6891 28747
rect 6977 28691 7033 28747
rect 7119 28691 7175 28747
rect 7261 28691 7317 28747
rect 7403 28691 7459 28747
rect 7545 28691 7601 28747
rect 7687 28691 7743 28747
rect 7829 28691 7885 28747
rect 7971 28691 8027 28747
rect 8113 28691 8169 28747
rect 8255 28691 8311 28747
rect 8397 28691 8453 28747
rect 8539 28691 8595 28747
rect 8681 28691 8737 28747
rect 8823 28691 8879 28747
rect 8965 28691 9021 28747
rect 9107 28691 9163 28747
rect 9249 28691 9305 28747
rect 9391 28691 9447 28747
rect 9533 28691 9589 28747
rect 9675 28691 9731 28747
rect 9817 28691 9873 28747
rect 9959 28691 10015 28747
rect 10101 28691 10157 28747
rect 10243 28691 10299 28747
rect 10385 28691 10441 28747
rect 10527 28691 10583 28747
rect 10669 28691 10725 28747
rect 10811 28691 10867 28747
rect 10953 28691 11009 28747
rect 11095 28691 11151 28747
rect 11237 28691 11293 28747
rect 11379 28691 11435 28747
rect 11521 28691 11577 28747
rect 11663 28691 11719 28747
rect 11805 28691 11861 28747
rect 11947 28691 12003 28747
rect 12089 28691 12145 28747
rect 12231 28691 12287 28747
rect 12373 28691 12429 28747
rect 12515 28691 12571 28747
rect 12657 28691 12713 28747
rect 12799 28691 12855 28747
rect 12941 28691 12997 28747
rect 13083 28691 13139 28747
rect 13225 28691 13281 28747
rect 13367 28691 13423 28747
rect 13509 28691 13565 28747
rect 13651 28691 13707 28747
rect 13793 28691 13849 28747
rect 13935 28691 13991 28747
rect 14077 28691 14133 28747
rect 14219 28691 14275 28747
rect 14361 28691 14417 28747
rect 14503 28691 14559 28747
rect 14645 28691 14701 28747
rect 14787 28691 14843 28747
rect 161 28549 217 28605
rect 303 28549 359 28605
rect 445 28549 501 28605
rect 587 28549 643 28605
rect 729 28549 785 28605
rect 871 28549 927 28605
rect 1013 28549 1069 28605
rect 1155 28549 1211 28605
rect 1297 28549 1353 28605
rect 1439 28549 1495 28605
rect 1581 28549 1637 28605
rect 1723 28549 1779 28605
rect 1865 28549 1921 28605
rect 2007 28549 2063 28605
rect 2149 28549 2205 28605
rect 2291 28549 2347 28605
rect 2433 28549 2489 28605
rect 2575 28549 2631 28605
rect 2717 28549 2773 28605
rect 2859 28549 2915 28605
rect 3001 28549 3057 28605
rect 3143 28549 3199 28605
rect 3285 28549 3341 28605
rect 3427 28549 3483 28605
rect 3569 28549 3625 28605
rect 3711 28549 3767 28605
rect 3853 28549 3909 28605
rect 3995 28549 4051 28605
rect 4137 28549 4193 28605
rect 4279 28549 4335 28605
rect 4421 28549 4477 28605
rect 4563 28549 4619 28605
rect 4705 28549 4761 28605
rect 4847 28549 4903 28605
rect 4989 28549 5045 28605
rect 5131 28549 5187 28605
rect 5273 28549 5329 28605
rect 5415 28549 5471 28605
rect 5557 28549 5613 28605
rect 5699 28549 5755 28605
rect 5841 28549 5897 28605
rect 5983 28549 6039 28605
rect 6125 28549 6181 28605
rect 6267 28549 6323 28605
rect 6409 28549 6465 28605
rect 6551 28549 6607 28605
rect 6693 28549 6749 28605
rect 6835 28549 6891 28605
rect 6977 28549 7033 28605
rect 7119 28549 7175 28605
rect 7261 28549 7317 28605
rect 7403 28549 7459 28605
rect 7545 28549 7601 28605
rect 7687 28549 7743 28605
rect 7829 28549 7885 28605
rect 7971 28549 8027 28605
rect 8113 28549 8169 28605
rect 8255 28549 8311 28605
rect 8397 28549 8453 28605
rect 8539 28549 8595 28605
rect 8681 28549 8737 28605
rect 8823 28549 8879 28605
rect 8965 28549 9021 28605
rect 9107 28549 9163 28605
rect 9249 28549 9305 28605
rect 9391 28549 9447 28605
rect 9533 28549 9589 28605
rect 9675 28549 9731 28605
rect 9817 28549 9873 28605
rect 9959 28549 10015 28605
rect 10101 28549 10157 28605
rect 10243 28549 10299 28605
rect 10385 28549 10441 28605
rect 10527 28549 10583 28605
rect 10669 28549 10725 28605
rect 10811 28549 10867 28605
rect 10953 28549 11009 28605
rect 11095 28549 11151 28605
rect 11237 28549 11293 28605
rect 11379 28549 11435 28605
rect 11521 28549 11577 28605
rect 11663 28549 11719 28605
rect 11805 28549 11861 28605
rect 11947 28549 12003 28605
rect 12089 28549 12145 28605
rect 12231 28549 12287 28605
rect 12373 28549 12429 28605
rect 12515 28549 12571 28605
rect 12657 28549 12713 28605
rect 12799 28549 12855 28605
rect 12941 28549 12997 28605
rect 13083 28549 13139 28605
rect 13225 28549 13281 28605
rect 13367 28549 13423 28605
rect 13509 28549 13565 28605
rect 13651 28549 13707 28605
rect 13793 28549 13849 28605
rect 13935 28549 13991 28605
rect 14077 28549 14133 28605
rect 14219 28549 14275 28605
rect 14361 28549 14417 28605
rect 14503 28549 14559 28605
rect 14645 28549 14701 28605
rect 14787 28549 14843 28605
rect 161 28407 217 28463
rect 303 28407 359 28463
rect 445 28407 501 28463
rect 587 28407 643 28463
rect 729 28407 785 28463
rect 871 28407 927 28463
rect 1013 28407 1069 28463
rect 1155 28407 1211 28463
rect 1297 28407 1353 28463
rect 1439 28407 1495 28463
rect 1581 28407 1637 28463
rect 1723 28407 1779 28463
rect 1865 28407 1921 28463
rect 2007 28407 2063 28463
rect 2149 28407 2205 28463
rect 2291 28407 2347 28463
rect 2433 28407 2489 28463
rect 2575 28407 2631 28463
rect 2717 28407 2773 28463
rect 2859 28407 2915 28463
rect 3001 28407 3057 28463
rect 3143 28407 3199 28463
rect 3285 28407 3341 28463
rect 3427 28407 3483 28463
rect 3569 28407 3625 28463
rect 3711 28407 3767 28463
rect 3853 28407 3909 28463
rect 3995 28407 4051 28463
rect 4137 28407 4193 28463
rect 4279 28407 4335 28463
rect 4421 28407 4477 28463
rect 4563 28407 4619 28463
rect 4705 28407 4761 28463
rect 4847 28407 4903 28463
rect 4989 28407 5045 28463
rect 5131 28407 5187 28463
rect 5273 28407 5329 28463
rect 5415 28407 5471 28463
rect 5557 28407 5613 28463
rect 5699 28407 5755 28463
rect 5841 28407 5897 28463
rect 5983 28407 6039 28463
rect 6125 28407 6181 28463
rect 6267 28407 6323 28463
rect 6409 28407 6465 28463
rect 6551 28407 6607 28463
rect 6693 28407 6749 28463
rect 6835 28407 6891 28463
rect 6977 28407 7033 28463
rect 7119 28407 7175 28463
rect 7261 28407 7317 28463
rect 7403 28407 7459 28463
rect 7545 28407 7601 28463
rect 7687 28407 7743 28463
rect 7829 28407 7885 28463
rect 7971 28407 8027 28463
rect 8113 28407 8169 28463
rect 8255 28407 8311 28463
rect 8397 28407 8453 28463
rect 8539 28407 8595 28463
rect 8681 28407 8737 28463
rect 8823 28407 8879 28463
rect 8965 28407 9021 28463
rect 9107 28407 9163 28463
rect 9249 28407 9305 28463
rect 9391 28407 9447 28463
rect 9533 28407 9589 28463
rect 9675 28407 9731 28463
rect 9817 28407 9873 28463
rect 9959 28407 10015 28463
rect 10101 28407 10157 28463
rect 10243 28407 10299 28463
rect 10385 28407 10441 28463
rect 10527 28407 10583 28463
rect 10669 28407 10725 28463
rect 10811 28407 10867 28463
rect 10953 28407 11009 28463
rect 11095 28407 11151 28463
rect 11237 28407 11293 28463
rect 11379 28407 11435 28463
rect 11521 28407 11577 28463
rect 11663 28407 11719 28463
rect 11805 28407 11861 28463
rect 11947 28407 12003 28463
rect 12089 28407 12145 28463
rect 12231 28407 12287 28463
rect 12373 28407 12429 28463
rect 12515 28407 12571 28463
rect 12657 28407 12713 28463
rect 12799 28407 12855 28463
rect 12941 28407 12997 28463
rect 13083 28407 13139 28463
rect 13225 28407 13281 28463
rect 13367 28407 13423 28463
rect 13509 28407 13565 28463
rect 13651 28407 13707 28463
rect 13793 28407 13849 28463
rect 13935 28407 13991 28463
rect 14077 28407 14133 28463
rect 14219 28407 14275 28463
rect 14361 28407 14417 28463
rect 14503 28407 14559 28463
rect 14645 28407 14701 28463
rect 14787 28407 14843 28463
rect 161 28265 217 28321
rect 303 28265 359 28321
rect 445 28265 501 28321
rect 587 28265 643 28321
rect 729 28265 785 28321
rect 871 28265 927 28321
rect 1013 28265 1069 28321
rect 1155 28265 1211 28321
rect 1297 28265 1353 28321
rect 1439 28265 1495 28321
rect 1581 28265 1637 28321
rect 1723 28265 1779 28321
rect 1865 28265 1921 28321
rect 2007 28265 2063 28321
rect 2149 28265 2205 28321
rect 2291 28265 2347 28321
rect 2433 28265 2489 28321
rect 2575 28265 2631 28321
rect 2717 28265 2773 28321
rect 2859 28265 2915 28321
rect 3001 28265 3057 28321
rect 3143 28265 3199 28321
rect 3285 28265 3341 28321
rect 3427 28265 3483 28321
rect 3569 28265 3625 28321
rect 3711 28265 3767 28321
rect 3853 28265 3909 28321
rect 3995 28265 4051 28321
rect 4137 28265 4193 28321
rect 4279 28265 4335 28321
rect 4421 28265 4477 28321
rect 4563 28265 4619 28321
rect 4705 28265 4761 28321
rect 4847 28265 4903 28321
rect 4989 28265 5045 28321
rect 5131 28265 5187 28321
rect 5273 28265 5329 28321
rect 5415 28265 5471 28321
rect 5557 28265 5613 28321
rect 5699 28265 5755 28321
rect 5841 28265 5897 28321
rect 5983 28265 6039 28321
rect 6125 28265 6181 28321
rect 6267 28265 6323 28321
rect 6409 28265 6465 28321
rect 6551 28265 6607 28321
rect 6693 28265 6749 28321
rect 6835 28265 6891 28321
rect 6977 28265 7033 28321
rect 7119 28265 7175 28321
rect 7261 28265 7317 28321
rect 7403 28265 7459 28321
rect 7545 28265 7601 28321
rect 7687 28265 7743 28321
rect 7829 28265 7885 28321
rect 7971 28265 8027 28321
rect 8113 28265 8169 28321
rect 8255 28265 8311 28321
rect 8397 28265 8453 28321
rect 8539 28265 8595 28321
rect 8681 28265 8737 28321
rect 8823 28265 8879 28321
rect 8965 28265 9021 28321
rect 9107 28265 9163 28321
rect 9249 28265 9305 28321
rect 9391 28265 9447 28321
rect 9533 28265 9589 28321
rect 9675 28265 9731 28321
rect 9817 28265 9873 28321
rect 9959 28265 10015 28321
rect 10101 28265 10157 28321
rect 10243 28265 10299 28321
rect 10385 28265 10441 28321
rect 10527 28265 10583 28321
rect 10669 28265 10725 28321
rect 10811 28265 10867 28321
rect 10953 28265 11009 28321
rect 11095 28265 11151 28321
rect 11237 28265 11293 28321
rect 11379 28265 11435 28321
rect 11521 28265 11577 28321
rect 11663 28265 11719 28321
rect 11805 28265 11861 28321
rect 11947 28265 12003 28321
rect 12089 28265 12145 28321
rect 12231 28265 12287 28321
rect 12373 28265 12429 28321
rect 12515 28265 12571 28321
rect 12657 28265 12713 28321
rect 12799 28265 12855 28321
rect 12941 28265 12997 28321
rect 13083 28265 13139 28321
rect 13225 28265 13281 28321
rect 13367 28265 13423 28321
rect 13509 28265 13565 28321
rect 13651 28265 13707 28321
rect 13793 28265 13849 28321
rect 13935 28265 13991 28321
rect 14077 28265 14133 28321
rect 14219 28265 14275 28321
rect 14361 28265 14417 28321
rect 14503 28265 14559 28321
rect 14645 28265 14701 28321
rect 14787 28265 14843 28321
rect 161 28123 217 28179
rect 303 28123 359 28179
rect 445 28123 501 28179
rect 587 28123 643 28179
rect 729 28123 785 28179
rect 871 28123 927 28179
rect 1013 28123 1069 28179
rect 1155 28123 1211 28179
rect 1297 28123 1353 28179
rect 1439 28123 1495 28179
rect 1581 28123 1637 28179
rect 1723 28123 1779 28179
rect 1865 28123 1921 28179
rect 2007 28123 2063 28179
rect 2149 28123 2205 28179
rect 2291 28123 2347 28179
rect 2433 28123 2489 28179
rect 2575 28123 2631 28179
rect 2717 28123 2773 28179
rect 2859 28123 2915 28179
rect 3001 28123 3057 28179
rect 3143 28123 3199 28179
rect 3285 28123 3341 28179
rect 3427 28123 3483 28179
rect 3569 28123 3625 28179
rect 3711 28123 3767 28179
rect 3853 28123 3909 28179
rect 3995 28123 4051 28179
rect 4137 28123 4193 28179
rect 4279 28123 4335 28179
rect 4421 28123 4477 28179
rect 4563 28123 4619 28179
rect 4705 28123 4761 28179
rect 4847 28123 4903 28179
rect 4989 28123 5045 28179
rect 5131 28123 5187 28179
rect 5273 28123 5329 28179
rect 5415 28123 5471 28179
rect 5557 28123 5613 28179
rect 5699 28123 5755 28179
rect 5841 28123 5897 28179
rect 5983 28123 6039 28179
rect 6125 28123 6181 28179
rect 6267 28123 6323 28179
rect 6409 28123 6465 28179
rect 6551 28123 6607 28179
rect 6693 28123 6749 28179
rect 6835 28123 6891 28179
rect 6977 28123 7033 28179
rect 7119 28123 7175 28179
rect 7261 28123 7317 28179
rect 7403 28123 7459 28179
rect 7545 28123 7601 28179
rect 7687 28123 7743 28179
rect 7829 28123 7885 28179
rect 7971 28123 8027 28179
rect 8113 28123 8169 28179
rect 8255 28123 8311 28179
rect 8397 28123 8453 28179
rect 8539 28123 8595 28179
rect 8681 28123 8737 28179
rect 8823 28123 8879 28179
rect 8965 28123 9021 28179
rect 9107 28123 9163 28179
rect 9249 28123 9305 28179
rect 9391 28123 9447 28179
rect 9533 28123 9589 28179
rect 9675 28123 9731 28179
rect 9817 28123 9873 28179
rect 9959 28123 10015 28179
rect 10101 28123 10157 28179
rect 10243 28123 10299 28179
rect 10385 28123 10441 28179
rect 10527 28123 10583 28179
rect 10669 28123 10725 28179
rect 10811 28123 10867 28179
rect 10953 28123 11009 28179
rect 11095 28123 11151 28179
rect 11237 28123 11293 28179
rect 11379 28123 11435 28179
rect 11521 28123 11577 28179
rect 11663 28123 11719 28179
rect 11805 28123 11861 28179
rect 11947 28123 12003 28179
rect 12089 28123 12145 28179
rect 12231 28123 12287 28179
rect 12373 28123 12429 28179
rect 12515 28123 12571 28179
rect 12657 28123 12713 28179
rect 12799 28123 12855 28179
rect 12941 28123 12997 28179
rect 13083 28123 13139 28179
rect 13225 28123 13281 28179
rect 13367 28123 13423 28179
rect 13509 28123 13565 28179
rect 13651 28123 13707 28179
rect 13793 28123 13849 28179
rect 13935 28123 13991 28179
rect 14077 28123 14133 28179
rect 14219 28123 14275 28179
rect 14361 28123 14417 28179
rect 14503 28123 14559 28179
rect 14645 28123 14701 28179
rect 14787 28123 14843 28179
rect 161 27981 217 28037
rect 303 27981 359 28037
rect 445 27981 501 28037
rect 587 27981 643 28037
rect 729 27981 785 28037
rect 871 27981 927 28037
rect 1013 27981 1069 28037
rect 1155 27981 1211 28037
rect 1297 27981 1353 28037
rect 1439 27981 1495 28037
rect 1581 27981 1637 28037
rect 1723 27981 1779 28037
rect 1865 27981 1921 28037
rect 2007 27981 2063 28037
rect 2149 27981 2205 28037
rect 2291 27981 2347 28037
rect 2433 27981 2489 28037
rect 2575 27981 2631 28037
rect 2717 27981 2773 28037
rect 2859 27981 2915 28037
rect 3001 27981 3057 28037
rect 3143 27981 3199 28037
rect 3285 27981 3341 28037
rect 3427 27981 3483 28037
rect 3569 27981 3625 28037
rect 3711 27981 3767 28037
rect 3853 27981 3909 28037
rect 3995 27981 4051 28037
rect 4137 27981 4193 28037
rect 4279 27981 4335 28037
rect 4421 27981 4477 28037
rect 4563 27981 4619 28037
rect 4705 27981 4761 28037
rect 4847 27981 4903 28037
rect 4989 27981 5045 28037
rect 5131 27981 5187 28037
rect 5273 27981 5329 28037
rect 5415 27981 5471 28037
rect 5557 27981 5613 28037
rect 5699 27981 5755 28037
rect 5841 27981 5897 28037
rect 5983 27981 6039 28037
rect 6125 27981 6181 28037
rect 6267 27981 6323 28037
rect 6409 27981 6465 28037
rect 6551 27981 6607 28037
rect 6693 27981 6749 28037
rect 6835 27981 6891 28037
rect 6977 27981 7033 28037
rect 7119 27981 7175 28037
rect 7261 27981 7317 28037
rect 7403 27981 7459 28037
rect 7545 27981 7601 28037
rect 7687 27981 7743 28037
rect 7829 27981 7885 28037
rect 7971 27981 8027 28037
rect 8113 27981 8169 28037
rect 8255 27981 8311 28037
rect 8397 27981 8453 28037
rect 8539 27981 8595 28037
rect 8681 27981 8737 28037
rect 8823 27981 8879 28037
rect 8965 27981 9021 28037
rect 9107 27981 9163 28037
rect 9249 27981 9305 28037
rect 9391 27981 9447 28037
rect 9533 27981 9589 28037
rect 9675 27981 9731 28037
rect 9817 27981 9873 28037
rect 9959 27981 10015 28037
rect 10101 27981 10157 28037
rect 10243 27981 10299 28037
rect 10385 27981 10441 28037
rect 10527 27981 10583 28037
rect 10669 27981 10725 28037
rect 10811 27981 10867 28037
rect 10953 27981 11009 28037
rect 11095 27981 11151 28037
rect 11237 27981 11293 28037
rect 11379 27981 11435 28037
rect 11521 27981 11577 28037
rect 11663 27981 11719 28037
rect 11805 27981 11861 28037
rect 11947 27981 12003 28037
rect 12089 27981 12145 28037
rect 12231 27981 12287 28037
rect 12373 27981 12429 28037
rect 12515 27981 12571 28037
rect 12657 27981 12713 28037
rect 12799 27981 12855 28037
rect 12941 27981 12997 28037
rect 13083 27981 13139 28037
rect 13225 27981 13281 28037
rect 13367 27981 13423 28037
rect 13509 27981 13565 28037
rect 13651 27981 13707 28037
rect 13793 27981 13849 28037
rect 13935 27981 13991 28037
rect 14077 27981 14133 28037
rect 14219 27981 14275 28037
rect 14361 27981 14417 28037
rect 14503 27981 14559 28037
rect 14645 27981 14701 28037
rect 14787 27981 14843 28037
rect 161 27839 217 27895
rect 303 27839 359 27895
rect 445 27839 501 27895
rect 587 27839 643 27895
rect 729 27839 785 27895
rect 871 27839 927 27895
rect 1013 27839 1069 27895
rect 1155 27839 1211 27895
rect 1297 27839 1353 27895
rect 1439 27839 1495 27895
rect 1581 27839 1637 27895
rect 1723 27839 1779 27895
rect 1865 27839 1921 27895
rect 2007 27839 2063 27895
rect 2149 27839 2205 27895
rect 2291 27839 2347 27895
rect 2433 27839 2489 27895
rect 2575 27839 2631 27895
rect 2717 27839 2773 27895
rect 2859 27839 2915 27895
rect 3001 27839 3057 27895
rect 3143 27839 3199 27895
rect 3285 27839 3341 27895
rect 3427 27839 3483 27895
rect 3569 27839 3625 27895
rect 3711 27839 3767 27895
rect 3853 27839 3909 27895
rect 3995 27839 4051 27895
rect 4137 27839 4193 27895
rect 4279 27839 4335 27895
rect 4421 27839 4477 27895
rect 4563 27839 4619 27895
rect 4705 27839 4761 27895
rect 4847 27839 4903 27895
rect 4989 27839 5045 27895
rect 5131 27839 5187 27895
rect 5273 27839 5329 27895
rect 5415 27839 5471 27895
rect 5557 27839 5613 27895
rect 5699 27839 5755 27895
rect 5841 27839 5897 27895
rect 5983 27839 6039 27895
rect 6125 27839 6181 27895
rect 6267 27839 6323 27895
rect 6409 27839 6465 27895
rect 6551 27839 6607 27895
rect 6693 27839 6749 27895
rect 6835 27839 6891 27895
rect 6977 27839 7033 27895
rect 7119 27839 7175 27895
rect 7261 27839 7317 27895
rect 7403 27839 7459 27895
rect 7545 27839 7601 27895
rect 7687 27839 7743 27895
rect 7829 27839 7885 27895
rect 7971 27839 8027 27895
rect 8113 27839 8169 27895
rect 8255 27839 8311 27895
rect 8397 27839 8453 27895
rect 8539 27839 8595 27895
rect 8681 27839 8737 27895
rect 8823 27839 8879 27895
rect 8965 27839 9021 27895
rect 9107 27839 9163 27895
rect 9249 27839 9305 27895
rect 9391 27839 9447 27895
rect 9533 27839 9589 27895
rect 9675 27839 9731 27895
rect 9817 27839 9873 27895
rect 9959 27839 10015 27895
rect 10101 27839 10157 27895
rect 10243 27839 10299 27895
rect 10385 27839 10441 27895
rect 10527 27839 10583 27895
rect 10669 27839 10725 27895
rect 10811 27839 10867 27895
rect 10953 27839 11009 27895
rect 11095 27839 11151 27895
rect 11237 27839 11293 27895
rect 11379 27839 11435 27895
rect 11521 27839 11577 27895
rect 11663 27839 11719 27895
rect 11805 27839 11861 27895
rect 11947 27839 12003 27895
rect 12089 27839 12145 27895
rect 12231 27839 12287 27895
rect 12373 27839 12429 27895
rect 12515 27839 12571 27895
rect 12657 27839 12713 27895
rect 12799 27839 12855 27895
rect 12941 27839 12997 27895
rect 13083 27839 13139 27895
rect 13225 27839 13281 27895
rect 13367 27839 13423 27895
rect 13509 27839 13565 27895
rect 13651 27839 13707 27895
rect 13793 27839 13849 27895
rect 13935 27839 13991 27895
rect 14077 27839 14133 27895
rect 14219 27839 14275 27895
rect 14361 27839 14417 27895
rect 14503 27839 14559 27895
rect 14645 27839 14701 27895
rect 14787 27839 14843 27895
rect 161 27697 217 27753
rect 303 27697 359 27753
rect 445 27697 501 27753
rect 587 27697 643 27753
rect 729 27697 785 27753
rect 871 27697 927 27753
rect 1013 27697 1069 27753
rect 1155 27697 1211 27753
rect 1297 27697 1353 27753
rect 1439 27697 1495 27753
rect 1581 27697 1637 27753
rect 1723 27697 1779 27753
rect 1865 27697 1921 27753
rect 2007 27697 2063 27753
rect 2149 27697 2205 27753
rect 2291 27697 2347 27753
rect 2433 27697 2489 27753
rect 2575 27697 2631 27753
rect 2717 27697 2773 27753
rect 2859 27697 2915 27753
rect 3001 27697 3057 27753
rect 3143 27697 3199 27753
rect 3285 27697 3341 27753
rect 3427 27697 3483 27753
rect 3569 27697 3625 27753
rect 3711 27697 3767 27753
rect 3853 27697 3909 27753
rect 3995 27697 4051 27753
rect 4137 27697 4193 27753
rect 4279 27697 4335 27753
rect 4421 27697 4477 27753
rect 4563 27697 4619 27753
rect 4705 27697 4761 27753
rect 4847 27697 4903 27753
rect 4989 27697 5045 27753
rect 5131 27697 5187 27753
rect 5273 27697 5329 27753
rect 5415 27697 5471 27753
rect 5557 27697 5613 27753
rect 5699 27697 5755 27753
rect 5841 27697 5897 27753
rect 5983 27697 6039 27753
rect 6125 27697 6181 27753
rect 6267 27697 6323 27753
rect 6409 27697 6465 27753
rect 6551 27697 6607 27753
rect 6693 27697 6749 27753
rect 6835 27697 6891 27753
rect 6977 27697 7033 27753
rect 7119 27697 7175 27753
rect 7261 27697 7317 27753
rect 7403 27697 7459 27753
rect 7545 27697 7601 27753
rect 7687 27697 7743 27753
rect 7829 27697 7885 27753
rect 7971 27697 8027 27753
rect 8113 27697 8169 27753
rect 8255 27697 8311 27753
rect 8397 27697 8453 27753
rect 8539 27697 8595 27753
rect 8681 27697 8737 27753
rect 8823 27697 8879 27753
rect 8965 27697 9021 27753
rect 9107 27697 9163 27753
rect 9249 27697 9305 27753
rect 9391 27697 9447 27753
rect 9533 27697 9589 27753
rect 9675 27697 9731 27753
rect 9817 27697 9873 27753
rect 9959 27697 10015 27753
rect 10101 27697 10157 27753
rect 10243 27697 10299 27753
rect 10385 27697 10441 27753
rect 10527 27697 10583 27753
rect 10669 27697 10725 27753
rect 10811 27697 10867 27753
rect 10953 27697 11009 27753
rect 11095 27697 11151 27753
rect 11237 27697 11293 27753
rect 11379 27697 11435 27753
rect 11521 27697 11577 27753
rect 11663 27697 11719 27753
rect 11805 27697 11861 27753
rect 11947 27697 12003 27753
rect 12089 27697 12145 27753
rect 12231 27697 12287 27753
rect 12373 27697 12429 27753
rect 12515 27697 12571 27753
rect 12657 27697 12713 27753
rect 12799 27697 12855 27753
rect 12941 27697 12997 27753
rect 13083 27697 13139 27753
rect 13225 27697 13281 27753
rect 13367 27697 13423 27753
rect 13509 27697 13565 27753
rect 13651 27697 13707 27753
rect 13793 27697 13849 27753
rect 13935 27697 13991 27753
rect 14077 27697 14133 27753
rect 14219 27697 14275 27753
rect 14361 27697 14417 27753
rect 14503 27697 14559 27753
rect 14645 27697 14701 27753
rect 14787 27697 14843 27753
rect 161 27555 217 27611
rect 303 27555 359 27611
rect 445 27555 501 27611
rect 587 27555 643 27611
rect 729 27555 785 27611
rect 871 27555 927 27611
rect 1013 27555 1069 27611
rect 1155 27555 1211 27611
rect 1297 27555 1353 27611
rect 1439 27555 1495 27611
rect 1581 27555 1637 27611
rect 1723 27555 1779 27611
rect 1865 27555 1921 27611
rect 2007 27555 2063 27611
rect 2149 27555 2205 27611
rect 2291 27555 2347 27611
rect 2433 27555 2489 27611
rect 2575 27555 2631 27611
rect 2717 27555 2773 27611
rect 2859 27555 2915 27611
rect 3001 27555 3057 27611
rect 3143 27555 3199 27611
rect 3285 27555 3341 27611
rect 3427 27555 3483 27611
rect 3569 27555 3625 27611
rect 3711 27555 3767 27611
rect 3853 27555 3909 27611
rect 3995 27555 4051 27611
rect 4137 27555 4193 27611
rect 4279 27555 4335 27611
rect 4421 27555 4477 27611
rect 4563 27555 4619 27611
rect 4705 27555 4761 27611
rect 4847 27555 4903 27611
rect 4989 27555 5045 27611
rect 5131 27555 5187 27611
rect 5273 27555 5329 27611
rect 5415 27555 5471 27611
rect 5557 27555 5613 27611
rect 5699 27555 5755 27611
rect 5841 27555 5897 27611
rect 5983 27555 6039 27611
rect 6125 27555 6181 27611
rect 6267 27555 6323 27611
rect 6409 27555 6465 27611
rect 6551 27555 6607 27611
rect 6693 27555 6749 27611
rect 6835 27555 6891 27611
rect 6977 27555 7033 27611
rect 7119 27555 7175 27611
rect 7261 27555 7317 27611
rect 7403 27555 7459 27611
rect 7545 27555 7601 27611
rect 7687 27555 7743 27611
rect 7829 27555 7885 27611
rect 7971 27555 8027 27611
rect 8113 27555 8169 27611
rect 8255 27555 8311 27611
rect 8397 27555 8453 27611
rect 8539 27555 8595 27611
rect 8681 27555 8737 27611
rect 8823 27555 8879 27611
rect 8965 27555 9021 27611
rect 9107 27555 9163 27611
rect 9249 27555 9305 27611
rect 9391 27555 9447 27611
rect 9533 27555 9589 27611
rect 9675 27555 9731 27611
rect 9817 27555 9873 27611
rect 9959 27555 10015 27611
rect 10101 27555 10157 27611
rect 10243 27555 10299 27611
rect 10385 27555 10441 27611
rect 10527 27555 10583 27611
rect 10669 27555 10725 27611
rect 10811 27555 10867 27611
rect 10953 27555 11009 27611
rect 11095 27555 11151 27611
rect 11237 27555 11293 27611
rect 11379 27555 11435 27611
rect 11521 27555 11577 27611
rect 11663 27555 11719 27611
rect 11805 27555 11861 27611
rect 11947 27555 12003 27611
rect 12089 27555 12145 27611
rect 12231 27555 12287 27611
rect 12373 27555 12429 27611
rect 12515 27555 12571 27611
rect 12657 27555 12713 27611
rect 12799 27555 12855 27611
rect 12941 27555 12997 27611
rect 13083 27555 13139 27611
rect 13225 27555 13281 27611
rect 13367 27555 13423 27611
rect 13509 27555 13565 27611
rect 13651 27555 13707 27611
rect 13793 27555 13849 27611
rect 13935 27555 13991 27611
rect 14077 27555 14133 27611
rect 14219 27555 14275 27611
rect 14361 27555 14417 27611
rect 14503 27555 14559 27611
rect 14645 27555 14701 27611
rect 14787 27555 14843 27611
rect 161 27413 217 27469
rect 303 27413 359 27469
rect 445 27413 501 27469
rect 587 27413 643 27469
rect 729 27413 785 27469
rect 871 27413 927 27469
rect 1013 27413 1069 27469
rect 1155 27413 1211 27469
rect 1297 27413 1353 27469
rect 1439 27413 1495 27469
rect 1581 27413 1637 27469
rect 1723 27413 1779 27469
rect 1865 27413 1921 27469
rect 2007 27413 2063 27469
rect 2149 27413 2205 27469
rect 2291 27413 2347 27469
rect 2433 27413 2489 27469
rect 2575 27413 2631 27469
rect 2717 27413 2773 27469
rect 2859 27413 2915 27469
rect 3001 27413 3057 27469
rect 3143 27413 3199 27469
rect 3285 27413 3341 27469
rect 3427 27413 3483 27469
rect 3569 27413 3625 27469
rect 3711 27413 3767 27469
rect 3853 27413 3909 27469
rect 3995 27413 4051 27469
rect 4137 27413 4193 27469
rect 4279 27413 4335 27469
rect 4421 27413 4477 27469
rect 4563 27413 4619 27469
rect 4705 27413 4761 27469
rect 4847 27413 4903 27469
rect 4989 27413 5045 27469
rect 5131 27413 5187 27469
rect 5273 27413 5329 27469
rect 5415 27413 5471 27469
rect 5557 27413 5613 27469
rect 5699 27413 5755 27469
rect 5841 27413 5897 27469
rect 5983 27413 6039 27469
rect 6125 27413 6181 27469
rect 6267 27413 6323 27469
rect 6409 27413 6465 27469
rect 6551 27413 6607 27469
rect 6693 27413 6749 27469
rect 6835 27413 6891 27469
rect 6977 27413 7033 27469
rect 7119 27413 7175 27469
rect 7261 27413 7317 27469
rect 7403 27413 7459 27469
rect 7545 27413 7601 27469
rect 7687 27413 7743 27469
rect 7829 27413 7885 27469
rect 7971 27413 8027 27469
rect 8113 27413 8169 27469
rect 8255 27413 8311 27469
rect 8397 27413 8453 27469
rect 8539 27413 8595 27469
rect 8681 27413 8737 27469
rect 8823 27413 8879 27469
rect 8965 27413 9021 27469
rect 9107 27413 9163 27469
rect 9249 27413 9305 27469
rect 9391 27413 9447 27469
rect 9533 27413 9589 27469
rect 9675 27413 9731 27469
rect 9817 27413 9873 27469
rect 9959 27413 10015 27469
rect 10101 27413 10157 27469
rect 10243 27413 10299 27469
rect 10385 27413 10441 27469
rect 10527 27413 10583 27469
rect 10669 27413 10725 27469
rect 10811 27413 10867 27469
rect 10953 27413 11009 27469
rect 11095 27413 11151 27469
rect 11237 27413 11293 27469
rect 11379 27413 11435 27469
rect 11521 27413 11577 27469
rect 11663 27413 11719 27469
rect 11805 27413 11861 27469
rect 11947 27413 12003 27469
rect 12089 27413 12145 27469
rect 12231 27413 12287 27469
rect 12373 27413 12429 27469
rect 12515 27413 12571 27469
rect 12657 27413 12713 27469
rect 12799 27413 12855 27469
rect 12941 27413 12997 27469
rect 13083 27413 13139 27469
rect 13225 27413 13281 27469
rect 13367 27413 13423 27469
rect 13509 27413 13565 27469
rect 13651 27413 13707 27469
rect 13793 27413 13849 27469
rect 13935 27413 13991 27469
rect 14077 27413 14133 27469
rect 14219 27413 14275 27469
rect 14361 27413 14417 27469
rect 14503 27413 14559 27469
rect 14645 27413 14701 27469
rect 14787 27413 14843 27469
rect 161 27271 217 27327
rect 303 27271 359 27327
rect 445 27271 501 27327
rect 587 27271 643 27327
rect 729 27271 785 27327
rect 871 27271 927 27327
rect 1013 27271 1069 27327
rect 1155 27271 1211 27327
rect 1297 27271 1353 27327
rect 1439 27271 1495 27327
rect 1581 27271 1637 27327
rect 1723 27271 1779 27327
rect 1865 27271 1921 27327
rect 2007 27271 2063 27327
rect 2149 27271 2205 27327
rect 2291 27271 2347 27327
rect 2433 27271 2489 27327
rect 2575 27271 2631 27327
rect 2717 27271 2773 27327
rect 2859 27271 2915 27327
rect 3001 27271 3057 27327
rect 3143 27271 3199 27327
rect 3285 27271 3341 27327
rect 3427 27271 3483 27327
rect 3569 27271 3625 27327
rect 3711 27271 3767 27327
rect 3853 27271 3909 27327
rect 3995 27271 4051 27327
rect 4137 27271 4193 27327
rect 4279 27271 4335 27327
rect 4421 27271 4477 27327
rect 4563 27271 4619 27327
rect 4705 27271 4761 27327
rect 4847 27271 4903 27327
rect 4989 27271 5045 27327
rect 5131 27271 5187 27327
rect 5273 27271 5329 27327
rect 5415 27271 5471 27327
rect 5557 27271 5613 27327
rect 5699 27271 5755 27327
rect 5841 27271 5897 27327
rect 5983 27271 6039 27327
rect 6125 27271 6181 27327
rect 6267 27271 6323 27327
rect 6409 27271 6465 27327
rect 6551 27271 6607 27327
rect 6693 27271 6749 27327
rect 6835 27271 6891 27327
rect 6977 27271 7033 27327
rect 7119 27271 7175 27327
rect 7261 27271 7317 27327
rect 7403 27271 7459 27327
rect 7545 27271 7601 27327
rect 7687 27271 7743 27327
rect 7829 27271 7885 27327
rect 7971 27271 8027 27327
rect 8113 27271 8169 27327
rect 8255 27271 8311 27327
rect 8397 27271 8453 27327
rect 8539 27271 8595 27327
rect 8681 27271 8737 27327
rect 8823 27271 8879 27327
rect 8965 27271 9021 27327
rect 9107 27271 9163 27327
rect 9249 27271 9305 27327
rect 9391 27271 9447 27327
rect 9533 27271 9589 27327
rect 9675 27271 9731 27327
rect 9817 27271 9873 27327
rect 9959 27271 10015 27327
rect 10101 27271 10157 27327
rect 10243 27271 10299 27327
rect 10385 27271 10441 27327
rect 10527 27271 10583 27327
rect 10669 27271 10725 27327
rect 10811 27271 10867 27327
rect 10953 27271 11009 27327
rect 11095 27271 11151 27327
rect 11237 27271 11293 27327
rect 11379 27271 11435 27327
rect 11521 27271 11577 27327
rect 11663 27271 11719 27327
rect 11805 27271 11861 27327
rect 11947 27271 12003 27327
rect 12089 27271 12145 27327
rect 12231 27271 12287 27327
rect 12373 27271 12429 27327
rect 12515 27271 12571 27327
rect 12657 27271 12713 27327
rect 12799 27271 12855 27327
rect 12941 27271 12997 27327
rect 13083 27271 13139 27327
rect 13225 27271 13281 27327
rect 13367 27271 13423 27327
rect 13509 27271 13565 27327
rect 13651 27271 13707 27327
rect 13793 27271 13849 27327
rect 13935 27271 13991 27327
rect 14077 27271 14133 27327
rect 14219 27271 14275 27327
rect 14361 27271 14417 27327
rect 14503 27271 14559 27327
rect 14645 27271 14701 27327
rect 14787 27271 14843 27327
rect 161 27129 217 27185
rect 303 27129 359 27185
rect 445 27129 501 27185
rect 587 27129 643 27185
rect 729 27129 785 27185
rect 871 27129 927 27185
rect 1013 27129 1069 27185
rect 1155 27129 1211 27185
rect 1297 27129 1353 27185
rect 1439 27129 1495 27185
rect 1581 27129 1637 27185
rect 1723 27129 1779 27185
rect 1865 27129 1921 27185
rect 2007 27129 2063 27185
rect 2149 27129 2205 27185
rect 2291 27129 2347 27185
rect 2433 27129 2489 27185
rect 2575 27129 2631 27185
rect 2717 27129 2773 27185
rect 2859 27129 2915 27185
rect 3001 27129 3057 27185
rect 3143 27129 3199 27185
rect 3285 27129 3341 27185
rect 3427 27129 3483 27185
rect 3569 27129 3625 27185
rect 3711 27129 3767 27185
rect 3853 27129 3909 27185
rect 3995 27129 4051 27185
rect 4137 27129 4193 27185
rect 4279 27129 4335 27185
rect 4421 27129 4477 27185
rect 4563 27129 4619 27185
rect 4705 27129 4761 27185
rect 4847 27129 4903 27185
rect 4989 27129 5045 27185
rect 5131 27129 5187 27185
rect 5273 27129 5329 27185
rect 5415 27129 5471 27185
rect 5557 27129 5613 27185
rect 5699 27129 5755 27185
rect 5841 27129 5897 27185
rect 5983 27129 6039 27185
rect 6125 27129 6181 27185
rect 6267 27129 6323 27185
rect 6409 27129 6465 27185
rect 6551 27129 6607 27185
rect 6693 27129 6749 27185
rect 6835 27129 6891 27185
rect 6977 27129 7033 27185
rect 7119 27129 7175 27185
rect 7261 27129 7317 27185
rect 7403 27129 7459 27185
rect 7545 27129 7601 27185
rect 7687 27129 7743 27185
rect 7829 27129 7885 27185
rect 7971 27129 8027 27185
rect 8113 27129 8169 27185
rect 8255 27129 8311 27185
rect 8397 27129 8453 27185
rect 8539 27129 8595 27185
rect 8681 27129 8737 27185
rect 8823 27129 8879 27185
rect 8965 27129 9021 27185
rect 9107 27129 9163 27185
rect 9249 27129 9305 27185
rect 9391 27129 9447 27185
rect 9533 27129 9589 27185
rect 9675 27129 9731 27185
rect 9817 27129 9873 27185
rect 9959 27129 10015 27185
rect 10101 27129 10157 27185
rect 10243 27129 10299 27185
rect 10385 27129 10441 27185
rect 10527 27129 10583 27185
rect 10669 27129 10725 27185
rect 10811 27129 10867 27185
rect 10953 27129 11009 27185
rect 11095 27129 11151 27185
rect 11237 27129 11293 27185
rect 11379 27129 11435 27185
rect 11521 27129 11577 27185
rect 11663 27129 11719 27185
rect 11805 27129 11861 27185
rect 11947 27129 12003 27185
rect 12089 27129 12145 27185
rect 12231 27129 12287 27185
rect 12373 27129 12429 27185
rect 12515 27129 12571 27185
rect 12657 27129 12713 27185
rect 12799 27129 12855 27185
rect 12941 27129 12997 27185
rect 13083 27129 13139 27185
rect 13225 27129 13281 27185
rect 13367 27129 13423 27185
rect 13509 27129 13565 27185
rect 13651 27129 13707 27185
rect 13793 27129 13849 27185
rect 13935 27129 13991 27185
rect 14077 27129 14133 27185
rect 14219 27129 14275 27185
rect 14361 27129 14417 27185
rect 14503 27129 14559 27185
rect 14645 27129 14701 27185
rect 14787 27129 14843 27185
rect 161 26987 217 27043
rect 303 26987 359 27043
rect 445 26987 501 27043
rect 587 26987 643 27043
rect 729 26987 785 27043
rect 871 26987 927 27043
rect 1013 26987 1069 27043
rect 1155 26987 1211 27043
rect 1297 26987 1353 27043
rect 1439 26987 1495 27043
rect 1581 26987 1637 27043
rect 1723 26987 1779 27043
rect 1865 26987 1921 27043
rect 2007 26987 2063 27043
rect 2149 26987 2205 27043
rect 2291 26987 2347 27043
rect 2433 26987 2489 27043
rect 2575 26987 2631 27043
rect 2717 26987 2773 27043
rect 2859 26987 2915 27043
rect 3001 26987 3057 27043
rect 3143 26987 3199 27043
rect 3285 26987 3341 27043
rect 3427 26987 3483 27043
rect 3569 26987 3625 27043
rect 3711 26987 3767 27043
rect 3853 26987 3909 27043
rect 3995 26987 4051 27043
rect 4137 26987 4193 27043
rect 4279 26987 4335 27043
rect 4421 26987 4477 27043
rect 4563 26987 4619 27043
rect 4705 26987 4761 27043
rect 4847 26987 4903 27043
rect 4989 26987 5045 27043
rect 5131 26987 5187 27043
rect 5273 26987 5329 27043
rect 5415 26987 5471 27043
rect 5557 26987 5613 27043
rect 5699 26987 5755 27043
rect 5841 26987 5897 27043
rect 5983 26987 6039 27043
rect 6125 26987 6181 27043
rect 6267 26987 6323 27043
rect 6409 26987 6465 27043
rect 6551 26987 6607 27043
rect 6693 26987 6749 27043
rect 6835 26987 6891 27043
rect 6977 26987 7033 27043
rect 7119 26987 7175 27043
rect 7261 26987 7317 27043
rect 7403 26987 7459 27043
rect 7545 26987 7601 27043
rect 7687 26987 7743 27043
rect 7829 26987 7885 27043
rect 7971 26987 8027 27043
rect 8113 26987 8169 27043
rect 8255 26987 8311 27043
rect 8397 26987 8453 27043
rect 8539 26987 8595 27043
rect 8681 26987 8737 27043
rect 8823 26987 8879 27043
rect 8965 26987 9021 27043
rect 9107 26987 9163 27043
rect 9249 26987 9305 27043
rect 9391 26987 9447 27043
rect 9533 26987 9589 27043
rect 9675 26987 9731 27043
rect 9817 26987 9873 27043
rect 9959 26987 10015 27043
rect 10101 26987 10157 27043
rect 10243 26987 10299 27043
rect 10385 26987 10441 27043
rect 10527 26987 10583 27043
rect 10669 26987 10725 27043
rect 10811 26987 10867 27043
rect 10953 26987 11009 27043
rect 11095 26987 11151 27043
rect 11237 26987 11293 27043
rect 11379 26987 11435 27043
rect 11521 26987 11577 27043
rect 11663 26987 11719 27043
rect 11805 26987 11861 27043
rect 11947 26987 12003 27043
rect 12089 26987 12145 27043
rect 12231 26987 12287 27043
rect 12373 26987 12429 27043
rect 12515 26987 12571 27043
rect 12657 26987 12713 27043
rect 12799 26987 12855 27043
rect 12941 26987 12997 27043
rect 13083 26987 13139 27043
rect 13225 26987 13281 27043
rect 13367 26987 13423 27043
rect 13509 26987 13565 27043
rect 13651 26987 13707 27043
rect 13793 26987 13849 27043
rect 13935 26987 13991 27043
rect 14077 26987 14133 27043
rect 14219 26987 14275 27043
rect 14361 26987 14417 27043
rect 14503 26987 14559 27043
rect 14645 26987 14701 27043
rect 14787 26987 14843 27043
rect 161 26845 217 26901
rect 303 26845 359 26901
rect 445 26845 501 26901
rect 587 26845 643 26901
rect 729 26845 785 26901
rect 871 26845 927 26901
rect 1013 26845 1069 26901
rect 1155 26845 1211 26901
rect 1297 26845 1353 26901
rect 1439 26845 1495 26901
rect 1581 26845 1637 26901
rect 1723 26845 1779 26901
rect 1865 26845 1921 26901
rect 2007 26845 2063 26901
rect 2149 26845 2205 26901
rect 2291 26845 2347 26901
rect 2433 26845 2489 26901
rect 2575 26845 2631 26901
rect 2717 26845 2773 26901
rect 2859 26845 2915 26901
rect 3001 26845 3057 26901
rect 3143 26845 3199 26901
rect 3285 26845 3341 26901
rect 3427 26845 3483 26901
rect 3569 26845 3625 26901
rect 3711 26845 3767 26901
rect 3853 26845 3909 26901
rect 3995 26845 4051 26901
rect 4137 26845 4193 26901
rect 4279 26845 4335 26901
rect 4421 26845 4477 26901
rect 4563 26845 4619 26901
rect 4705 26845 4761 26901
rect 4847 26845 4903 26901
rect 4989 26845 5045 26901
rect 5131 26845 5187 26901
rect 5273 26845 5329 26901
rect 5415 26845 5471 26901
rect 5557 26845 5613 26901
rect 5699 26845 5755 26901
rect 5841 26845 5897 26901
rect 5983 26845 6039 26901
rect 6125 26845 6181 26901
rect 6267 26845 6323 26901
rect 6409 26845 6465 26901
rect 6551 26845 6607 26901
rect 6693 26845 6749 26901
rect 6835 26845 6891 26901
rect 6977 26845 7033 26901
rect 7119 26845 7175 26901
rect 7261 26845 7317 26901
rect 7403 26845 7459 26901
rect 7545 26845 7601 26901
rect 7687 26845 7743 26901
rect 7829 26845 7885 26901
rect 7971 26845 8027 26901
rect 8113 26845 8169 26901
rect 8255 26845 8311 26901
rect 8397 26845 8453 26901
rect 8539 26845 8595 26901
rect 8681 26845 8737 26901
rect 8823 26845 8879 26901
rect 8965 26845 9021 26901
rect 9107 26845 9163 26901
rect 9249 26845 9305 26901
rect 9391 26845 9447 26901
rect 9533 26845 9589 26901
rect 9675 26845 9731 26901
rect 9817 26845 9873 26901
rect 9959 26845 10015 26901
rect 10101 26845 10157 26901
rect 10243 26845 10299 26901
rect 10385 26845 10441 26901
rect 10527 26845 10583 26901
rect 10669 26845 10725 26901
rect 10811 26845 10867 26901
rect 10953 26845 11009 26901
rect 11095 26845 11151 26901
rect 11237 26845 11293 26901
rect 11379 26845 11435 26901
rect 11521 26845 11577 26901
rect 11663 26845 11719 26901
rect 11805 26845 11861 26901
rect 11947 26845 12003 26901
rect 12089 26845 12145 26901
rect 12231 26845 12287 26901
rect 12373 26845 12429 26901
rect 12515 26845 12571 26901
rect 12657 26845 12713 26901
rect 12799 26845 12855 26901
rect 12941 26845 12997 26901
rect 13083 26845 13139 26901
rect 13225 26845 13281 26901
rect 13367 26845 13423 26901
rect 13509 26845 13565 26901
rect 13651 26845 13707 26901
rect 13793 26845 13849 26901
rect 13935 26845 13991 26901
rect 14077 26845 14133 26901
rect 14219 26845 14275 26901
rect 14361 26845 14417 26901
rect 14503 26845 14559 26901
rect 14645 26845 14701 26901
rect 14787 26845 14843 26901
rect 161 26507 217 26563
rect 303 26507 359 26563
rect 445 26507 501 26563
rect 587 26507 643 26563
rect 729 26507 785 26563
rect 871 26507 927 26563
rect 1013 26507 1069 26563
rect 1155 26507 1211 26563
rect 1297 26507 1353 26563
rect 1439 26507 1495 26563
rect 1581 26507 1637 26563
rect 1723 26507 1779 26563
rect 1865 26507 1921 26563
rect 2007 26507 2063 26563
rect 2149 26507 2205 26563
rect 2291 26507 2347 26563
rect 2433 26507 2489 26563
rect 2575 26507 2631 26563
rect 2717 26507 2773 26563
rect 2859 26507 2915 26563
rect 3001 26507 3057 26563
rect 3143 26507 3199 26563
rect 3285 26507 3341 26563
rect 3427 26507 3483 26563
rect 3569 26507 3625 26563
rect 3711 26507 3767 26563
rect 3853 26507 3909 26563
rect 3995 26507 4051 26563
rect 4137 26507 4193 26563
rect 4279 26507 4335 26563
rect 4421 26507 4477 26563
rect 4563 26507 4619 26563
rect 4705 26507 4761 26563
rect 4847 26507 4903 26563
rect 4989 26507 5045 26563
rect 5131 26507 5187 26563
rect 5273 26507 5329 26563
rect 5415 26507 5471 26563
rect 5557 26507 5613 26563
rect 5699 26507 5755 26563
rect 5841 26507 5897 26563
rect 5983 26507 6039 26563
rect 6125 26507 6181 26563
rect 6267 26507 6323 26563
rect 6409 26507 6465 26563
rect 6551 26507 6607 26563
rect 6693 26507 6749 26563
rect 6835 26507 6891 26563
rect 6977 26507 7033 26563
rect 7119 26507 7175 26563
rect 7261 26507 7317 26563
rect 7403 26507 7459 26563
rect 7545 26507 7601 26563
rect 7687 26507 7743 26563
rect 7829 26507 7885 26563
rect 7971 26507 8027 26563
rect 8113 26507 8169 26563
rect 8255 26507 8311 26563
rect 8397 26507 8453 26563
rect 8539 26507 8595 26563
rect 8681 26507 8737 26563
rect 8823 26507 8879 26563
rect 8965 26507 9021 26563
rect 9107 26507 9163 26563
rect 9249 26507 9305 26563
rect 9391 26507 9447 26563
rect 9533 26507 9589 26563
rect 9675 26507 9731 26563
rect 9817 26507 9873 26563
rect 9959 26507 10015 26563
rect 10101 26507 10157 26563
rect 10243 26507 10299 26563
rect 10385 26507 10441 26563
rect 10527 26507 10583 26563
rect 10669 26507 10725 26563
rect 10811 26507 10867 26563
rect 10953 26507 11009 26563
rect 11095 26507 11151 26563
rect 11237 26507 11293 26563
rect 11379 26507 11435 26563
rect 11521 26507 11577 26563
rect 11663 26507 11719 26563
rect 11805 26507 11861 26563
rect 11947 26507 12003 26563
rect 12089 26507 12145 26563
rect 12231 26507 12287 26563
rect 12373 26507 12429 26563
rect 12515 26507 12571 26563
rect 12657 26507 12713 26563
rect 12799 26507 12855 26563
rect 12941 26507 12997 26563
rect 13083 26507 13139 26563
rect 13225 26507 13281 26563
rect 13367 26507 13423 26563
rect 13509 26507 13565 26563
rect 13651 26507 13707 26563
rect 13793 26507 13849 26563
rect 13935 26507 13991 26563
rect 14077 26507 14133 26563
rect 14219 26507 14275 26563
rect 14361 26507 14417 26563
rect 14503 26507 14559 26563
rect 14645 26507 14701 26563
rect 14787 26507 14843 26563
rect 161 26365 217 26421
rect 303 26365 359 26421
rect 445 26365 501 26421
rect 587 26365 643 26421
rect 729 26365 785 26421
rect 871 26365 927 26421
rect 1013 26365 1069 26421
rect 1155 26365 1211 26421
rect 1297 26365 1353 26421
rect 1439 26365 1495 26421
rect 1581 26365 1637 26421
rect 1723 26365 1779 26421
rect 1865 26365 1921 26421
rect 2007 26365 2063 26421
rect 2149 26365 2205 26421
rect 2291 26365 2347 26421
rect 2433 26365 2489 26421
rect 2575 26365 2631 26421
rect 2717 26365 2773 26421
rect 2859 26365 2915 26421
rect 3001 26365 3057 26421
rect 3143 26365 3199 26421
rect 3285 26365 3341 26421
rect 3427 26365 3483 26421
rect 3569 26365 3625 26421
rect 3711 26365 3767 26421
rect 3853 26365 3909 26421
rect 3995 26365 4051 26421
rect 4137 26365 4193 26421
rect 4279 26365 4335 26421
rect 4421 26365 4477 26421
rect 4563 26365 4619 26421
rect 4705 26365 4761 26421
rect 4847 26365 4903 26421
rect 4989 26365 5045 26421
rect 5131 26365 5187 26421
rect 5273 26365 5329 26421
rect 5415 26365 5471 26421
rect 5557 26365 5613 26421
rect 5699 26365 5755 26421
rect 5841 26365 5897 26421
rect 5983 26365 6039 26421
rect 6125 26365 6181 26421
rect 6267 26365 6323 26421
rect 6409 26365 6465 26421
rect 6551 26365 6607 26421
rect 6693 26365 6749 26421
rect 6835 26365 6891 26421
rect 6977 26365 7033 26421
rect 7119 26365 7175 26421
rect 7261 26365 7317 26421
rect 7403 26365 7459 26421
rect 7545 26365 7601 26421
rect 7687 26365 7743 26421
rect 7829 26365 7885 26421
rect 7971 26365 8027 26421
rect 8113 26365 8169 26421
rect 8255 26365 8311 26421
rect 8397 26365 8453 26421
rect 8539 26365 8595 26421
rect 8681 26365 8737 26421
rect 8823 26365 8879 26421
rect 8965 26365 9021 26421
rect 9107 26365 9163 26421
rect 9249 26365 9305 26421
rect 9391 26365 9447 26421
rect 9533 26365 9589 26421
rect 9675 26365 9731 26421
rect 9817 26365 9873 26421
rect 9959 26365 10015 26421
rect 10101 26365 10157 26421
rect 10243 26365 10299 26421
rect 10385 26365 10441 26421
rect 10527 26365 10583 26421
rect 10669 26365 10725 26421
rect 10811 26365 10867 26421
rect 10953 26365 11009 26421
rect 11095 26365 11151 26421
rect 11237 26365 11293 26421
rect 11379 26365 11435 26421
rect 11521 26365 11577 26421
rect 11663 26365 11719 26421
rect 11805 26365 11861 26421
rect 11947 26365 12003 26421
rect 12089 26365 12145 26421
rect 12231 26365 12287 26421
rect 12373 26365 12429 26421
rect 12515 26365 12571 26421
rect 12657 26365 12713 26421
rect 12799 26365 12855 26421
rect 12941 26365 12997 26421
rect 13083 26365 13139 26421
rect 13225 26365 13281 26421
rect 13367 26365 13423 26421
rect 13509 26365 13565 26421
rect 13651 26365 13707 26421
rect 13793 26365 13849 26421
rect 13935 26365 13991 26421
rect 14077 26365 14133 26421
rect 14219 26365 14275 26421
rect 14361 26365 14417 26421
rect 14503 26365 14559 26421
rect 14645 26365 14701 26421
rect 14787 26365 14843 26421
rect 161 26223 217 26279
rect 303 26223 359 26279
rect 445 26223 501 26279
rect 587 26223 643 26279
rect 729 26223 785 26279
rect 871 26223 927 26279
rect 1013 26223 1069 26279
rect 1155 26223 1211 26279
rect 1297 26223 1353 26279
rect 1439 26223 1495 26279
rect 1581 26223 1637 26279
rect 1723 26223 1779 26279
rect 1865 26223 1921 26279
rect 2007 26223 2063 26279
rect 2149 26223 2205 26279
rect 2291 26223 2347 26279
rect 2433 26223 2489 26279
rect 2575 26223 2631 26279
rect 2717 26223 2773 26279
rect 2859 26223 2915 26279
rect 3001 26223 3057 26279
rect 3143 26223 3199 26279
rect 3285 26223 3341 26279
rect 3427 26223 3483 26279
rect 3569 26223 3625 26279
rect 3711 26223 3767 26279
rect 3853 26223 3909 26279
rect 3995 26223 4051 26279
rect 4137 26223 4193 26279
rect 4279 26223 4335 26279
rect 4421 26223 4477 26279
rect 4563 26223 4619 26279
rect 4705 26223 4761 26279
rect 4847 26223 4903 26279
rect 4989 26223 5045 26279
rect 5131 26223 5187 26279
rect 5273 26223 5329 26279
rect 5415 26223 5471 26279
rect 5557 26223 5613 26279
rect 5699 26223 5755 26279
rect 5841 26223 5897 26279
rect 5983 26223 6039 26279
rect 6125 26223 6181 26279
rect 6267 26223 6323 26279
rect 6409 26223 6465 26279
rect 6551 26223 6607 26279
rect 6693 26223 6749 26279
rect 6835 26223 6891 26279
rect 6977 26223 7033 26279
rect 7119 26223 7175 26279
rect 7261 26223 7317 26279
rect 7403 26223 7459 26279
rect 7545 26223 7601 26279
rect 7687 26223 7743 26279
rect 7829 26223 7885 26279
rect 7971 26223 8027 26279
rect 8113 26223 8169 26279
rect 8255 26223 8311 26279
rect 8397 26223 8453 26279
rect 8539 26223 8595 26279
rect 8681 26223 8737 26279
rect 8823 26223 8879 26279
rect 8965 26223 9021 26279
rect 9107 26223 9163 26279
rect 9249 26223 9305 26279
rect 9391 26223 9447 26279
rect 9533 26223 9589 26279
rect 9675 26223 9731 26279
rect 9817 26223 9873 26279
rect 9959 26223 10015 26279
rect 10101 26223 10157 26279
rect 10243 26223 10299 26279
rect 10385 26223 10441 26279
rect 10527 26223 10583 26279
rect 10669 26223 10725 26279
rect 10811 26223 10867 26279
rect 10953 26223 11009 26279
rect 11095 26223 11151 26279
rect 11237 26223 11293 26279
rect 11379 26223 11435 26279
rect 11521 26223 11577 26279
rect 11663 26223 11719 26279
rect 11805 26223 11861 26279
rect 11947 26223 12003 26279
rect 12089 26223 12145 26279
rect 12231 26223 12287 26279
rect 12373 26223 12429 26279
rect 12515 26223 12571 26279
rect 12657 26223 12713 26279
rect 12799 26223 12855 26279
rect 12941 26223 12997 26279
rect 13083 26223 13139 26279
rect 13225 26223 13281 26279
rect 13367 26223 13423 26279
rect 13509 26223 13565 26279
rect 13651 26223 13707 26279
rect 13793 26223 13849 26279
rect 13935 26223 13991 26279
rect 14077 26223 14133 26279
rect 14219 26223 14275 26279
rect 14361 26223 14417 26279
rect 14503 26223 14559 26279
rect 14645 26223 14701 26279
rect 14787 26223 14843 26279
rect 161 26081 217 26137
rect 303 26081 359 26137
rect 445 26081 501 26137
rect 587 26081 643 26137
rect 729 26081 785 26137
rect 871 26081 927 26137
rect 1013 26081 1069 26137
rect 1155 26081 1211 26137
rect 1297 26081 1353 26137
rect 1439 26081 1495 26137
rect 1581 26081 1637 26137
rect 1723 26081 1779 26137
rect 1865 26081 1921 26137
rect 2007 26081 2063 26137
rect 2149 26081 2205 26137
rect 2291 26081 2347 26137
rect 2433 26081 2489 26137
rect 2575 26081 2631 26137
rect 2717 26081 2773 26137
rect 2859 26081 2915 26137
rect 3001 26081 3057 26137
rect 3143 26081 3199 26137
rect 3285 26081 3341 26137
rect 3427 26081 3483 26137
rect 3569 26081 3625 26137
rect 3711 26081 3767 26137
rect 3853 26081 3909 26137
rect 3995 26081 4051 26137
rect 4137 26081 4193 26137
rect 4279 26081 4335 26137
rect 4421 26081 4477 26137
rect 4563 26081 4619 26137
rect 4705 26081 4761 26137
rect 4847 26081 4903 26137
rect 4989 26081 5045 26137
rect 5131 26081 5187 26137
rect 5273 26081 5329 26137
rect 5415 26081 5471 26137
rect 5557 26081 5613 26137
rect 5699 26081 5755 26137
rect 5841 26081 5897 26137
rect 5983 26081 6039 26137
rect 6125 26081 6181 26137
rect 6267 26081 6323 26137
rect 6409 26081 6465 26137
rect 6551 26081 6607 26137
rect 6693 26081 6749 26137
rect 6835 26081 6891 26137
rect 6977 26081 7033 26137
rect 7119 26081 7175 26137
rect 7261 26081 7317 26137
rect 7403 26081 7459 26137
rect 7545 26081 7601 26137
rect 7687 26081 7743 26137
rect 7829 26081 7885 26137
rect 7971 26081 8027 26137
rect 8113 26081 8169 26137
rect 8255 26081 8311 26137
rect 8397 26081 8453 26137
rect 8539 26081 8595 26137
rect 8681 26081 8737 26137
rect 8823 26081 8879 26137
rect 8965 26081 9021 26137
rect 9107 26081 9163 26137
rect 9249 26081 9305 26137
rect 9391 26081 9447 26137
rect 9533 26081 9589 26137
rect 9675 26081 9731 26137
rect 9817 26081 9873 26137
rect 9959 26081 10015 26137
rect 10101 26081 10157 26137
rect 10243 26081 10299 26137
rect 10385 26081 10441 26137
rect 10527 26081 10583 26137
rect 10669 26081 10725 26137
rect 10811 26081 10867 26137
rect 10953 26081 11009 26137
rect 11095 26081 11151 26137
rect 11237 26081 11293 26137
rect 11379 26081 11435 26137
rect 11521 26081 11577 26137
rect 11663 26081 11719 26137
rect 11805 26081 11861 26137
rect 11947 26081 12003 26137
rect 12089 26081 12145 26137
rect 12231 26081 12287 26137
rect 12373 26081 12429 26137
rect 12515 26081 12571 26137
rect 12657 26081 12713 26137
rect 12799 26081 12855 26137
rect 12941 26081 12997 26137
rect 13083 26081 13139 26137
rect 13225 26081 13281 26137
rect 13367 26081 13423 26137
rect 13509 26081 13565 26137
rect 13651 26081 13707 26137
rect 13793 26081 13849 26137
rect 13935 26081 13991 26137
rect 14077 26081 14133 26137
rect 14219 26081 14275 26137
rect 14361 26081 14417 26137
rect 14503 26081 14559 26137
rect 14645 26081 14701 26137
rect 14787 26081 14843 26137
rect 161 25939 217 25995
rect 303 25939 359 25995
rect 445 25939 501 25995
rect 587 25939 643 25995
rect 729 25939 785 25995
rect 871 25939 927 25995
rect 1013 25939 1069 25995
rect 1155 25939 1211 25995
rect 1297 25939 1353 25995
rect 1439 25939 1495 25995
rect 1581 25939 1637 25995
rect 1723 25939 1779 25995
rect 1865 25939 1921 25995
rect 2007 25939 2063 25995
rect 2149 25939 2205 25995
rect 2291 25939 2347 25995
rect 2433 25939 2489 25995
rect 2575 25939 2631 25995
rect 2717 25939 2773 25995
rect 2859 25939 2915 25995
rect 3001 25939 3057 25995
rect 3143 25939 3199 25995
rect 3285 25939 3341 25995
rect 3427 25939 3483 25995
rect 3569 25939 3625 25995
rect 3711 25939 3767 25995
rect 3853 25939 3909 25995
rect 3995 25939 4051 25995
rect 4137 25939 4193 25995
rect 4279 25939 4335 25995
rect 4421 25939 4477 25995
rect 4563 25939 4619 25995
rect 4705 25939 4761 25995
rect 4847 25939 4903 25995
rect 4989 25939 5045 25995
rect 5131 25939 5187 25995
rect 5273 25939 5329 25995
rect 5415 25939 5471 25995
rect 5557 25939 5613 25995
rect 5699 25939 5755 25995
rect 5841 25939 5897 25995
rect 5983 25939 6039 25995
rect 6125 25939 6181 25995
rect 6267 25939 6323 25995
rect 6409 25939 6465 25995
rect 6551 25939 6607 25995
rect 6693 25939 6749 25995
rect 6835 25939 6891 25995
rect 6977 25939 7033 25995
rect 7119 25939 7175 25995
rect 7261 25939 7317 25995
rect 7403 25939 7459 25995
rect 7545 25939 7601 25995
rect 7687 25939 7743 25995
rect 7829 25939 7885 25995
rect 7971 25939 8027 25995
rect 8113 25939 8169 25995
rect 8255 25939 8311 25995
rect 8397 25939 8453 25995
rect 8539 25939 8595 25995
rect 8681 25939 8737 25995
rect 8823 25939 8879 25995
rect 8965 25939 9021 25995
rect 9107 25939 9163 25995
rect 9249 25939 9305 25995
rect 9391 25939 9447 25995
rect 9533 25939 9589 25995
rect 9675 25939 9731 25995
rect 9817 25939 9873 25995
rect 9959 25939 10015 25995
rect 10101 25939 10157 25995
rect 10243 25939 10299 25995
rect 10385 25939 10441 25995
rect 10527 25939 10583 25995
rect 10669 25939 10725 25995
rect 10811 25939 10867 25995
rect 10953 25939 11009 25995
rect 11095 25939 11151 25995
rect 11237 25939 11293 25995
rect 11379 25939 11435 25995
rect 11521 25939 11577 25995
rect 11663 25939 11719 25995
rect 11805 25939 11861 25995
rect 11947 25939 12003 25995
rect 12089 25939 12145 25995
rect 12231 25939 12287 25995
rect 12373 25939 12429 25995
rect 12515 25939 12571 25995
rect 12657 25939 12713 25995
rect 12799 25939 12855 25995
rect 12941 25939 12997 25995
rect 13083 25939 13139 25995
rect 13225 25939 13281 25995
rect 13367 25939 13423 25995
rect 13509 25939 13565 25995
rect 13651 25939 13707 25995
rect 13793 25939 13849 25995
rect 13935 25939 13991 25995
rect 14077 25939 14133 25995
rect 14219 25939 14275 25995
rect 14361 25939 14417 25995
rect 14503 25939 14559 25995
rect 14645 25939 14701 25995
rect 14787 25939 14843 25995
rect 161 25797 217 25853
rect 303 25797 359 25853
rect 445 25797 501 25853
rect 587 25797 643 25853
rect 729 25797 785 25853
rect 871 25797 927 25853
rect 1013 25797 1069 25853
rect 1155 25797 1211 25853
rect 1297 25797 1353 25853
rect 1439 25797 1495 25853
rect 1581 25797 1637 25853
rect 1723 25797 1779 25853
rect 1865 25797 1921 25853
rect 2007 25797 2063 25853
rect 2149 25797 2205 25853
rect 2291 25797 2347 25853
rect 2433 25797 2489 25853
rect 2575 25797 2631 25853
rect 2717 25797 2773 25853
rect 2859 25797 2915 25853
rect 3001 25797 3057 25853
rect 3143 25797 3199 25853
rect 3285 25797 3341 25853
rect 3427 25797 3483 25853
rect 3569 25797 3625 25853
rect 3711 25797 3767 25853
rect 3853 25797 3909 25853
rect 3995 25797 4051 25853
rect 4137 25797 4193 25853
rect 4279 25797 4335 25853
rect 4421 25797 4477 25853
rect 4563 25797 4619 25853
rect 4705 25797 4761 25853
rect 4847 25797 4903 25853
rect 4989 25797 5045 25853
rect 5131 25797 5187 25853
rect 5273 25797 5329 25853
rect 5415 25797 5471 25853
rect 5557 25797 5613 25853
rect 5699 25797 5755 25853
rect 5841 25797 5897 25853
rect 5983 25797 6039 25853
rect 6125 25797 6181 25853
rect 6267 25797 6323 25853
rect 6409 25797 6465 25853
rect 6551 25797 6607 25853
rect 6693 25797 6749 25853
rect 6835 25797 6891 25853
rect 6977 25797 7033 25853
rect 7119 25797 7175 25853
rect 7261 25797 7317 25853
rect 7403 25797 7459 25853
rect 7545 25797 7601 25853
rect 7687 25797 7743 25853
rect 7829 25797 7885 25853
rect 7971 25797 8027 25853
rect 8113 25797 8169 25853
rect 8255 25797 8311 25853
rect 8397 25797 8453 25853
rect 8539 25797 8595 25853
rect 8681 25797 8737 25853
rect 8823 25797 8879 25853
rect 8965 25797 9021 25853
rect 9107 25797 9163 25853
rect 9249 25797 9305 25853
rect 9391 25797 9447 25853
rect 9533 25797 9589 25853
rect 9675 25797 9731 25853
rect 9817 25797 9873 25853
rect 9959 25797 10015 25853
rect 10101 25797 10157 25853
rect 10243 25797 10299 25853
rect 10385 25797 10441 25853
rect 10527 25797 10583 25853
rect 10669 25797 10725 25853
rect 10811 25797 10867 25853
rect 10953 25797 11009 25853
rect 11095 25797 11151 25853
rect 11237 25797 11293 25853
rect 11379 25797 11435 25853
rect 11521 25797 11577 25853
rect 11663 25797 11719 25853
rect 11805 25797 11861 25853
rect 11947 25797 12003 25853
rect 12089 25797 12145 25853
rect 12231 25797 12287 25853
rect 12373 25797 12429 25853
rect 12515 25797 12571 25853
rect 12657 25797 12713 25853
rect 12799 25797 12855 25853
rect 12941 25797 12997 25853
rect 13083 25797 13139 25853
rect 13225 25797 13281 25853
rect 13367 25797 13423 25853
rect 13509 25797 13565 25853
rect 13651 25797 13707 25853
rect 13793 25797 13849 25853
rect 13935 25797 13991 25853
rect 14077 25797 14133 25853
rect 14219 25797 14275 25853
rect 14361 25797 14417 25853
rect 14503 25797 14559 25853
rect 14645 25797 14701 25853
rect 14787 25797 14843 25853
rect 161 25655 217 25711
rect 303 25655 359 25711
rect 445 25655 501 25711
rect 587 25655 643 25711
rect 729 25655 785 25711
rect 871 25655 927 25711
rect 1013 25655 1069 25711
rect 1155 25655 1211 25711
rect 1297 25655 1353 25711
rect 1439 25655 1495 25711
rect 1581 25655 1637 25711
rect 1723 25655 1779 25711
rect 1865 25655 1921 25711
rect 2007 25655 2063 25711
rect 2149 25655 2205 25711
rect 2291 25655 2347 25711
rect 2433 25655 2489 25711
rect 2575 25655 2631 25711
rect 2717 25655 2773 25711
rect 2859 25655 2915 25711
rect 3001 25655 3057 25711
rect 3143 25655 3199 25711
rect 3285 25655 3341 25711
rect 3427 25655 3483 25711
rect 3569 25655 3625 25711
rect 3711 25655 3767 25711
rect 3853 25655 3909 25711
rect 3995 25655 4051 25711
rect 4137 25655 4193 25711
rect 4279 25655 4335 25711
rect 4421 25655 4477 25711
rect 4563 25655 4619 25711
rect 4705 25655 4761 25711
rect 4847 25655 4903 25711
rect 4989 25655 5045 25711
rect 5131 25655 5187 25711
rect 5273 25655 5329 25711
rect 5415 25655 5471 25711
rect 5557 25655 5613 25711
rect 5699 25655 5755 25711
rect 5841 25655 5897 25711
rect 5983 25655 6039 25711
rect 6125 25655 6181 25711
rect 6267 25655 6323 25711
rect 6409 25655 6465 25711
rect 6551 25655 6607 25711
rect 6693 25655 6749 25711
rect 6835 25655 6891 25711
rect 6977 25655 7033 25711
rect 7119 25655 7175 25711
rect 7261 25655 7317 25711
rect 7403 25655 7459 25711
rect 7545 25655 7601 25711
rect 7687 25655 7743 25711
rect 7829 25655 7885 25711
rect 7971 25655 8027 25711
rect 8113 25655 8169 25711
rect 8255 25655 8311 25711
rect 8397 25655 8453 25711
rect 8539 25655 8595 25711
rect 8681 25655 8737 25711
rect 8823 25655 8879 25711
rect 8965 25655 9021 25711
rect 9107 25655 9163 25711
rect 9249 25655 9305 25711
rect 9391 25655 9447 25711
rect 9533 25655 9589 25711
rect 9675 25655 9731 25711
rect 9817 25655 9873 25711
rect 9959 25655 10015 25711
rect 10101 25655 10157 25711
rect 10243 25655 10299 25711
rect 10385 25655 10441 25711
rect 10527 25655 10583 25711
rect 10669 25655 10725 25711
rect 10811 25655 10867 25711
rect 10953 25655 11009 25711
rect 11095 25655 11151 25711
rect 11237 25655 11293 25711
rect 11379 25655 11435 25711
rect 11521 25655 11577 25711
rect 11663 25655 11719 25711
rect 11805 25655 11861 25711
rect 11947 25655 12003 25711
rect 12089 25655 12145 25711
rect 12231 25655 12287 25711
rect 12373 25655 12429 25711
rect 12515 25655 12571 25711
rect 12657 25655 12713 25711
rect 12799 25655 12855 25711
rect 12941 25655 12997 25711
rect 13083 25655 13139 25711
rect 13225 25655 13281 25711
rect 13367 25655 13423 25711
rect 13509 25655 13565 25711
rect 13651 25655 13707 25711
rect 13793 25655 13849 25711
rect 13935 25655 13991 25711
rect 14077 25655 14133 25711
rect 14219 25655 14275 25711
rect 14361 25655 14417 25711
rect 14503 25655 14559 25711
rect 14645 25655 14701 25711
rect 14787 25655 14843 25711
rect 161 25513 217 25569
rect 303 25513 359 25569
rect 445 25513 501 25569
rect 587 25513 643 25569
rect 729 25513 785 25569
rect 871 25513 927 25569
rect 1013 25513 1069 25569
rect 1155 25513 1211 25569
rect 1297 25513 1353 25569
rect 1439 25513 1495 25569
rect 1581 25513 1637 25569
rect 1723 25513 1779 25569
rect 1865 25513 1921 25569
rect 2007 25513 2063 25569
rect 2149 25513 2205 25569
rect 2291 25513 2347 25569
rect 2433 25513 2489 25569
rect 2575 25513 2631 25569
rect 2717 25513 2773 25569
rect 2859 25513 2915 25569
rect 3001 25513 3057 25569
rect 3143 25513 3199 25569
rect 3285 25513 3341 25569
rect 3427 25513 3483 25569
rect 3569 25513 3625 25569
rect 3711 25513 3767 25569
rect 3853 25513 3909 25569
rect 3995 25513 4051 25569
rect 4137 25513 4193 25569
rect 4279 25513 4335 25569
rect 4421 25513 4477 25569
rect 4563 25513 4619 25569
rect 4705 25513 4761 25569
rect 4847 25513 4903 25569
rect 4989 25513 5045 25569
rect 5131 25513 5187 25569
rect 5273 25513 5329 25569
rect 5415 25513 5471 25569
rect 5557 25513 5613 25569
rect 5699 25513 5755 25569
rect 5841 25513 5897 25569
rect 5983 25513 6039 25569
rect 6125 25513 6181 25569
rect 6267 25513 6323 25569
rect 6409 25513 6465 25569
rect 6551 25513 6607 25569
rect 6693 25513 6749 25569
rect 6835 25513 6891 25569
rect 6977 25513 7033 25569
rect 7119 25513 7175 25569
rect 7261 25513 7317 25569
rect 7403 25513 7459 25569
rect 7545 25513 7601 25569
rect 7687 25513 7743 25569
rect 7829 25513 7885 25569
rect 7971 25513 8027 25569
rect 8113 25513 8169 25569
rect 8255 25513 8311 25569
rect 8397 25513 8453 25569
rect 8539 25513 8595 25569
rect 8681 25513 8737 25569
rect 8823 25513 8879 25569
rect 8965 25513 9021 25569
rect 9107 25513 9163 25569
rect 9249 25513 9305 25569
rect 9391 25513 9447 25569
rect 9533 25513 9589 25569
rect 9675 25513 9731 25569
rect 9817 25513 9873 25569
rect 9959 25513 10015 25569
rect 10101 25513 10157 25569
rect 10243 25513 10299 25569
rect 10385 25513 10441 25569
rect 10527 25513 10583 25569
rect 10669 25513 10725 25569
rect 10811 25513 10867 25569
rect 10953 25513 11009 25569
rect 11095 25513 11151 25569
rect 11237 25513 11293 25569
rect 11379 25513 11435 25569
rect 11521 25513 11577 25569
rect 11663 25513 11719 25569
rect 11805 25513 11861 25569
rect 11947 25513 12003 25569
rect 12089 25513 12145 25569
rect 12231 25513 12287 25569
rect 12373 25513 12429 25569
rect 12515 25513 12571 25569
rect 12657 25513 12713 25569
rect 12799 25513 12855 25569
rect 12941 25513 12997 25569
rect 13083 25513 13139 25569
rect 13225 25513 13281 25569
rect 13367 25513 13423 25569
rect 13509 25513 13565 25569
rect 13651 25513 13707 25569
rect 13793 25513 13849 25569
rect 13935 25513 13991 25569
rect 14077 25513 14133 25569
rect 14219 25513 14275 25569
rect 14361 25513 14417 25569
rect 14503 25513 14559 25569
rect 14645 25513 14701 25569
rect 14787 25513 14843 25569
rect 161 25371 217 25427
rect 303 25371 359 25427
rect 445 25371 501 25427
rect 587 25371 643 25427
rect 729 25371 785 25427
rect 871 25371 927 25427
rect 1013 25371 1069 25427
rect 1155 25371 1211 25427
rect 1297 25371 1353 25427
rect 1439 25371 1495 25427
rect 1581 25371 1637 25427
rect 1723 25371 1779 25427
rect 1865 25371 1921 25427
rect 2007 25371 2063 25427
rect 2149 25371 2205 25427
rect 2291 25371 2347 25427
rect 2433 25371 2489 25427
rect 2575 25371 2631 25427
rect 2717 25371 2773 25427
rect 2859 25371 2915 25427
rect 3001 25371 3057 25427
rect 3143 25371 3199 25427
rect 3285 25371 3341 25427
rect 3427 25371 3483 25427
rect 3569 25371 3625 25427
rect 3711 25371 3767 25427
rect 3853 25371 3909 25427
rect 3995 25371 4051 25427
rect 4137 25371 4193 25427
rect 4279 25371 4335 25427
rect 4421 25371 4477 25427
rect 4563 25371 4619 25427
rect 4705 25371 4761 25427
rect 4847 25371 4903 25427
rect 4989 25371 5045 25427
rect 5131 25371 5187 25427
rect 5273 25371 5329 25427
rect 5415 25371 5471 25427
rect 5557 25371 5613 25427
rect 5699 25371 5755 25427
rect 5841 25371 5897 25427
rect 5983 25371 6039 25427
rect 6125 25371 6181 25427
rect 6267 25371 6323 25427
rect 6409 25371 6465 25427
rect 6551 25371 6607 25427
rect 6693 25371 6749 25427
rect 6835 25371 6891 25427
rect 6977 25371 7033 25427
rect 7119 25371 7175 25427
rect 7261 25371 7317 25427
rect 7403 25371 7459 25427
rect 7545 25371 7601 25427
rect 7687 25371 7743 25427
rect 7829 25371 7885 25427
rect 7971 25371 8027 25427
rect 8113 25371 8169 25427
rect 8255 25371 8311 25427
rect 8397 25371 8453 25427
rect 8539 25371 8595 25427
rect 8681 25371 8737 25427
rect 8823 25371 8879 25427
rect 8965 25371 9021 25427
rect 9107 25371 9163 25427
rect 9249 25371 9305 25427
rect 9391 25371 9447 25427
rect 9533 25371 9589 25427
rect 9675 25371 9731 25427
rect 9817 25371 9873 25427
rect 9959 25371 10015 25427
rect 10101 25371 10157 25427
rect 10243 25371 10299 25427
rect 10385 25371 10441 25427
rect 10527 25371 10583 25427
rect 10669 25371 10725 25427
rect 10811 25371 10867 25427
rect 10953 25371 11009 25427
rect 11095 25371 11151 25427
rect 11237 25371 11293 25427
rect 11379 25371 11435 25427
rect 11521 25371 11577 25427
rect 11663 25371 11719 25427
rect 11805 25371 11861 25427
rect 11947 25371 12003 25427
rect 12089 25371 12145 25427
rect 12231 25371 12287 25427
rect 12373 25371 12429 25427
rect 12515 25371 12571 25427
rect 12657 25371 12713 25427
rect 12799 25371 12855 25427
rect 12941 25371 12997 25427
rect 13083 25371 13139 25427
rect 13225 25371 13281 25427
rect 13367 25371 13423 25427
rect 13509 25371 13565 25427
rect 13651 25371 13707 25427
rect 13793 25371 13849 25427
rect 13935 25371 13991 25427
rect 14077 25371 14133 25427
rect 14219 25371 14275 25427
rect 14361 25371 14417 25427
rect 14503 25371 14559 25427
rect 14645 25371 14701 25427
rect 14787 25371 14843 25427
rect 161 25229 217 25285
rect 303 25229 359 25285
rect 445 25229 501 25285
rect 587 25229 643 25285
rect 729 25229 785 25285
rect 871 25229 927 25285
rect 1013 25229 1069 25285
rect 1155 25229 1211 25285
rect 1297 25229 1353 25285
rect 1439 25229 1495 25285
rect 1581 25229 1637 25285
rect 1723 25229 1779 25285
rect 1865 25229 1921 25285
rect 2007 25229 2063 25285
rect 2149 25229 2205 25285
rect 2291 25229 2347 25285
rect 2433 25229 2489 25285
rect 2575 25229 2631 25285
rect 2717 25229 2773 25285
rect 2859 25229 2915 25285
rect 3001 25229 3057 25285
rect 3143 25229 3199 25285
rect 3285 25229 3341 25285
rect 3427 25229 3483 25285
rect 3569 25229 3625 25285
rect 3711 25229 3767 25285
rect 3853 25229 3909 25285
rect 3995 25229 4051 25285
rect 4137 25229 4193 25285
rect 4279 25229 4335 25285
rect 4421 25229 4477 25285
rect 4563 25229 4619 25285
rect 4705 25229 4761 25285
rect 4847 25229 4903 25285
rect 4989 25229 5045 25285
rect 5131 25229 5187 25285
rect 5273 25229 5329 25285
rect 5415 25229 5471 25285
rect 5557 25229 5613 25285
rect 5699 25229 5755 25285
rect 5841 25229 5897 25285
rect 5983 25229 6039 25285
rect 6125 25229 6181 25285
rect 6267 25229 6323 25285
rect 6409 25229 6465 25285
rect 6551 25229 6607 25285
rect 6693 25229 6749 25285
rect 6835 25229 6891 25285
rect 6977 25229 7033 25285
rect 7119 25229 7175 25285
rect 7261 25229 7317 25285
rect 7403 25229 7459 25285
rect 7545 25229 7601 25285
rect 7687 25229 7743 25285
rect 7829 25229 7885 25285
rect 7971 25229 8027 25285
rect 8113 25229 8169 25285
rect 8255 25229 8311 25285
rect 8397 25229 8453 25285
rect 8539 25229 8595 25285
rect 8681 25229 8737 25285
rect 8823 25229 8879 25285
rect 8965 25229 9021 25285
rect 9107 25229 9163 25285
rect 9249 25229 9305 25285
rect 9391 25229 9447 25285
rect 9533 25229 9589 25285
rect 9675 25229 9731 25285
rect 9817 25229 9873 25285
rect 9959 25229 10015 25285
rect 10101 25229 10157 25285
rect 10243 25229 10299 25285
rect 10385 25229 10441 25285
rect 10527 25229 10583 25285
rect 10669 25229 10725 25285
rect 10811 25229 10867 25285
rect 10953 25229 11009 25285
rect 11095 25229 11151 25285
rect 11237 25229 11293 25285
rect 11379 25229 11435 25285
rect 11521 25229 11577 25285
rect 11663 25229 11719 25285
rect 11805 25229 11861 25285
rect 11947 25229 12003 25285
rect 12089 25229 12145 25285
rect 12231 25229 12287 25285
rect 12373 25229 12429 25285
rect 12515 25229 12571 25285
rect 12657 25229 12713 25285
rect 12799 25229 12855 25285
rect 12941 25229 12997 25285
rect 13083 25229 13139 25285
rect 13225 25229 13281 25285
rect 13367 25229 13423 25285
rect 13509 25229 13565 25285
rect 13651 25229 13707 25285
rect 13793 25229 13849 25285
rect 13935 25229 13991 25285
rect 14077 25229 14133 25285
rect 14219 25229 14275 25285
rect 14361 25229 14417 25285
rect 14503 25229 14559 25285
rect 14645 25229 14701 25285
rect 14787 25229 14843 25285
rect 161 24907 217 24963
rect 303 24907 359 24963
rect 445 24907 501 24963
rect 587 24907 643 24963
rect 729 24907 785 24963
rect 871 24907 927 24963
rect 1013 24907 1069 24963
rect 1155 24907 1211 24963
rect 1297 24907 1353 24963
rect 1439 24907 1495 24963
rect 1581 24907 1637 24963
rect 1723 24907 1779 24963
rect 1865 24907 1921 24963
rect 2007 24907 2063 24963
rect 2149 24907 2205 24963
rect 2291 24907 2347 24963
rect 2433 24907 2489 24963
rect 2575 24907 2631 24963
rect 2717 24907 2773 24963
rect 2859 24907 2915 24963
rect 3001 24907 3057 24963
rect 3143 24907 3199 24963
rect 3285 24907 3341 24963
rect 3427 24907 3483 24963
rect 3569 24907 3625 24963
rect 3711 24907 3767 24963
rect 3853 24907 3909 24963
rect 3995 24907 4051 24963
rect 4137 24907 4193 24963
rect 4279 24907 4335 24963
rect 4421 24907 4477 24963
rect 4563 24907 4619 24963
rect 4705 24907 4761 24963
rect 4847 24907 4903 24963
rect 4989 24907 5045 24963
rect 5131 24907 5187 24963
rect 5273 24907 5329 24963
rect 5415 24907 5471 24963
rect 5557 24907 5613 24963
rect 5699 24907 5755 24963
rect 5841 24907 5897 24963
rect 5983 24907 6039 24963
rect 6125 24907 6181 24963
rect 6267 24907 6323 24963
rect 6409 24907 6465 24963
rect 6551 24907 6607 24963
rect 6693 24907 6749 24963
rect 6835 24907 6891 24963
rect 6977 24907 7033 24963
rect 7119 24907 7175 24963
rect 7261 24907 7317 24963
rect 7403 24907 7459 24963
rect 7545 24907 7601 24963
rect 7687 24907 7743 24963
rect 7829 24907 7885 24963
rect 7971 24907 8027 24963
rect 8113 24907 8169 24963
rect 8255 24907 8311 24963
rect 8397 24907 8453 24963
rect 8539 24907 8595 24963
rect 8681 24907 8737 24963
rect 8823 24907 8879 24963
rect 8965 24907 9021 24963
rect 9107 24907 9163 24963
rect 9249 24907 9305 24963
rect 9391 24907 9447 24963
rect 9533 24907 9589 24963
rect 9675 24907 9731 24963
rect 9817 24907 9873 24963
rect 9959 24907 10015 24963
rect 10101 24907 10157 24963
rect 10243 24907 10299 24963
rect 10385 24907 10441 24963
rect 10527 24907 10583 24963
rect 10669 24907 10725 24963
rect 10811 24907 10867 24963
rect 10953 24907 11009 24963
rect 11095 24907 11151 24963
rect 11237 24907 11293 24963
rect 11379 24907 11435 24963
rect 11521 24907 11577 24963
rect 11663 24907 11719 24963
rect 11805 24907 11861 24963
rect 11947 24907 12003 24963
rect 12089 24907 12145 24963
rect 12231 24907 12287 24963
rect 12373 24907 12429 24963
rect 12515 24907 12571 24963
rect 12657 24907 12713 24963
rect 12799 24907 12855 24963
rect 12941 24907 12997 24963
rect 13083 24907 13139 24963
rect 13225 24907 13281 24963
rect 13367 24907 13423 24963
rect 13509 24907 13565 24963
rect 13651 24907 13707 24963
rect 13793 24907 13849 24963
rect 13935 24907 13991 24963
rect 14077 24907 14133 24963
rect 14219 24907 14275 24963
rect 14361 24907 14417 24963
rect 14503 24907 14559 24963
rect 14645 24907 14701 24963
rect 14787 24907 14843 24963
rect 161 24765 217 24821
rect 303 24765 359 24821
rect 445 24765 501 24821
rect 587 24765 643 24821
rect 729 24765 785 24821
rect 871 24765 927 24821
rect 1013 24765 1069 24821
rect 1155 24765 1211 24821
rect 1297 24765 1353 24821
rect 1439 24765 1495 24821
rect 1581 24765 1637 24821
rect 1723 24765 1779 24821
rect 1865 24765 1921 24821
rect 2007 24765 2063 24821
rect 2149 24765 2205 24821
rect 2291 24765 2347 24821
rect 2433 24765 2489 24821
rect 2575 24765 2631 24821
rect 2717 24765 2773 24821
rect 2859 24765 2915 24821
rect 3001 24765 3057 24821
rect 3143 24765 3199 24821
rect 3285 24765 3341 24821
rect 3427 24765 3483 24821
rect 3569 24765 3625 24821
rect 3711 24765 3767 24821
rect 3853 24765 3909 24821
rect 3995 24765 4051 24821
rect 4137 24765 4193 24821
rect 4279 24765 4335 24821
rect 4421 24765 4477 24821
rect 4563 24765 4619 24821
rect 4705 24765 4761 24821
rect 4847 24765 4903 24821
rect 4989 24765 5045 24821
rect 5131 24765 5187 24821
rect 5273 24765 5329 24821
rect 5415 24765 5471 24821
rect 5557 24765 5613 24821
rect 5699 24765 5755 24821
rect 5841 24765 5897 24821
rect 5983 24765 6039 24821
rect 6125 24765 6181 24821
rect 6267 24765 6323 24821
rect 6409 24765 6465 24821
rect 6551 24765 6607 24821
rect 6693 24765 6749 24821
rect 6835 24765 6891 24821
rect 6977 24765 7033 24821
rect 7119 24765 7175 24821
rect 7261 24765 7317 24821
rect 7403 24765 7459 24821
rect 7545 24765 7601 24821
rect 7687 24765 7743 24821
rect 7829 24765 7885 24821
rect 7971 24765 8027 24821
rect 8113 24765 8169 24821
rect 8255 24765 8311 24821
rect 8397 24765 8453 24821
rect 8539 24765 8595 24821
rect 8681 24765 8737 24821
rect 8823 24765 8879 24821
rect 8965 24765 9021 24821
rect 9107 24765 9163 24821
rect 9249 24765 9305 24821
rect 9391 24765 9447 24821
rect 9533 24765 9589 24821
rect 9675 24765 9731 24821
rect 9817 24765 9873 24821
rect 9959 24765 10015 24821
rect 10101 24765 10157 24821
rect 10243 24765 10299 24821
rect 10385 24765 10441 24821
rect 10527 24765 10583 24821
rect 10669 24765 10725 24821
rect 10811 24765 10867 24821
rect 10953 24765 11009 24821
rect 11095 24765 11151 24821
rect 11237 24765 11293 24821
rect 11379 24765 11435 24821
rect 11521 24765 11577 24821
rect 11663 24765 11719 24821
rect 11805 24765 11861 24821
rect 11947 24765 12003 24821
rect 12089 24765 12145 24821
rect 12231 24765 12287 24821
rect 12373 24765 12429 24821
rect 12515 24765 12571 24821
rect 12657 24765 12713 24821
rect 12799 24765 12855 24821
rect 12941 24765 12997 24821
rect 13083 24765 13139 24821
rect 13225 24765 13281 24821
rect 13367 24765 13423 24821
rect 13509 24765 13565 24821
rect 13651 24765 13707 24821
rect 13793 24765 13849 24821
rect 13935 24765 13991 24821
rect 14077 24765 14133 24821
rect 14219 24765 14275 24821
rect 14361 24765 14417 24821
rect 14503 24765 14559 24821
rect 14645 24765 14701 24821
rect 14787 24765 14843 24821
rect 161 24623 217 24679
rect 303 24623 359 24679
rect 445 24623 501 24679
rect 587 24623 643 24679
rect 729 24623 785 24679
rect 871 24623 927 24679
rect 1013 24623 1069 24679
rect 1155 24623 1211 24679
rect 1297 24623 1353 24679
rect 1439 24623 1495 24679
rect 1581 24623 1637 24679
rect 1723 24623 1779 24679
rect 1865 24623 1921 24679
rect 2007 24623 2063 24679
rect 2149 24623 2205 24679
rect 2291 24623 2347 24679
rect 2433 24623 2489 24679
rect 2575 24623 2631 24679
rect 2717 24623 2773 24679
rect 2859 24623 2915 24679
rect 3001 24623 3057 24679
rect 3143 24623 3199 24679
rect 3285 24623 3341 24679
rect 3427 24623 3483 24679
rect 3569 24623 3625 24679
rect 3711 24623 3767 24679
rect 3853 24623 3909 24679
rect 3995 24623 4051 24679
rect 4137 24623 4193 24679
rect 4279 24623 4335 24679
rect 4421 24623 4477 24679
rect 4563 24623 4619 24679
rect 4705 24623 4761 24679
rect 4847 24623 4903 24679
rect 4989 24623 5045 24679
rect 5131 24623 5187 24679
rect 5273 24623 5329 24679
rect 5415 24623 5471 24679
rect 5557 24623 5613 24679
rect 5699 24623 5755 24679
rect 5841 24623 5897 24679
rect 5983 24623 6039 24679
rect 6125 24623 6181 24679
rect 6267 24623 6323 24679
rect 6409 24623 6465 24679
rect 6551 24623 6607 24679
rect 6693 24623 6749 24679
rect 6835 24623 6891 24679
rect 6977 24623 7033 24679
rect 7119 24623 7175 24679
rect 7261 24623 7317 24679
rect 7403 24623 7459 24679
rect 7545 24623 7601 24679
rect 7687 24623 7743 24679
rect 7829 24623 7885 24679
rect 7971 24623 8027 24679
rect 8113 24623 8169 24679
rect 8255 24623 8311 24679
rect 8397 24623 8453 24679
rect 8539 24623 8595 24679
rect 8681 24623 8737 24679
rect 8823 24623 8879 24679
rect 8965 24623 9021 24679
rect 9107 24623 9163 24679
rect 9249 24623 9305 24679
rect 9391 24623 9447 24679
rect 9533 24623 9589 24679
rect 9675 24623 9731 24679
rect 9817 24623 9873 24679
rect 9959 24623 10015 24679
rect 10101 24623 10157 24679
rect 10243 24623 10299 24679
rect 10385 24623 10441 24679
rect 10527 24623 10583 24679
rect 10669 24623 10725 24679
rect 10811 24623 10867 24679
rect 10953 24623 11009 24679
rect 11095 24623 11151 24679
rect 11237 24623 11293 24679
rect 11379 24623 11435 24679
rect 11521 24623 11577 24679
rect 11663 24623 11719 24679
rect 11805 24623 11861 24679
rect 11947 24623 12003 24679
rect 12089 24623 12145 24679
rect 12231 24623 12287 24679
rect 12373 24623 12429 24679
rect 12515 24623 12571 24679
rect 12657 24623 12713 24679
rect 12799 24623 12855 24679
rect 12941 24623 12997 24679
rect 13083 24623 13139 24679
rect 13225 24623 13281 24679
rect 13367 24623 13423 24679
rect 13509 24623 13565 24679
rect 13651 24623 13707 24679
rect 13793 24623 13849 24679
rect 13935 24623 13991 24679
rect 14077 24623 14133 24679
rect 14219 24623 14275 24679
rect 14361 24623 14417 24679
rect 14503 24623 14559 24679
rect 14645 24623 14701 24679
rect 14787 24623 14843 24679
rect 161 24481 217 24537
rect 303 24481 359 24537
rect 445 24481 501 24537
rect 587 24481 643 24537
rect 729 24481 785 24537
rect 871 24481 927 24537
rect 1013 24481 1069 24537
rect 1155 24481 1211 24537
rect 1297 24481 1353 24537
rect 1439 24481 1495 24537
rect 1581 24481 1637 24537
rect 1723 24481 1779 24537
rect 1865 24481 1921 24537
rect 2007 24481 2063 24537
rect 2149 24481 2205 24537
rect 2291 24481 2347 24537
rect 2433 24481 2489 24537
rect 2575 24481 2631 24537
rect 2717 24481 2773 24537
rect 2859 24481 2915 24537
rect 3001 24481 3057 24537
rect 3143 24481 3199 24537
rect 3285 24481 3341 24537
rect 3427 24481 3483 24537
rect 3569 24481 3625 24537
rect 3711 24481 3767 24537
rect 3853 24481 3909 24537
rect 3995 24481 4051 24537
rect 4137 24481 4193 24537
rect 4279 24481 4335 24537
rect 4421 24481 4477 24537
rect 4563 24481 4619 24537
rect 4705 24481 4761 24537
rect 4847 24481 4903 24537
rect 4989 24481 5045 24537
rect 5131 24481 5187 24537
rect 5273 24481 5329 24537
rect 5415 24481 5471 24537
rect 5557 24481 5613 24537
rect 5699 24481 5755 24537
rect 5841 24481 5897 24537
rect 5983 24481 6039 24537
rect 6125 24481 6181 24537
rect 6267 24481 6323 24537
rect 6409 24481 6465 24537
rect 6551 24481 6607 24537
rect 6693 24481 6749 24537
rect 6835 24481 6891 24537
rect 6977 24481 7033 24537
rect 7119 24481 7175 24537
rect 7261 24481 7317 24537
rect 7403 24481 7459 24537
rect 7545 24481 7601 24537
rect 7687 24481 7743 24537
rect 7829 24481 7885 24537
rect 7971 24481 8027 24537
rect 8113 24481 8169 24537
rect 8255 24481 8311 24537
rect 8397 24481 8453 24537
rect 8539 24481 8595 24537
rect 8681 24481 8737 24537
rect 8823 24481 8879 24537
rect 8965 24481 9021 24537
rect 9107 24481 9163 24537
rect 9249 24481 9305 24537
rect 9391 24481 9447 24537
rect 9533 24481 9589 24537
rect 9675 24481 9731 24537
rect 9817 24481 9873 24537
rect 9959 24481 10015 24537
rect 10101 24481 10157 24537
rect 10243 24481 10299 24537
rect 10385 24481 10441 24537
rect 10527 24481 10583 24537
rect 10669 24481 10725 24537
rect 10811 24481 10867 24537
rect 10953 24481 11009 24537
rect 11095 24481 11151 24537
rect 11237 24481 11293 24537
rect 11379 24481 11435 24537
rect 11521 24481 11577 24537
rect 11663 24481 11719 24537
rect 11805 24481 11861 24537
rect 11947 24481 12003 24537
rect 12089 24481 12145 24537
rect 12231 24481 12287 24537
rect 12373 24481 12429 24537
rect 12515 24481 12571 24537
rect 12657 24481 12713 24537
rect 12799 24481 12855 24537
rect 12941 24481 12997 24537
rect 13083 24481 13139 24537
rect 13225 24481 13281 24537
rect 13367 24481 13423 24537
rect 13509 24481 13565 24537
rect 13651 24481 13707 24537
rect 13793 24481 13849 24537
rect 13935 24481 13991 24537
rect 14077 24481 14133 24537
rect 14219 24481 14275 24537
rect 14361 24481 14417 24537
rect 14503 24481 14559 24537
rect 14645 24481 14701 24537
rect 14787 24481 14843 24537
rect 161 24339 217 24395
rect 303 24339 359 24395
rect 445 24339 501 24395
rect 587 24339 643 24395
rect 729 24339 785 24395
rect 871 24339 927 24395
rect 1013 24339 1069 24395
rect 1155 24339 1211 24395
rect 1297 24339 1353 24395
rect 1439 24339 1495 24395
rect 1581 24339 1637 24395
rect 1723 24339 1779 24395
rect 1865 24339 1921 24395
rect 2007 24339 2063 24395
rect 2149 24339 2205 24395
rect 2291 24339 2347 24395
rect 2433 24339 2489 24395
rect 2575 24339 2631 24395
rect 2717 24339 2773 24395
rect 2859 24339 2915 24395
rect 3001 24339 3057 24395
rect 3143 24339 3199 24395
rect 3285 24339 3341 24395
rect 3427 24339 3483 24395
rect 3569 24339 3625 24395
rect 3711 24339 3767 24395
rect 3853 24339 3909 24395
rect 3995 24339 4051 24395
rect 4137 24339 4193 24395
rect 4279 24339 4335 24395
rect 4421 24339 4477 24395
rect 4563 24339 4619 24395
rect 4705 24339 4761 24395
rect 4847 24339 4903 24395
rect 4989 24339 5045 24395
rect 5131 24339 5187 24395
rect 5273 24339 5329 24395
rect 5415 24339 5471 24395
rect 5557 24339 5613 24395
rect 5699 24339 5755 24395
rect 5841 24339 5897 24395
rect 5983 24339 6039 24395
rect 6125 24339 6181 24395
rect 6267 24339 6323 24395
rect 6409 24339 6465 24395
rect 6551 24339 6607 24395
rect 6693 24339 6749 24395
rect 6835 24339 6891 24395
rect 6977 24339 7033 24395
rect 7119 24339 7175 24395
rect 7261 24339 7317 24395
rect 7403 24339 7459 24395
rect 7545 24339 7601 24395
rect 7687 24339 7743 24395
rect 7829 24339 7885 24395
rect 7971 24339 8027 24395
rect 8113 24339 8169 24395
rect 8255 24339 8311 24395
rect 8397 24339 8453 24395
rect 8539 24339 8595 24395
rect 8681 24339 8737 24395
rect 8823 24339 8879 24395
rect 8965 24339 9021 24395
rect 9107 24339 9163 24395
rect 9249 24339 9305 24395
rect 9391 24339 9447 24395
rect 9533 24339 9589 24395
rect 9675 24339 9731 24395
rect 9817 24339 9873 24395
rect 9959 24339 10015 24395
rect 10101 24339 10157 24395
rect 10243 24339 10299 24395
rect 10385 24339 10441 24395
rect 10527 24339 10583 24395
rect 10669 24339 10725 24395
rect 10811 24339 10867 24395
rect 10953 24339 11009 24395
rect 11095 24339 11151 24395
rect 11237 24339 11293 24395
rect 11379 24339 11435 24395
rect 11521 24339 11577 24395
rect 11663 24339 11719 24395
rect 11805 24339 11861 24395
rect 11947 24339 12003 24395
rect 12089 24339 12145 24395
rect 12231 24339 12287 24395
rect 12373 24339 12429 24395
rect 12515 24339 12571 24395
rect 12657 24339 12713 24395
rect 12799 24339 12855 24395
rect 12941 24339 12997 24395
rect 13083 24339 13139 24395
rect 13225 24339 13281 24395
rect 13367 24339 13423 24395
rect 13509 24339 13565 24395
rect 13651 24339 13707 24395
rect 13793 24339 13849 24395
rect 13935 24339 13991 24395
rect 14077 24339 14133 24395
rect 14219 24339 14275 24395
rect 14361 24339 14417 24395
rect 14503 24339 14559 24395
rect 14645 24339 14701 24395
rect 14787 24339 14843 24395
rect 161 24197 217 24253
rect 303 24197 359 24253
rect 445 24197 501 24253
rect 587 24197 643 24253
rect 729 24197 785 24253
rect 871 24197 927 24253
rect 1013 24197 1069 24253
rect 1155 24197 1211 24253
rect 1297 24197 1353 24253
rect 1439 24197 1495 24253
rect 1581 24197 1637 24253
rect 1723 24197 1779 24253
rect 1865 24197 1921 24253
rect 2007 24197 2063 24253
rect 2149 24197 2205 24253
rect 2291 24197 2347 24253
rect 2433 24197 2489 24253
rect 2575 24197 2631 24253
rect 2717 24197 2773 24253
rect 2859 24197 2915 24253
rect 3001 24197 3057 24253
rect 3143 24197 3199 24253
rect 3285 24197 3341 24253
rect 3427 24197 3483 24253
rect 3569 24197 3625 24253
rect 3711 24197 3767 24253
rect 3853 24197 3909 24253
rect 3995 24197 4051 24253
rect 4137 24197 4193 24253
rect 4279 24197 4335 24253
rect 4421 24197 4477 24253
rect 4563 24197 4619 24253
rect 4705 24197 4761 24253
rect 4847 24197 4903 24253
rect 4989 24197 5045 24253
rect 5131 24197 5187 24253
rect 5273 24197 5329 24253
rect 5415 24197 5471 24253
rect 5557 24197 5613 24253
rect 5699 24197 5755 24253
rect 5841 24197 5897 24253
rect 5983 24197 6039 24253
rect 6125 24197 6181 24253
rect 6267 24197 6323 24253
rect 6409 24197 6465 24253
rect 6551 24197 6607 24253
rect 6693 24197 6749 24253
rect 6835 24197 6891 24253
rect 6977 24197 7033 24253
rect 7119 24197 7175 24253
rect 7261 24197 7317 24253
rect 7403 24197 7459 24253
rect 7545 24197 7601 24253
rect 7687 24197 7743 24253
rect 7829 24197 7885 24253
rect 7971 24197 8027 24253
rect 8113 24197 8169 24253
rect 8255 24197 8311 24253
rect 8397 24197 8453 24253
rect 8539 24197 8595 24253
rect 8681 24197 8737 24253
rect 8823 24197 8879 24253
rect 8965 24197 9021 24253
rect 9107 24197 9163 24253
rect 9249 24197 9305 24253
rect 9391 24197 9447 24253
rect 9533 24197 9589 24253
rect 9675 24197 9731 24253
rect 9817 24197 9873 24253
rect 9959 24197 10015 24253
rect 10101 24197 10157 24253
rect 10243 24197 10299 24253
rect 10385 24197 10441 24253
rect 10527 24197 10583 24253
rect 10669 24197 10725 24253
rect 10811 24197 10867 24253
rect 10953 24197 11009 24253
rect 11095 24197 11151 24253
rect 11237 24197 11293 24253
rect 11379 24197 11435 24253
rect 11521 24197 11577 24253
rect 11663 24197 11719 24253
rect 11805 24197 11861 24253
rect 11947 24197 12003 24253
rect 12089 24197 12145 24253
rect 12231 24197 12287 24253
rect 12373 24197 12429 24253
rect 12515 24197 12571 24253
rect 12657 24197 12713 24253
rect 12799 24197 12855 24253
rect 12941 24197 12997 24253
rect 13083 24197 13139 24253
rect 13225 24197 13281 24253
rect 13367 24197 13423 24253
rect 13509 24197 13565 24253
rect 13651 24197 13707 24253
rect 13793 24197 13849 24253
rect 13935 24197 13991 24253
rect 14077 24197 14133 24253
rect 14219 24197 14275 24253
rect 14361 24197 14417 24253
rect 14503 24197 14559 24253
rect 14645 24197 14701 24253
rect 14787 24197 14843 24253
rect 161 24055 217 24111
rect 303 24055 359 24111
rect 445 24055 501 24111
rect 587 24055 643 24111
rect 729 24055 785 24111
rect 871 24055 927 24111
rect 1013 24055 1069 24111
rect 1155 24055 1211 24111
rect 1297 24055 1353 24111
rect 1439 24055 1495 24111
rect 1581 24055 1637 24111
rect 1723 24055 1779 24111
rect 1865 24055 1921 24111
rect 2007 24055 2063 24111
rect 2149 24055 2205 24111
rect 2291 24055 2347 24111
rect 2433 24055 2489 24111
rect 2575 24055 2631 24111
rect 2717 24055 2773 24111
rect 2859 24055 2915 24111
rect 3001 24055 3057 24111
rect 3143 24055 3199 24111
rect 3285 24055 3341 24111
rect 3427 24055 3483 24111
rect 3569 24055 3625 24111
rect 3711 24055 3767 24111
rect 3853 24055 3909 24111
rect 3995 24055 4051 24111
rect 4137 24055 4193 24111
rect 4279 24055 4335 24111
rect 4421 24055 4477 24111
rect 4563 24055 4619 24111
rect 4705 24055 4761 24111
rect 4847 24055 4903 24111
rect 4989 24055 5045 24111
rect 5131 24055 5187 24111
rect 5273 24055 5329 24111
rect 5415 24055 5471 24111
rect 5557 24055 5613 24111
rect 5699 24055 5755 24111
rect 5841 24055 5897 24111
rect 5983 24055 6039 24111
rect 6125 24055 6181 24111
rect 6267 24055 6323 24111
rect 6409 24055 6465 24111
rect 6551 24055 6607 24111
rect 6693 24055 6749 24111
rect 6835 24055 6891 24111
rect 6977 24055 7033 24111
rect 7119 24055 7175 24111
rect 7261 24055 7317 24111
rect 7403 24055 7459 24111
rect 7545 24055 7601 24111
rect 7687 24055 7743 24111
rect 7829 24055 7885 24111
rect 7971 24055 8027 24111
rect 8113 24055 8169 24111
rect 8255 24055 8311 24111
rect 8397 24055 8453 24111
rect 8539 24055 8595 24111
rect 8681 24055 8737 24111
rect 8823 24055 8879 24111
rect 8965 24055 9021 24111
rect 9107 24055 9163 24111
rect 9249 24055 9305 24111
rect 9391 24055 9447 24111
rect 9533 24055 9589 24111
rect 9675 24055 9731 24111
rect 9817 24055 9873 24111
rect 9959 24055 10015 24111
rect 10101 24055 10157 24111
rect 10243 24055 10299 24111
rect 10385 24055 10441 24111
rect 10527 24055 10583 24111
rect 10669 24055 10725 24111
rect 10811 24055 10867 24111
rect 10953 24055 11009 24111
rect 11095 24055 11151 24111
rect 11237 24055 11293 24111
rect 11379 24055 11435 24111
rect 11521 24055 11577 24111
rect 11663 24055 11719 24111
rect 11805 24055 11861 24111
rect 11947 24055 12003 24111
rect 12089 24055 12145 24111
rect 12231 24055 12287 24111
rect 12373 24055 12429 24111
rect 12515 24055 12571 24111
rect 12657 24055 12713 24111
rect 12799 24055 12855 24111
rect 12941 24055 12997 24111
rect 13083 24055 13139 24111
rect 13225 24055 13281 24111
rect 13367 24055 13423 24111
rect 13509 24055 13565 24111
rect 13651 24055 13707 24111
rect 13793 24055 13849 24111
rect 13935 24055 13991 24111
rect 14077 24055 14133 24111
rect 14219 24055 14275 24111
rect 14361 24055 14417 24111
rect 14503 24055 14559 24111
rect 14645 24055 14701 24111
rect 14787 24055 14843 24111
rect 161 23913 217 23969
rect 303 23913 359 23969
rect 445 23913 501 23969
rect 587 23913 643 23969
rect 729 23913 785 23969
rect 871 23913 927 23969
rect 1013 23913 1069 23969
rect 1155 23913 1211 23969
rect 1297 23913 1353 23969
rect 1439 23913 1495 23969
rect 1581 23913 1637 23969
rect 1723 23913 1779 23969
rect 1865 23913 1921 23969
rect 2007 23913 2063 23969
rect 2149 23913 2205 23969
rect 2291 23913 2347 23969
rect 2433 23913 2489 23969
rect 2575 23913 2631 23969
rect 2717 23913 2773 23969
rect 2859 23913 2915 23969
rect 3001 23913 3057 23969
rect 3143 23913 3199 23969
rect 3285 23913 3341 23969
rect 3427 23913 3483 23969
rect 3569 23913 3625 23969
rect 3711 23913 3767 23969
rect 3853 23913 3909 23969
rect 3995 23913 4051 23969
rect 4137 23913 4193 23969
rect 4279 23913 4335 23969
rect 4421 23913 4477 23969
rect 4563 23913 4619 23969
rect 4705 23913 4761 23969
rect 4847 23913 4903 23969
rect 4989 23913 5045 23969
rect 5131 23913 5187 23969
rect 5273 23913 5329 23969
rect 5415 23913 5471 23969
rect 5557 23913 5613 23969
rect 5699 23913 5755 23969
rect 5841 23913 5897 23969
rect 5983 23913 6039 23969
rect 6125 23913 6181 23969
rect 6267 23913 6323 23969
rect 6409 23913 6465 23969
rect 6551 23913 6607 23969
rect 6693 23913 6749 23969
rect 6835 23913 6891 23969
rect 6977 23913 7033 23969
rect 7119 23913 7175 23969
rect 7261 23913 7317 23969
rect 7403 23913 7459 23969
rect 7545 23913 7601 23969
rect 7687 23913 7743 23969
rect 7829 23913 7885 23969
rect 7971 23913 8027 23969
rect 8113 23913 8169 23969
rect 8255 23913 8311 23969
rect 8397 23913 8453 23969
rect 8539 23913 8595 23969
rect 8681 23913 8737 23969
rect 8823 23913 8879 23969
rect 8965 23913 9021 23969
rect 9107 23913 9163 23969
rect 9249 23913 9305 23969
rect 9391 23913 9447 23969
rect 9533 23913 9589 23969
rect 9675 23913 9731 23969
rect 9817 23913 9873 23969
rect 9959 23913 10015 23969
rect 10101 23913 10157 23969
rect 10243 23913 10299 23969
rect 10385 23913 10441 23969
rect 10527 23913 10583 23969
rect 10669 23913 10725 23969
rect 10811 23913 10867 23969
rect 10953 23913 11009 23969
rect 11095 23913 11151 23969
rect 11237 23913 11293 23969
rect 11379 23913 11435 23969
rect 11521 23913 11577 23969
rect 11663 23913 11719 23969
rect 11805 23913 11861 23969
rect 11947 23913 12003 23969
rect 12089 23913 12145 23969
rect 12231 23913 12287 23969
rect 12373 23913 12429 23969
rect 12515 23913 12571 23969
rect 12657 23913 12713 23969
rect 12799 23913 12855 23969
rect 12941 23913 12997 23969
rect 13083 23913 13139 23969
rect 13225 23913 13281 23969
rect 13367 23913 13423 23969
rect 13509 23913 13565 23969
rect 13651 23913 13707 23969
rect 13793 23913 13849 23969
rect 13935 23913 13991 23969
rect 14077 23913 14133 23969
rect 14219 23913 14275 23969
rect 14361 23913 14417 23969
rect 14503 23913 14559 23969
rect 14645 23913 14701 23969
rect 14787 23913 14843 23969
rect 161 23771 217 23827
rect 303 23771 359 23827
rect 445 23771 501 23827
rect 587 23771 643 23827
rect 729 23771 785 23827
rect 871 23771 927 23827
rect 1013 23771 1069 23827
rect 1155 23771 1211 23827
rect 1297 23771 1353 23827
rect 1439 23771 1495 23827
rect 1581 23771 1637 23827
rect 1723 23771 1779 23827
rect 1865 23771 1921 23827
rect 2007 23771 2063 23827
rect 2149 23771 2205 23827
rect 2291 23771 2347 23827
rect 2433 23771 2489 23827
rect 2575 23771 2631 23827
rect 2717 23771 2773 23827
rect 2859 23771 2915 23827
rect 3001 23771 3057 23827
rect 3143 23771 3199 23827
rect 3285 23771 3341 23827
rect 3427 23771 3483 23827
rect 3569 23771 3625 23827
rect 3711 23771 3767 23827
rect 3853 23771 3909 23827
rect 3995 23771 4051 23827
rect 4137 23771 4193 23827
rect 4279 23771 4335 23827
rect 4421 23771 4477 23827
rect 4563 23771 4619 23827
rect 4705 23771 4761 23827
rect 4847 23771 4903 23827
rect 4989 23771 5045 23827
rect 5131 23771 5187 23827
rect 5273 23771 5329 23827
rect 5415 23771 5471 23827
rect 5557 23771 5613 23827
rect 5699 23771 5755 23827
rect 5841 23771 5897 23827
rect 5983 23771 6039 23827
rect 6125 23771 6181 23827
rect 6267 23771 6323 23827
rect 6409 23771 6465 23827
rect 6551 23771 6607 23827
rect 6693 23771 6749 23827
rect 6835 23771 6891 23827
rect 6977 23771 7033 23827
rect 7119 23771 7175 23827
rect 7261 23771 7317 23827
rect 7403 23771 7459 23827
rect 7545 23771 7601 23827
rect 7687 23771 7743 23827
rect 7829 23771 7885 23827
rect 7971 23771 8027 23827
rect 8113 23771 8169 23827
rect 8255 23771 8311 23827
rect 8397 23771 8453 23827
rect 8539 23771 8595 23827
rect 8681 23771 8737 23827
rect 8823 23771 8879 23827
rect 8965 23771 9021 23827
rect 9107 23771 9163 23827
rect 9249 23771 9305 23827
rect 9391 23771 9447 23827
rect 9533 23771 9589 23827
rect 9675 23771 9731 23827
rect 9817 23771 9873 23827
rect 9959 23771 10015 23827
rect 10101 23771 10157 23827
rect 10243 23771 10299 23827
rect 10385 23771 10441 23827
rect 10527 23771 10583 23827
rect 10669 23771 10725 23827
rect 10811 23771 10867 23827
rect 10953 23771 11009 23827
rect 11095 23771 11151 23827
rect 11237 23771 11293 23827
rect 11379 23771 11435 23827
rect 11521 23771 11577 23827
rect 11663 23771 11719 23827
rect 11805 23771 11861 23827
rect 11947 23771 12003 23827
rect 12089 23771 12145 23827
rect 12231 23771 12287 23827
rect 12373 23771 12429 23827
rect 12515 23771 12571 23827
rect 12657 23771 12713 23827
rect 12799 23771 12855 23827
rect 12941 23771 12997 23827
rect 13083 23771 13139 23827
rect 13225 23771 13281 23827
rect 13367 23771 13423 23827
rect 13509 23771 13565 23827
rect 13651 23771 13707 23827
rect 13793 23771 13849 23827
rect 13935 23771 13991 23827
rect 14077 23771 14133 23827
rect 14219 23771 14275 23827
rect 14361 23771 14417 23827
rect 14503 23771 14559 23827
rect 14645 23771 14701 23827
rect 14787 23771 14843 23827
rect 161 23629 217 23685
rect 303 23629 359 23685
rect 445 23629 501 23685
rect 587 23629 643 23685
rect 729 23629 785 23685
rect 871 23629 927 23685
rect 1013 23629 1069 23685
rect 1155 23629 1211 23685
rect 1297 23629 1353 23685
rect 1439 23629 1495 23685
rect 1581 23629 1637 23685
rect 1723 23629 1779 23685
rect 1865 23629 1921 23685
rect 2007 23629 2063 23685
rect 2149 23629 2205 23685
rect 2291 23629 2347 23685
rect 2433 23629 2489 23685
rect 2575 23629 2631 23685
rect 2717 23629 2773 23685
rect 2859 23629 2915 23685
rect 3001 23629 3057 23685
rect 3143 23629 3199 23685
rect 3285 23629 3341 23685
rect 3427 23629 3483 23685
rect 3569 23629 3625 23685
rect 3711 23629 3767 23685
rect 3853 23629 3909 23685
rect 3995 23629 4051 23685
rect 4137 23629 4193 23685
rect 4279 23629 4335 23685
rect 4421 23629 4477 23685
rect 4563 23629 4619 23685
rect 4705 23629 4761 23685
rect 4847 23629 4903 23685
rect 4989 23629 5045 23685
rect 5131 23629 5187 23685
rect 5273 23629 5329 23685
rect 5415 23629 5471 23685
rect 5557 23629 5613 23685
rect 5699 23629 5755 23685
rect 5841 23629 5897 23685
rect 5983 23629 6039 23685
rect 6125 23629 6181 23685
rect 6267 23629 6323 23685
rect 6409 23629 6465 23685
rect 6551 23629 6607 23685
rect 6693 23629 6749 23685
rect 6835 23629 6891 23685
rect 6977 23629 7033 23685
rect 7119 23629 7175 23685
rect 7261 23629 7317 23685
rect 7403 23629 7459 23685
rect 7545 23629 7601 23685
rect 7687 23629 7743 23685
rect 7829 23629 7885 23685
rect 7971 23629 8027 23685
rect 8113 23629 8169 23685
rect 8255 23629 8311 23685
rect 8397 23629 8453 23685
rect 8539 23629 8595 23685
rect 8681 23629 8737 23685
rect 8823 23629 8879 23685
rect 8965 23629 9021 23685
rect 9107 23629 9163 23685
rect 9249 23629 9305 23685
rect 9391 23629 9447 23685
rect 9533 23629 9589 23685
rect 9675 23629 9731 23685
rect 9817 23629 9873 23685
rect 9959 23629 10015 23685
rect 10101 23629 10157 23685
rect 10243 23629 10299 23685
rect 10385 23629 10441 23685
rect 10527 23629 10583 23685
rect 10669 23629 10725 23685
rect 10811 23629 10867 23685
rect 10953 23629 11009 23685
rect 11095 23629 11151 23685
rect 11237 23629 11293 23685
rect 11379 23629 11435 23685
rect 11521 23629 11577 23685
rect 11663 23629 11719 23685
rect 11805 23629 11861 23685
rect 11947 23629 12003 23685
rect 12089 23629 12145 23685
rect 12231 23629 12287 23685
rect 12373 23629 12429 23685
rect 12515 23629 12571 23685
rect 12657 23629 12713 23685
rect 12799 23629 12855 23685
rect 12941 23629 12997 23685
rect 13083 23629 13139 23685
rect 13225 23629 13281 23685
rect 13367 23629 13423 23685
rect 13509 23629 13565 23685
rect 13651 23629 13707 23685
rect 13793 23629 13849 23685
rect 13935 23629 13991 23685
rect 14077 23629 14133 23685
rect 14219 23629 14275 23685
rect 14361 23629 14417 23685
rect 14503 23629 14559 23685
rect 14645 23629 14701 23685
rect 14787 23629 14843 23685
rect 161 23285 217 23341
rect 303 23285 359 23341
rect 445 23285 501 23341
rect 587 23285 643 23341
rect 729 23285 785 23341
rect 871 23285 927 23341
rect 1013 23285 1069 23341
rect 1155 23285 1211 23341
rect 1297 23285 1353 23341
rect 1439 23285 1495 23341
rect 1581 23285 1637 23341
rect 1723 23285 1779 23341
rect 1865 23285 1921 23341
rect 2007 23285 2063 23341
rect 2149 23285 2205 23341
rect 2291 23285 2347 23341
rect 2433 23285 2489 23341
rect 2575 23285 2631 23341
rect 2717 23285 2773 23341
rect 2859 23285 2915 23341
rect 3001 23285 3057 23341
rect 3143 23285 3199 23341
rect 3285 23285 3341 23341
rect 3427 23285 3483 23341
rect 3569 23285 3625 23341
rect 3711 23285 3767 23341
rect 3853 23285 3909 23341
rect 3995 23285 4051 23341
rect 4137 23285 4193 23341
rect 4279 23285 4335 23341
rect 4421 23285 4477 23341
rect 4563 23285 4619 23341
rect 4705 23285 4761 23341
rect 4847 23285 4903 23341
rect 4989 23285 5045 23341
rect 5131 23285 5187 23341
rect 5273 23285 5329 23341
rect 5415 23285 5471 23341
rect 5557 23285 5613 23341
rect 5699 23285 5755 23341
rect 5841 23285 5897 23341
rect 5983 23285 6039 23341
rect 6125 23285 6181 23341
rect 6267 23285 6323 23341
rect 6409 23285 6465 23341
rect 6551 23285 6607 23341
rect 6693 23285 6749 23341
rect 6835 23285 6891 23341
rect 6977 23285 7033 23341
rect 7119 23285 7175 23341
rect 7261 23285 7317 23341
rect 7403 23285 7459 23341
rect 7545 23285 7601 23341
rect 7687 23285 7743 23341
rect 7829 23285 7885 23341
rect 7971 23285 8027 23341
rect 8113 23285 8169 23341
rect 8255 23285 8311 23341
rect 8397 23285 8453 23341
rect 8539 23285 8595 23341
rect 8681 23285 8737 23341
rect 8823 23285 8879 23341
rect 8965 23285 9021 23341
rect 9107 23285 9163 23341
rect 9249 23285 9305 23341
rect 9391 23285 9447 23341
rect 9533 23285 9589 23341
rect 9675 23285 9731 23341
rect 9817 23285 9873 23341
rect 9959 23285 10015 23341
rect 10101 23285 10157 23341
rect 10243 23285 10299 23341
rect 10385 23285 10441 23341
rect 10527 23285 10583 23341
rect 10669 23285 10725 23341
rect 10811 23285 10867 23341
rect 10953 23285 11009 23341
rect 11095 23285 11151 23341
rect 11237 23285 11293 23341
rect 11379 23285 11435 23341
rect 11521 23285 11577 23341
rect 11663 23285 11719 23341
rect 11805 23285 11861 23341
rect 11947 23285 12003 23341
rect 12089 23285 12145 23341
rect 12231 23285 12287 23341
rect 12373 23285 12429 23341
rect 12515 23285 12571 23341
rect 12657 23285 12713 23341
rect 12799 23285 12855 23341
rect 12941 23285 12997 23341
rect 13083 23285 13139 23341
rect 13225 23285 13281 23341
rect 13367 23285 13423 23341
rect 13509 23285 13565 23341
rect 13651 23285 13707 23341
rect 13793 23285 13849 23341
rect 13935 23285 13991 23341
rect 14077 23285 14133 23341
rect 14219 23285 14275 23341
rect 14361 23285 14417 23341
rect 14503 23285 14559 23341
rect 14645 23285 14701 23341
rect 14787 23285 14843 23341
rect 161 23143 217 23199
rect 303 23143 359 23199
rect 445 23143 501 23199
rect 587 23143 643 23199
rect 729 23143 785 23199
rect 871 23143 927 23199
rect 1013 23143 1069 23199
rect 1155 23143 1211 23199
rect 1297 23143 1353 23199
rect 1439 23143 1495 23199
rect 1581 23143 1637 23199
rect 1723 23143 1779 23199
rect 1865 23143 1921 23199
rect 2007 23143 2063 23199
rect 2149 23143 2205 23199
rect 2291 23143 2347 23199
rect 2433 23143 2489 23199
rect 2575 23143 2631 23199
rect 2717 23143 2773 23199
rect 2859 23143 2915 23199
rect 3001 23143 3057 23199
rect 3143 23143 3199 23199
rect 3285 23143 3341 23199
rect 3427 23143 3483 23199
rect 3569 23143 3625 23199
rect 3711 23143 3767 23199
rect 3853 23143 3909 23199
rect 3995 23143 4051 23199
rect 4137 23143 4193 23199
rect 4279 23143 4335 23199
rect 4421 23143 4477 23199
rect 4563 23143 4619 23199
rect 4705 23143 4761 23199
rect 4847 23143 4903 23199
rect 4989 23143 5045 23199
rect 5131 23143 5187 23199
rect 5273 23143 5329 23199
rect 5415 23143 5471 23199
rect 5557 23143 5613 23199
rect 5699 23143 5755 23199
rect 5841 23143 5897 23199
rect 5983 23143 6039 23199
rect 6125 23143 6181 23199
rect 6267 23143 6323 23199
rect 6409 23143 6465 23199
rect 6551 23143 6607 23199
rect 6693 23143 6749 23199
rect 6835 23143 6891 23199
rect 6977 23143 7033 23199
rect 7119 23143 7175 23199
rect 7261 23143 7317 23199
rect 7403 23143 7459 23199
rect 7545 23143 7601 23199
rect 7687 23143 7743 23199
rect 7829 23143 7885 23199
rect 7971 23143 8027 23199
rect 8113 23143 8169 23199
rect 8255 23143 8311 23199
rect 8397 23143 8453 23199
rect 8539 23143 8595 23199
rect 8681 23143 8737 23199
rect 8823 23143 8879 23199
rect 8965 23143 9021 23199
rect 9107 23143 9163 23199
rect 9249 23143 9305 23199
rect 9391 23143 9447 23199
rect 9533 23143 9589 23199
rect 9675 23143 9731 23199
rect 9817 23143 9873 23199
rect 9959 23143 10015 23199
rect 10101 23143 10157 23199
rect 10243 23143 10299 23199
rect 10385 23143 10441 23199
rect 10527 23143 10583 23199
rect 10669 23143 10725 23199
rect 10811 23143 10867 23199
rect 10953 23143 11009 23199
rect 11095 23143 11151 23199
rect 11237 23143 11293 23199
rect 11379 23143 11435 23199
rect 11521 23143 11577 23199
rect 11663 23143 11719 23199
rect 11805 23143 11861 23199
rect 11947 23143 12003 23199
rect 12089 23143 12145 23199
rect 12231 23143 12287 23199
rect 12373 23143 12429 23199
rect 12515 23143 12571 23199
rect 12657 23143 12713 23199
rect 12799 23143 12855 23199
rect 12941 23143 12997 23199
rect 13083 23143 13139 23199
rect 13225 23143 13281 23199
rect 13367 23143 13423 23199
rect 13509 23143 13565 23199
rect 13651 23143 13707 23199
rect 13793 23143 13849 23199
rect 13935 23143 13991 23199
rect 14077 23143 14133 23199
rect 14219 23143 14275 23199
rect 14361 23143 14417 23199
rect 14503 23143 14559 23199
rect 14645 23143 14701 23199
rect 14787 23143 14843 23199
rect 161 23001 217 23057
rect 303 23001 359 23057
rect 445 23001 501 23057
rect 587 23001 643 23057
rect 729 23001 785 23057
rect 871 23001 927 23057
rect 1013 23001 1069 23057
rect 1155 23001 1211 23057
rect 1297 23001 1353 23057
rect 1439 23001 1495 23057
rect 1581 23001 1637 23057
rect 1723 23001 1779 23057
rect 1865 23001 1921 23057
rect 2007 23001 2063 23057
rect 2149 23001 2205 23057
rect 2291 23001 2347 23057
rect 2433 23001 2489 23057
rect 2575 23001 2631 23057
rect 2717 23001 2773 23057
rect 2859 23001 2915 23057
rect 3001 23001 3057 23057
rect 3143 23001 3199 23057
rect 3285 23001 3341 23057
rect 3427 23001 3483 23057
rect 3569 23001 3625 23057
rect 3711 23001 3767 23057
rect 3853 23001 3909 23057
rect 3995 23001 4051 23057
rect 4137 23001 4193 23057
rect 4279 23001 4335 23057
rect 4421 23001 4477 23057
rect 4563 23001 4619 23057
rect 4705 23001 4761 23057
rect 4847 23001 4903 23057
rect 4989 23001 5045 23057
rect 5131 23001 5187 23057
rect 5273 23001 5329 23057
rect 5415 23001 5471 23057
rect 5557 23001 5613 23057
rect 5699 23001 5755 23057
rect 5841 23001 5897 23057
rect 5983 23001 6039 23057
rect 6125 23001 6181 23057
rect 6267 23001 6323 23057
rect 6409 23001 6465 23057
rect 6551 23001 6607 23057
rect 6693 23001 6749 23057
rect 6835 23001 6891 23057
rect 6977 23001 7033 23057
rect 7119 23001 7175 23057
rect 7261 23001 7317 23057
rect 7403 23001 7459 23057
rect 7545 23001 7601 23057
rect 7687 23001 7743 23057
rect 7829 23001 7885 23057
rect 7971 23001 8027 23057
rect 8113 23001 8169 23057
rect 8255 23001 8311 23057
rect 8397 23001 8453 23057
rect 8539 23001 8595 23057
rect 8681 23001 8737 23057
rect 8823 23001 8879 23057
rect 8965 23001 9021 23057
rect 9107 23001 9163 23057
rect 9249 23001 9305 23057
rect 9391 23001 9447 23057
rect 9533 23001 9589 23057
rect 9675 23001 9731 23057
rect 9817 23001 9873 23057
rect 9959 23001 10015 23057
rect 10101 23001 10157 23057
rect 10243 23001 10299 23057
rect 10385 23001 10441 23057
rect 10527 23001 10583 23057
rect 10669 23001 10725 23057
rect 10811 23001 10867 23057
rect 10953 23001 11009 23057
rect 11095 23001 11151 23057
rect 11237 23001 11293 23057
rect 11379 23001 11435 23057
rect 11521 23001 11577 23057
rect 11663 23001 11719 23057
rect 11805 23001 11861 23057
rect 11947 23001 12003 23057
rect 12089 23001 12145 23057
rect 12231 23001 12287 23057
rect 12373 23001 12429 23057
rect 12515 23001 12571 23057
rect 12657 23001 12713 23057
rect 12799 23001 12855 23057
rect 12941 23001 12997 23057
rect 13083 23001 13139 23057
rect 13225 23001 13281 23057
rect 13367 23001 13423 23057
rect 13509 23001 13565 23057
rect 13651 23001 13707 23057
rect 13793 23001 13849 23057
rect 13935 23001 13991 23057
rect 14077 23001 14133 23057
rect 14219 23001 14275 23057
rect 14361 23001 14417 23057
rect 14503 23001 14559 23057
rect 14645 23001 14701 23057
rect 14787 23001 14843 23057
rect 161 22859 217 22915
rect 303 22859 359 22915
rect 445 22859 501 22915
rect 587 22859 643 22915
rect 729 22859 785 22915
rect 871 22859 927 22915
rect 1013 22859 1069 22915
rect 1155 22859 1211 22915
rect 1297 22859 1353 22915
rect 1439 22859 1495 22915
rect 1581 22859 1637 22915
rect 1723 22859 1779 22915
rect 1865 22859 1921 22915
rect 2007 22859 2063 22915
rect 2149 22859 2205 22915
rect 2291 22859 2347 22915
rect 2433 22859 2489 22915
rect 2575 22859 2631 22915
rect 2717 22859 2773 22915
rect 2859 22859 2915 22915
rect 3001 22859 3057 22915
rect 3143 22859 3199 22915
rect 3285 22859 3341 22915
rect 3427 22859 3483 22915
rect 3569 22859 3625 22915
rect 3711 22859 3767 22915
rect 3853 22859 3909 22915
rect 3995 22859 4051 22915
rect 4137 22859 4193 22915
rect 4279 22859 4335 22915
rect 4421 22859 4477 22915
rect 4563 22859 4619 22915
rect 4705 22859 4761 22915
rect 4847 22859 4903 22915
rect 4989 22859 5045 22915
rect 5131 22859 5187 22915
rect 5273 22859 5329 22915
rect 5415 22859 5471 22915
rect 5557 22859 5613 22915
rect 5699 22859 5755 22915
rect 5841 22859 5897 22915
rect 5983 22859 6039 22915
rect 6125 22859 6181 22915
rect 6267 22859 6323 22915
rect 6409 22859 6465 22915
rect 6551 22859 6607 22915
rect 6693 22859 6749 22915
rect 6835 22859 6891 22915
rect 6977 22859 7033 22915
rect 7119 22859 7175 22915
rect 7261 22859 7317 22915
rect 7403 22859 7459 22915
rect 7545 22859 7601 22915
rect 7687 22859 7743 22915
rect 7829 22859 7885 22915
rect 7971 22859 8027 22915
rect 8113 22859 8169 22915
rect 8255 22859 8311 22915
rect 8397 22859 8453 22915
rect 8539 22859 8595 22915
rect 8681 22859 8737 22915
rect 8823 22859 8879 22915
rect 8965 22859 9021 22915
rect 9107 22859 9163 22915
rect 9249 22859 9305 22915
rect 9391 22859 9447 22915
rect 9533 22859 9589 22915
rect 9675 22859 9731 22915
rect 9817 22859 9873 22915
rect 9959 22859 10015 22915
rect 10101 22859 10157 22915
rect 10243 22859 10299 22915
rect 10385 22859 10441 22915
rect 10527 22859 10583 22915
rect 10669 22859 10725 22915
rect 10811 22859 10867 22915
rect 10953 22859 11009 22915
rect 11095 22859 11151 22915
rect 11237 22859 11293 22915
rect 11379 22859 11435 22915
rect 11521 22859 11577 22915
rect 11663 22859 11719 22915
rect 11805 22859 11861 22915
rect 11947 22859 12003 22915
rect 12089 22859 12145 22915
rect 12231 22859 12287 22915
rect 12373 22859 12429 22915
rect 12515 22859 12571 22915
rect 12657 22859 12713 22915
rect 12799 22859 12855 22915
rect 12941 22859 12997 22915
rect 13083 22859 13139 22915
rect 13225 22859 13281 22915
rect 13367 22859 13423 22915
rect 13509 22859 13565 22915
rect 13651 22859 13707 22915
rect 13793 22859 13849 22915
rect 13935 22859 13991 22915
rect 14077 22859 14133 22915
rect 14219 22859 14275 22915
rect 14361 22859 14417 22915
rect 14503 22859 14559 22915
rect 14645 22859 14701 22915
rect 14787 22859 14843 22915
rect 161 22717 217 22773
rect 303 22717 359 22773
rect 445 22717 501 22773
rect 587 22717 643 22773
rect 729 22717 785 22773
rect 871 22717 927 22773
rect 1013 22717 1069 22773
rect 1155 22717 1211 22773
rect 1297 22717 1353 22773
rect 1439 22717 1495 22773
rect 1581 22717 1637 22773
rect 1723 22717 1779 22773
rect 1865 22717 1921 22773
rect 2007 22717 2063 22773
rect 2149 22717 2205 22773
rect 2291 22717 2347 22773
rect 2433 22717 2489 22773
rect 2575 22717 2631 22773
rect 2717 22717 2773 22773
rect 2859 22717 2915 22773
rect 3001 22717 3057 22773
rect 3143 22717 3199 22773
rect 3285 22717 3341 22773
rect 3427 22717 3483 22773
rect 3569 22717 3625 22773
rect 3711 22717 3767 22773
rect 3853 22717 3909 22773
rect 3995 22717 4051 22773
rect 4137 22717 4193 22773
rect 4279 22717 4335 22773
rect 4421 22717 4477 22773
rect 4563 22717 4619 22773
rect 4705 22717 4761 22773
rect 4847 22717 4903 22773
rect 4989 22717 5045 22773
rect 5131 22717 5187 22773
rect 5273 22717 5329 22773
rect 5415 22717 5471 22773
rect 5557 22717 5613 22773
rect 5699 22717 5755 22773
rect 5841 22717 5897 22773
rect 5983 22717 6039 22773
rect 6125 22717 6181 22773
rect 6267 22717 6323 22773
rect 6409 22717 6465 22773
rect 6551 22717 6607 22773
rect 6693 22717 6749 22773
rect 6835 22717 6891 22773
rect 6977 22717 7033 22773
rect 7119 22717 7175 22773
rect 7261 22717 7317 22773
rect 7403 22717 7459 22773
rect 7545 22717 7601 22773
rect 7687 22717 7743 22773
rect 7829 22717 7885 22773
rect 7971 22717 8027 22773
rect 8113 22717 8169 22773
rect 8255 22717 8311 22773
rect 8397 22717 8453 22773
rect 8539 22717 8595 22773
rect 8681 22717 8737 22773
rect 8823 22717 8879 22773
rect 8965 22717 9021 22773
rect 9107 22717 9163 22773
rect 9249 22717 9305 22773
rect 9391 22717 9447 22773
rect 9533 22717 9589 22773
rect 9675 22717 9731 22773
rect 9817 22717 9873 22773
rect 9959 22717 10015 22773
rect 10101 22717 10157 22773
rect 10243 22717 10299 22773
rect 10385 22717 10441 22773
rect 10527 22717 10583 22773
rect 10669 22717 10725 22773
rect 10811 22717 10867 22773
rect 10953 22717 11009 22773
rect 11095 22717 11151 22773
rect 11237 22717 11293 22773
rect 11379 22717 11435 22773
rect 11521 22717 11577 22773
rect 11663 22717 11719 22773
rect 11805 22717 11861 22773
rect 11947 22717 12003 22773
rect 12089 22717 12145 22773
rect 12231 22717 12287 22773
rect 12373 22717 12429 22773
rect 12515 22717 12571 22773
rect 12657 22717 12713 22773
rect 12799 22717 12855 22773
rect 12941 22717 12997 22773
rect 13083 22717 13139 22773
rect 13225 22717 13281 22773
rect 13367 22717 13423 22773
rect 13509 22717 13565 22773
rect 13651 22717 13707 22773
rect 13793 22717 13849 22773
rect 13935 22717 13991 22773
rect 14077 22717 14133 22773
rect 14219 22717 14275 22773
rect 14361 22717 14417 22773
rect 14503 22717 14559 22773
rect 14645 22717 14701 22773
rect 14787 22717 14843 22773
rect 161 22575 217 22631
rect 303 22575 359 22631
rect 445 22575 501 22631
rect 587 22575 643 22631
rect 729 22575 785 22631
rect 871 22575 927 22631
rect 1013 22575 1069 22631
rect 1155 22575 1211 22631
rect 1297 22575 1353 22631
rect 1439 22575 1495 22631
rect 1581 22575 1637 22631
rect 1723 22575 1779 22631
rect 1865 22575 1921 22631
rect 2007 22575 2063 22631
rect 2149 22575 2205 22631
rect 2291 22575 2347 22631
rect 2433 22575 2489 22631
rect 2575 22575 2631 22631
rect 2717 22575 2773 22631
rect 2859 22575 2915 22631
rect 3001 22575 3057 22631
rect 3143 22575 3199 22631
rect 3285 22575 3341 22631
rect 3427 22575 3483 22631
rect 3569 22575 3625 22631
rect 3711 22575 3767 22631
rect 3853 22575 3909 22631
rect 3995 22575 4051 22631
rect 4137 22575 4193 22631
rect 4279 22575 4335 22631
rect 4421 22575 4477 22631
rect 4563 22575 4619 22631
rect 4705 22575 4761 22631
rect 4847 22575 4903 22631
rect 4989 22575 5045 22631
rect 5131 22575 5187 22631
rect 5273 22575 5329 22631
rect 5415 22575 5471 22631
rect 5557 22575 5613 22631
rect 5699 22575 5755 22631
rect 5841 22575 5897 22631
rect 5983 22575 6039 22631
rect 6125 22575 6181 22631
rect 6267 22575 6323 22631
rect 6409 22575 6465 22631
rect 6551 22575 6607 22631
rect 6693 22575 6749 22631
rect 6835 22575 6891 22631
rect 6977 22575 7033 22631
rect 7119 22575 7175 22631
rect 7261 22575 7317 22631
rect 7403 22575 7459 22631
rect 7545 22575 7601 22631
rect 7687 22575 7743 22631
rect 7829 22575 7885 22631
rect 7971 22575 8027 22631
rect 8113 22575 8169 22631
rect 8255 22575 8311 22631
rect 8397 22575 8453 22631
rect 8539 22575 8595 22631
rect 8681 22575 8737 22631
rect 8823 22575 8879 22631
rect 8965 22575 9021 22631
rect 9107 22575 9163 22631
rect 9249 22575 9305 22631
rect 9391 22575 9447 22631
rect 9533 22575 9589 22631
rect 9675 22575 9731 22631
rect 9817 22575 9873 22631
rect 9959 22575 10015 22631
rect 10101 22575 10157 22631
rect 10243 22575 10299 22631
rect 10385 22575 10441 22631
rect 10527 22575 10583 22631
rect 10669 22575 10725 22631
rect 10811 22575 10867 22631
rect 10953 22575 11009 22631
rect 11095 22575 11151 22631
rect 11237 22575 11293 22631
rect 11379 22575 11435 22631
rect 11521 22575 11577 22631
rect 11663 22575 11719 22631
rect 11805 22575 11861 22631
rect 11947 22575 12003 22631
rect 12089 22575 12145 22631
rect 12231 22575 12287 22631
rect 12373 22575 12429 22631
rect 12515 22575 12571 22631
rect 12657 22575 12713 22631
rect 12799 22575 12855 22631
rect 12941 22575 12997 22631
rect 13083 22575 13139 22631
rect 13225 22575 13281 22631
rect 13367 22575 13423 22631
rect 13509 22575 13565 22631
rect 13651 22575 13707 22631
rect 13793 22575 13849 22631
rect 13935 22575 13991 22631
rect 14077 22575 14133 22631
rect 14219 22575 14275 22631
rect 14361 22575 14417 22631
rect 14503 22575 14559 22631
rect 14645 22575 14701 22631
rect 14787 22575 14843 22631
rect 161 22433 217 22489
rect 303 22433 359 22489
rect 445 22433 501 22489
rect 587 22433 643 22489
rect 729 22433 785 22489
rect 871 22433 927 22489
rect 1013 22433 1069 22489
rect 1155 22433 1211 22489
rect 1297 22433 1353 22489
rect 1439 22433 1495 22489
rect 1581 22433 1637 22489
rect 1723 22433 1779 22489
rect 1865 22433 1921 22489
rect 2007 22433 2063 22489
rect 2149 22433 2205 22489
rect 2291 22433 2347 22489
rect 2433 22433 2489 22489
rect 2575 22433 2631 22489
rect 2717 22433 2773 22489
rect 2859 22433 2915 22489
rect 3001 22433 3057 22489
rect 3143 22433 3199 22489
rect 3285 22433 3341 22489
rect 3427 22433 3483 22489
rect 3569 22433 3625 22489
rect 3711 22433 3767 22489
rect 3853 22433 3909 22489
rect 3995 22433 4051 22489
rect 4137 22433 4193 22489
rect 4279 22433 4335 22489
rect 4421 22433 4477 22489
rect 4563 22433 4619 22489
rect 4705 22433 4761 22489
rect 4847 22433 4903 22489
rect 4989 22433 5045 22489
rect 5131 22433 5187 22489
rect 5273 22433 5329 22489
rect 5415 22433 5471 22489
rect 5557 22433 5613 22489
rect 5699 22433 5755 22489
rect 5841 22433 5897 22489
rect 5983 22433 6039 22489
rect 6125 22433 6181 22489
rect 6267 22433 6323 22489
rect 6409 22433 6465 22489
rect 6551 22433 6607 22489
rect 6693 22433 6749 22489
rect 6835 22433 6891 22489
rect 6977 22433 7033 22489
rect 7119 22433 7175 22489
rect 7261 22433 7317 22489
rect 7403 22433 7459 22489
rect 7545 22433 7601 22489
rect 7687 22433 7743 22489
rect 7829 22433 7885 22489
rect 7971 22433 8027 22489
rect 8113 22433 8169 22489
rect 8255 22433 8311 22489
rect 8397 22433 8453 22489
rect 8539 22433 8595 22489
rect 8681 22433 8737 22489
rect 8823 22433 8879 22489
rect 8965 22433 9021 22489
rect 9107 22433 9163 22489
rect 9249 22433 9305 22489
rect 9391 22433 9447 22489
rect 9533 22433 9589 22489
rect 9675 22433 9731 22489
rect 9817 22433 9873 22489
rect 9959 22433 10015 22489
rect 10101 22433 10157 22489
rect 10243 22433 10299 22489
rect 10385 22433 10441 22489
rect 10527 22433 10583 22489
rect 10669 22433 10725 22489
rect 10811 22433 10867 22489
rect 10953 22433 11009 22489
rect 11095 22433 11151 22489
rect 11237 22433 11293 22489
rect 11379 22433 11435 22489
rect 11521 22433 11577 22489
rect 11663 22433 11719 22489
rect 11805 22433 11861 22489
rect 11947 22433 12003 22489
rect 12089 22433 12145 22489
rect 12231 22433 12287 22489
rect 12373 22433 12429 22489
rect 12515 22433 12571 22489
rect 12657 22433 12713 22489
rect 12799 22433 12855 22489
rect 12941 22433 12997 22489
rect 13083 22433 13139 22489
rect 13225 22433 13281 22489
rect 13367 22433 13423 22489
rect 13509 22433 13565 22489
rect 13651 22433 13707 22489
rect 13793 22433 13849 22489
rect 13935 22433 13991 22489
rect 14077 22433 14133 22489
rect 14219 22433 14275 22489
rect 14361 22433 14417 22489
rect 14503 22433 14559 22489
rect 14645 22433 14701 22489
rect 14787 22433 14843 22489
rect 161 22291 217 22347
rect 303 22291 359 22347
rect 445 22291 501 22347
rect 587 22291 643 22347
rect 729 22291 785 22347
rect 871 22291 927 22347
rect 1013 22291 1069 22347
rect 1155 22291 1211 22347
rect 1297 22291 1353 22347
rect 1439 22291 1495 22347
rect 1581 22291 1637 22347
rect 1723 22291 1779 22347
rect 1865 22291 1921 22347
rect 2007 22291 2063 22347
rect 2149 22291 2205 22347
rect 2291 22291 2347 22347
rect 2433 22291 2489 22347
rect 2575 22291 2631 22347
rect 2717 22291 2773 22347
rect 2859 22291 2915 22347
rect 3001 22291 3057 22347
rect 3143 22291 3199 22347
rect 3285 22291 3341 22347
rect 3427 22291 3483 22347
rect 3569 22291 3625 22347
rect 3711 22291 3767 22347
rect 3853 22291 3909 22347
rect 3995 22291 4051 22347
rect 4137 22291 4193 22347
rect 4279 22291 4335 22347
rect 4421 22291 4477 22347
rect 4563 22291 4619 22347
rect 4705 22291 4761 22347
rect 4847 22291 4903 22347
rect 4989 22291 5045 22347
rect 5131 22291 5187 22347
rect 5273 22291 5329 22347
rect 5415 22291 5471 22347
rect 5557 22291 5613 22347
rect 5699 22291 5755 22347
rect 5841 22291 5897 22347
rect 5983 22291 6039 22347
rect 6125 22291 6181 22347
rect 6267 22291 6323 22347
rect 6409 22291 6465 22347
rect 6551 22291 6607 22347
rect 6693 22291 6749 22347
rect 6835 22291 6891 22347
rect 6977 22291 7033 22347
rect 7119 22291 7175 22347
rect 7261 22291 7317 22347
rect 7403 22291 7459 22347
rect 7545 22291 7601 22347
rect 7687 22291 7743 22347
rect 7829 22291 7885 22347
rect 7971 22291 8027 22347
rect 8113 22291 8169 22347
rect 8255 22291 8311 22347
rect 8397 22291 8453 22347
rect 8539 22291 8595 22347
rect 8681 22291 8737 22347
rect 8823 22291 8879 22347
rect 8965 22291 9021 22347
rect 9107 22291 9163 22347
rect 9249 22291 9305 22347
rect 9391 22291 9447 22347
rect 9533 22291 9589 22347
rect 9675 22291 9731 22347
rect 9817 22291 9873 22347
rect 9959 22291 10015 22347
rect 10101 22291 10157 22347
rect 10243 22291 10299 22347
rect 10385 22291 10441 22347
rect 10527 22291 10583 22347
rect 10669 22291 10725 22347
rect 10811 22291 10867 22347
rect 10953 22291 11009 22347
rect 11095 22291 11151 22347
rect 11237 22291 11293 22347
rect 11379 22291 11435 22347
rect 11521 22291 11577 22347
rect 11663 22291 11719 22347
rect 11805 22291 11861 22347
rect 11947 22291 12003 22347
rect 12089 22291 12145 22347
rect 12231 22291 12287 22347
rect 12373 22291 12429 22347
rect 12515 22291 12571 22347
rect 12657 22291 12713 22347
rect 12799 22291 12855 22347
rect 12941 22291 12997 22347
rect 13083 22291 13139 22347
rect 13225 22291 13281 22347
rect 13367 22291 13423 22347
rect 13509 22291 13565 22347
rect 13651 22291 13707 22347
rect 13793 22291 13849 22347
rect 13935 22291 13991 22347
rect 14077 22291 14133 22347
rect 14219 22291 14275 22347
rect 14361 22291 14417 22347
rect 14503 22291 14559 22347
rect 14645 22291 14701 22347
rect 14787 22291 14843 22347
rect 161 22149 217 22205
rect 303 22149 359 22205
rect 445 22149 501 22205
rect 587 22149 643 22205
rect 729 22149 785 22205
rect 871 22149 927 22205
rect 1013 22149 1069 22205
rect 1155 22149 1211 22205
rect 1297 22149 1353 22205
rect 1439 22149 1495 22205
rect 1581 22149 1637 22205
rect 1723 22149 1779 22205
rect 1865 22149 1921 22205
rect 2007 22149 2063 22205
rect 2149 22149 2205 22205
rect 2291 22149 2347 22205
rect 2433 22149 2489 22205
rect 2575 22149 2631 22205
rect 2717 22149 2773 22205
rect 2859 22149 2915 22205
rect 3001 22149 3057 22205
rect 3143 22149 3199 22205
rect 3285 22149 3341 22205
rect 3427 22149 3483 22205
rect 3569 22149 3625 22205
rect 3711 22149 3767 22205
rect 3853 22149 3909 22205
rect 3995 22149 4051 22205
rect 4137 22149 4193 22205
rect 4279 22149 4335 22205
rect 4421 22149 4477 22205
rect 4563 22149 4619 22205
rect 4705 22149 4761 22205
rect 4847 22149 4903 22205
rect 4989 22149 5045 22205
rect 5131 22149 5187 22205
rect 5273 22149 5329 22205
rect 5415 22149 5471 22205
rect 5557 22149 5613 22205
rect 5699 22149 5755 22205
rect 5841 22149 5897 22205
rect 5983 22149 6039 22205
rect 6125 22149 6181 22205
rect 6267 22149 6323 22205
rect 6409 22149 6465 22205
rect 6551 22149 6607 22205
rect 6693 22149 6749 22205
rect 6835 22149 6891 22205
rect 6977 22149 7033 22205
rect 7119 22149 7175 22205
rect 7261 22149 7317 22205
rect 7403 22149 7459 22205
rect 7545 22149 7601 22205
rect 7687 22149 7743 22205
rect 7829 22149 7885 22205
rect 7971 22149 8027 22205
rect 8113 22149 8169 22205
rect 8255 22149 8311 22205
rect 8397 22149 8453 22205
rect 8539 22149 8595 22205
rect 8681 22149 8737 22205
rect 8823 22149 8879 22205
rect 8965 22149 9021 22205
rect 9107 22149 9163 22205
rect 9249 22149 9305 22205
rect 9391 22149 9447 22205
rect 9533 22149 9589 22205
rect 9675 22149 9731 22205
rect 9817 22149 9873 22205
rect 9959 22149 10015 22205
rect 10101 22149 10157 22205
rect 10243 22149 10299 22205
rect 10385 22149 10441 22205
rect 10527 22149 10583 22205
rect 10669 22149 10725 22205
rect 10811 22149 10867 22205
rect 10953 22149 11009 22205
rect 11095 22149 11151 22205
rect 11237 22149 11293 22205
rect 11379 22149 11435 22205
rect 11521 22149 11577 22205
rect 11663 22149 11719 22205
rect 11805 22149 11861 22205
rect 11947 22149 12003 22205
rect 12089 22149 12145 22205
rect 12231 22149 12287 22205
rect 12373 22149 12429 22205
rect 12515 22149 12571 22205
rect 12657 22149 12713 22205
rect 12799 22149 12855 22205
rect 12941 22149 12997 22205
rect 13083 22149 13139 22205
rect 13225 22149 13281 22205
rect 13367 22149 13423 22205
rect 13509 22149 13565 22205
rect 13651 22149 13707 22205
rect 13793 22149 13849 22205
rect 13935 22149 13991 22205
rect 14077 22149 14133 22205
rect 14219 22149 14275 22205
rect 14361 22149 14417 22205
rect 14503 22149 14559 22205
rect 14645 22149 14701 22205
rect 14787 22149 14843 22205
rect 161 22007 217 22063
rect 303 22007 359 22063
rect 445 22007 501 22063
rect 587 22007 643 22063
rect 729 22007 785 22063
rect 871 22007 927 22063
rect 1013 22007 1069 22063
rect 1155 22007 1211 22063
rect 1297 22007 1353 22063
rect 1439 22007 1495 22063
rect 1581 22007 1637 22063
rect 1723 22007 1779 22063
rect 1865 22007 1921 22063
rect 2007 22007 2063 22063
rect 2149 22007 2205 22063
rect 2291 22007 2347 22063
rect 2433 22007 2489 22063
rect 2575 22007 2631 22063
rect 2717 22007 2773 22063
rect 2859 22007 2915 22063
rect 3001 22007 3057 22063
rect 3143 22007 3199 22063
rect 3285 22007 3341 22063
rect 3427 22007 3483 22063
rect 3569 22007 3625 22063
rect 3711 22007 3767 22063
rect 3853 22007 3909 22063
rect 3995 22007 4051 22063
rect 4137 22007 4193 22063
rect 4279 22007 4335 22063
rect 4421 22007 4477 22063
rect 4563 22007 4619 22063
rect 4705 22007 4761 22063
rect 4847 22007 4903 22063
rect 4989 22007 5045 22063
rect 5131 22007 5187 22063
rect 5273 22007 5329 22063
rect 5415 22007 5471 22063
rect 5557 22007 5613 22063
rect 5699 22007 5755 22063
rect 5841 22007 5897 22063
rect 5983 22007 6039 22063
rect 6125 22007 6181 22063
rect 6267 22007 6323 22063
rect 6409 22007 6465 22063
rect 6551 22007 6607 22063
rect 6693 22007 6749 22063
rect 6835 22007 6891 22063
rect 6977 22007 7033 22063
rect 7119 22007 7175 22063
rect 7261 22007 7317 22063
rect 7403 22007 7459 22063
rect 7545 22007 7601 22063
rect 7687 22007 7743 22063
rect 7829 22007 7885 22063
rect 7971 22007 8027 22063
rect 8113 22007 8169 22063
rect 8255 22007 8311 22063
rect 8397 22007 8453 22063
rect 8539 22007 8595 22063
rect 8681 22007 8737 22063
rect 8823 22007 8879 22063
rect 8965 22007 9021 22063
rect 9107 22007 9163 22063
rect 9249 22007 9305 22063
rect 9391 22007 9447 22063
rect 9533 22007 9589 22063
rect 9675 22007 9731 22063
rect 9817 22007 9873 22063
rect 9959 22007 10015 22063
rect 10101 22007 10157 22063
rect 10243 22007 10299 22063
rect 10385 22007 10441 22063
rect 10527 22007 10583 22063
rect 10669 22007 10725 22063
rect 10811 22007 10867 22063
rect 10953 22007 11009 22063
rect 11095 22007 11151 22063
rect 11237 22007 11293 22063
rect 11379 22007 11435 22063
rect 11521 22007 11577 22063
rect 11663 22007 11719 22063
rect 11805 22007 11861 22063
rect 11947 22007 12003 22063
rect 12089 22007 12145 22063
rect 12231 22007 12287 22063
rect 12373 22007 12429 22063
rect 12515 22007 12571 22063
rect 12657 22007 12713 22063
rect 12799 22007 12855 22063
rect 12941 22007 12997 22063
rect 13083 22007 13139 22063
rect 13225 22007 13281 22063
rect 13367 22007 13423 22063
rect 13509 22007 13565 22063
rect 13651 22007 13707 22063
rect 13793 22007 13849 22063
rect 13935 22007 13991 22063
rect 14077 22007 14133 22063
rect 14219 22007 14275 22063
rect 14361 22007 14417 22063
rect 14503 22007 14559 22063
rect 14645 22007 14701 22063
rect 14787 22007 14843 22063
rect 161 21865 217 21921
rect 303 21865 359 21921
rect 445 21865 501 21921
rect 587 21865 643 21921
rect 729 21865 785 21921
rect 871 21865 927 21921
rect 1013 21865 1069 21921
rect 1155 21865 1211 21921
rect 1297 21865 1353 21921
rect 1439 21865 1495 21921
rect 1581 21865 1637 21921
rect 1723 21865 1779 21921
rect 1865 21865 1921 21921
rect 2007 21865 2063 21921
rect 2149 21865 2205 21921
rect 2291 21865 2347 21921
rect 2433 21865 2489 21921
rect 2575 21865 2631 21921
rect 2717 21865 2773 21921
rect 2859 21865 2915 21921
rect 3001 21865 3057 21921
rect 3143 21865 3199 21921
rect 3285 21865 3341 21921
rect 3427 21865 3483 21921
rect 3569 21865 3625 21921
rect 3711 21865 3767 21921
rect 3853 21865 3909 21921
rect 3995 21865 4051 21921
rect 4137 21865 4193 21921
rect 4279 21865 4335 21921
rect 4421 21865 4477 21921
rect 4563 21865 4619 21921
rect 4705 21865 4761 21921
rect 4847 21865 4903 21921
rect 4989 21865 5045 21921
rect 5131 21865 5187 21921
rect 5273 21865 5329 21921
rect 5415 21865 5471 21921
rect 5557 21865 5613 21921
rect 5699 21865 5755 21921
rect 5841 21865 5897 21921
rect 5983 21865 6039 21921
rect 6125 21865 6181 21921
rect 6267 21865 6323 21921
rect 6409 21865 6465 21921
rect 6551 21865 6607 21921
rect 6693 21865 6749 21921
rect 6835 21865 6891 21921
rect 6977 21865 7033 21921
rect 7119 21865 7175 21921
rect 7261 21865 7317 21921
rect 7403 21865 7459 21921
rect 7545 21865 7601 21921
rect 7687 21865 7743 21921
rect 7829 21865 7885 21921
rect 7971 21865 8027 21921
rect 8113 21865 8169 21921
rect 8255 21865 8311 21921
rect 8397 21865 8453 21921
rect 8539 21865 8595 21921
rect 8681 21865 8737 21921
rect 8823 21865 8879 21921
rect 8965 21865 9021 21921
rect 9107 21865 9163 21921
rect 9249 21865 9305 21921
rect 9391 21865 9447 21921
rect 9533 21865 9589 21921
rect 9675 21865 9731 21921
rect 9817 21865 9873 21921
rect 9959 21865 10015 21921
rect 10101 21865 10157 21921
rect 10243 21865 10299 21921
rect 10385 21865 10441 21921
rect 10527 21865 10583 21921
rect 10669 21865 10725 21921
rect 10811 21865 10867 21921
rect 10953 21865 11009 21921
rect 11095 21865 11151 21921
rect 11237 21865 11293 21921
rect 11379 21865 11435 21921
rect 11521 21865 11577 21921
rect 11663 21865 11719 21921
rect 11805 21865 11861 21921
rect 11947 21865 12003 21921
rect 12089 21865 12145 21921
rect 12231 21865 12287 21921
rect 12373 21865 12429 21921
rect 12515 21865 12571 21921
rect 12657 21865 12713 21921
rect 12799 21865 12855 21921
rect 12941 21865 12997 21921
rect 13083 21865 13139 21921
rect 13225 21865 13281 21921
rect 13367 21865 13423 21921
rect 13509 21865 13565 21921
rect 13651 21865 13707 21921
rect 13793 21865 13849 21921
rect 13935 21865 13991 21921
rect 14077 21865 14133 21921
rect 14219 21865 14275 21921
rect 14361 21865 14417 21921
rect 14503 21865 14559 21921
rect 14645 21865 14701 21921
rect 14787 21865 14843 21921
rect 161 21723 217 21779
rect 303 21723 359 21779
rect 445 21723 501 21779
rect 587 21723 643 21779
rect 729 21723 785 21779
rect 871 21723 927 21779
rect 1013 21723 1069 21779
rect 1155 21723 1211 21779
rect 1297 21723 1353 21779
rect 1439 21723 1495 21779
rect 1581 21723 1637 21779
rect 1723 21723 1779 21779
rect 1865 21723 1921 21779
rect 2007 21723 2063 21779
rect 2149 21723 2205 21779
rect 2291 21723 2347 21779
rect 2433 21723 2489 21779
rect 2575 21723 2631 21779
rect 2717 21723 2773 21779
rect 2859 21723 2915 21779
rect 3001 21723 3057 21779
rect 3143 21723 3199 21779
rect 3285 21723 3341 21779
rect 3427 21723 3483 21779
rect 3569 21723 3625 21779
rect 3711 21723 3767 21779
rect 3853 21723 3909 21779
rect 3995 21723 4051 21779
rect 4137 21723 4193 21779
rect 4279 21723 4335 21779
rect 4421 21723 4477 21779
rect 4563 21723 4619 21779
rect 4705 21723 4761 21779
rect 4847 21723 4903 21779
rect 4989 21723 5045 21779
rect 5131 21723 5187 21779
rect 5273 21723 5329 21779
rect 5415 21723 5471 21779
rect 5557 21723 5613 21779
rect 5699 21723 5755 21779
rect 5841 21723 5897 21779
rect 5983 21723 6039 21779
rect 6125 21723 6181 21779
rect 6267 21723 6323 21779
rect 6409 21723 6465 21779
rect 6551 21723 6607 21779
rect 6693 21723 6749 21779
rect 6835 21723 6891 21779
rect 6977 21723 7033 21779
rect 7119 21723 7175 21779
rect 7261 21723 7317 21779
rect 7403 21723 7459 21779
rect 7545 21723 7601 21779
rect 7687 21723 7743 21779
rect 7829 21723 7885 21779
rect 7971 21723 8027 21779
rect 8113 21723 8169 21779
rect 8255 21723 8311 21779
rect 8397 21723 8453 21779
rect 8539 21723 8595 21779
rect 8681 21723 8737 21779
rect 8823 21723 8879 21779
rect 8965 21723 9021 21779
rect 9107 21723 9163 21779
rect 9249 21723 9305 21779
rect 9391 21723 9447 21779
rect 9533 21723 9589 21779
rect 9675 21723 9731 21779
rect 9817 21723 9873 21779
rect 9959 21723 10015 21779
rect 10101 21723 10157 21779
rect 10243 21723 10299 21779
rect 10385 21723 10441 21779
rect 10527 21723 10583 21779
rect 10669 21723 10725 21779
rect 10811 21723 10867 21779
rect 10953 21723 11009 21779
rect 11095 21723 11151 21779
rect 11237 21723 11293 21779
rect 11379 21723 11435 21779
rect 11521 21723 11577 21779
rect 11663 21723 11719 21779
rect 11805 21723 11861 21779
rect 11947 21723 12003 21779
rect 12089 21723 12145 21779
rect 12231 21723 12287 21779
rect 12373 21723 12429 21779
rect 12515 21723 12571 21779
rect 12657 21723 12713 21779
rect 12799 21723 12855 21779
rect 12941 21723 12997 21779
rect 13083 21723 13139 21779
rect 13225 21723 13281 21779
rect 13367 21723 13423 21779
rect 13509 21723 13565 21779
rect 13651 21723 13707 21779
rect 13793 21723 13849 21779
rect 13935 21723 13991 21779
rect 14077 21723 14133 21779
rect 14219 21723 14275 21779
rect 14361 21723 14417 21779
rect 14503 21723 14559 21779
rect 14645 21723 14701 21779
rect 14787 21723 14843 21779
rect 161 21581 217 21637
rect 303 21581 359 21637
rect 445 21581 501 21637
rect 587 21581 643 21637
rect 729 21581 785 21637
rect 871 21581 927 21637
rect 1013 21581 1069 21637
rect 1155 21581 1211 21637
rect 1297 21581 1353 21637
rect 1439 21581 1495 21637
rect 1581 21581 1637 21637
rect 1723 21581 1779 21637
rect 1865 21581 1921 21637
rect 2007 21581 2063 21637
rect 2149 21581 2205 21637
rect 2291 21581 2347 21637
rect 2433 21581 2489 21637
rect 2575 21581 2631 21637
rect 2717 21581 2773 21637
rect 2859 21581 2915 21637
rect 3001 21581 3057 21637
rect 3143 21581 3199 21637
rect 3285 21581 3341 21637
rect 3427 21581 3483 21637
rect 3569 21581 3625 21637
rect 3711 21581 3767 21637
rect 3853 21581 3909 21637
rect 3995 21581 4051 21637
rect 4137 21581 4193 21637
rect 4279 21581 4335 21637
rect 4421 21581 4477 21637
rect 4563 21581 4619 21637
rect 4705 21581 4761 21637
rect 4847 21581 4903 21637
rect 4989 21581 5045 21637
rect 5131 21581 5187 21637
rect 5273 21581 5329 21637
rect 5415 21581 5471 21637
rect 5557 21581 5613 21637
rect 5699 21581 5755 21637
rect 5841 21581 5897 21637
rect 5983 21581 6039 21637
rect 6125 21581 6181 21637
rect 6267 21581 6323 21637
rect 6409 21581 6465 21637
rect 6551 21581 6607 21637
rect 6693 21581 6749 21637
rect 6835 21581 6891 21637
rect 6977 21581 7033 21637
rect 7119 21581 7175 21637
rect 7261 21581 7317 21637
rect 7403 21581 7459 21637
rect 7545 21581 7601 21637
rect 7687 21581 7743 21637
rect 7829 21581 7885 21637
rect 7971 21581 8027 21637
rect 8113 21581 8169 21637
rect 8255 21581 8311 21637
rect 8397 21581 8453 21637
rect 8539 21581 8595 21637
rect 8681 21581 8737 21637
rect 8823 21581 8879 21637
rect 8965 21581 9021 21637
rect 9107 21581 9163 21637
rect 9249 21581 9305 21637
rect 9391 21581 9447 21637
rect 9533 21581 9589 21637
rect 9675 21581 9731 21637
rect 9817 21581 9873 21637
rect 9959 21581 10015 21637
rect 10101 21581 10157 21637
rect 10243 21581 10299 21637
rect 10385 21581 10441 21637
rect 10527 21581 10583 21637
rect 10669 21581 10725 21637
rect 10811 21581 10867 21637
rect 10953 21581 11009 21637
rect 11095 21581 11151 21637
rect 11237 21581 11293 21637
rect 11379 21581 11435 21637
rect 11521 21581 11577 21637
rect 11663 21581 11719 21637
rect 11805 21581 11861 21637
rect 11947 21581 12003 21637
rect 12089 21581 12145 21637
rect 12231 21581 12287 21637
rect 12373 21581 12429 21637
rect 12515 21581 12571 21637
rect 12657 21581 12713 21637
rect 12799 21581 12855 21637
rect 12941 21581 12997 21637
rect 13083 21581 13139 21637
rect 13225 21581 13281 21637
rect 13367 21581 13423 21637
rect 13509 21581 13565 21637
rect 13651 21581 13707 21637
rect 13793 21581 13849 21637
rect 13935 21581 13991 21637
rect 14077 21581 14133 21637
rect 14219 21581 14275 21637
rect 14361 21581 14417 21637
rect 14503 21581 14559 21637
rect 14645 21581 14701 21637
rect 14787 21581 14843 21637
rect 161 21439 217 21495
rect 303 21439 359 21495
rect 445 21439 501 21495
rect 587 21439 643 21495
rect 729 21439 785 21495
rect 871 21439 927 21495
rect 1013 21439 1069 21495
rect 1155 21439 1211 21495
rect 1297 21439 1353 21495
rect 1439 21439 1495 21495
rect 1581 21439 1637 21495
rect 1723 21439 1779 21495
rect 1865 21439 1921 21495
rect 2007 21439 2063 21495
rect 2149 21439 2205 21495
rect 2291 21439 2347 21495
rect 2433 21439 2489 21495
rect 2575 21439 2631 21495
rect 2717 21439 2773 21495
rect 2859 21439 2915 21495
rect 3001 21439 3057 21495
rect 3143 21439 3199 21495
rect 3285 21439 3341 21495
rect 3427 21439 3483 21495
rect 3569 21439 3625 21495
rect 3711 21439 3767 21495
rect 3853 21439 3909 21495
rect 3995 21439 4051 21495
rect 4137 21439 4193 21495
rect 4279 21439 4335 21495
rect 4421 21439 4477 21495
rect 4563 21439 4619 21495
rect 4705 21439 4761 21495
rect 4847 21439 4903 21495
rect 4989 21439 5045 21495
rect 5131 21439 5187 21495
rect 5273 21439 5329 21495
rect 5415 21439 5471 21495
rect 5557 21439 5613 21495
rect 5699 21439 5755 21495
rect 5841 21439 5897 21495
rect 5983 21439 6039 21495
rect 6125 21439 6181 21495
rect 6267 21439 6323 21495
rect 6409 21439 6465 21495
rect 6551 21439 6607 21495
rect 6693 21439 6749 21495
rect 6835 21439 6891 21495
rect 6977 21439 7033 21495
rect 7119 21439 7175 21495
rect 7261 21439 7317 21495
rect 7403 21439 7459 21495
rect 7545 21439 7601 21495
rect 7687 21439 7743 21495
rect 7829 21439 7885 21495
rect 7971 21439 8027 21495
rect 8113 21439 8169 21495
rect 8255 21439 8311 21495
rect 8397 21439 8453 21495
rect 8539 21439 8595 21495
rect 8681 21439 8737 21495
rect 8823 21439 8879 21495
rect 8965 21439 9021 21495
rect 9107 21439 9163 21495
rect 9249 21439 9305 21495
rect 9391 21439 9447 21495
rect 9533 21439 9589 21495
rect 9675 21439 9731 21495
rect 9817 21439 9873 21495
rect 9959 21439 10015 21495
rect 10101 21439 10157 21495
rect 10243 21439 10299 21495
rect 10385 21439 10441 21495
rect 10527 21439 10583 21495
rect 10669 21439 10725 21495
rect 10811 21439 10867 21495
rect 10953 21439 11009 21495
rect 11095 21439 11151 21495
rect 11237 21439 11293 21495
rect 11379 21439 11435 21495
rect 11521 21439 11577 21495
rect 11663 21439 11719 21495
rect 11805 21439 11861 21495
rect 11947 21439 12003 21495
rect 12089 21439 12145 21495
rect 12231 21439 12287 21495
rect 12373 21439 12429 21495
rect 12515 21439 12571 21495
rect 12657 21439 12713 21495
rect 12799 21439 12855 21495
rect 12941 21439 12997 21495
rect 13083 21439 13139 21495
rect 13225 21439 13281 21495
rect 13367 21439 13423 21495
rect 13509 21439 13565 21495
rect 13651 21439 13707 21495
rect 13793 21439 13849 21495
rect 13935 21439 13991 21495
rect 14077 21439 14133 21495
rect 14219 21439 14275 21495
rect 14361 21439 14417 21495
rect 14503 21439 14559 21495
rect 14645 21439 14701 21495
rect 14787 21439 14843 21495
rect 161 21297 217 21353
rect 303 21297 359 21353
rect 445 21297 501 21353
rect 587 21297 643 21353
rect 729 21297 785 21353
rect 871 21297 927 21353
rect 1013 21297 1069 21353
rect 1155 21297 1211 21353
rect 1297 21297 1353 21353
rect 1439 21297 1495 21353
rect 1581 21297 1637 21353
rect 1723 21297 1779 21353
rect 1865 21297 1921 21353
rect 2007 21297 2063 21353
rect 2149 21297 2205 21353
rect 2291 21297 2347 21353
rect 2433 21297 2489 21353
rect 2575 21297 2631 21353
rect 2717 21297 2773 21353
rect 2859 21297 2915 21353
rect 3001 21297 3057 21353
rect 3143 21297 3199 21353
rect 3285 21297 3341 21353
rect 3427 21297 3483 21353
rect 3569 21297 3625 21353
rect 3711 21297 3767 21353
rect 3853 21297 3909 21353
rect 3995 21297 4051 21353
rect 4137 21297 4193 21353
rect 4279 21297 4335 21353
rect 4421 21297 4477 21353
rect 4563 21297 4619 21353
rect 4705 21297 4761 21353
rect 4847 21297 4903 21353
rect 4989 21297 5045 21353
rect 5131 21297 5187 21353
rect 5273 21297 5329 21353
rect 5415 21297 5471 21353
rect 5557 21297 5613 21353
rect 5699 21297 5755 21353
rect 5841 21297 5897 21353
rect 5983 21297 6039 21353
rect 6125 21297 6181 21353
rect 6267 21297 6323 21353
rect 6409 21297 6465 21353
rect 6551 21297 6607 21353
rect 6693 21297 6749 21353
rect 6835 21297 6891 21353
rect 6977 21297 7033 21353
rect 7119 21297 7175 21353
rect 7261 21297 7317 21353
rect 7403 21297 7459 21353
rect 7545 21297 7601 21353
rect 7687 21297 7743 21353
rect 7829 21297 7885 21353
rect 7971 21297 8027 21353
rect 8113 21297 8169 21353
rect 8255 21297 8311 21353
rect 8397 21297 8453 21353
rect 8539 21297 8595 21353
rect 8681 21297 8737 21353
rect 8823 21297 8879 21353
rect 8965 21297 9021 21353
rect 9107 21297 9163 21353
rect 9249 21297 9305 21353
rect 9391 21297 9447 21353
rect 9533 21297 9589 21353
rect 9675 21297 9731 21353
rect 9817 21297 9873 21353
rect 9959 21297 10015 21353
rect 10101 21297 10157 21353
rect 10243 21297 10299 21353
rect 10385 21297 10441 21353
rect 10527 21297 10583 21353
rect 10669 21297 10725 21353
rect 10811 21297 10867 21353
rect 10953 21297 11009 21353
rect 11095 21297 11151 21353
rect 11237 21297 11293 21353
rect 11379 21297 11435 21353
rect 11521 21297 11577 21353
rect 11663 21297 11719 21353
rect 11805 21297 11861 21353
rect 11947 21297 12003 21353
rect 12089 21297 12145 21353
rect 12231 21297 12287 21353
rect 12373 21297 12429 21353
rect 12515 21297 12571 21353
rect 12657 21297 12713 21353
rect 12799 21297 12855 21353
rect 12941 21297 12997 21353
rect 13083 21297 13139 21353
rect 13225 21297 13281 21353
rect 13367 21297 13423 21353
rect 13509 21297 13565 21353
rect 13651 21297 13707 21353
rect 13793 21297 13849 21353
rect 13935 21297 13991 21353
rect 14077 21297 14133 21353
rect 14219 21297 14275 21353
rect 14361 21297 14417 21353
rect 14503 21297 14559 21353
rect 14645 21297 14701 21353
rect 14787 21297 14843 21353
rect 161 21155 217 21211
rect 303 21155 359 21211
rect 445 21155 501 21211
rect 587 21155 643 21211
rect 729 21155 785 21211
rect 871 21155 927 21211
rect 1013 21155 1069 21211
rect 1155 21155 1211 21211
rect 1297 21155 1353 21211
rect 1439 21155 1495 21211
rect 1581 21155 1637 21211
rect 1723 21155 1779 21211
rect 1865 21155 1921 21211
rect 2007 21155 2063 21211
rect 2149 21155 2205 21211
rect 2291 21155 2347 21211
rect 2433 21155 2489 21211
rect 2575 21155 2631 21211
rect 2717 21155 2773 21211
rect 2859 21155 2915 21211
rect 3001 21155 3057 21211
rect 3143 21155 3199 21211
rect 3285 21155 3341 21211
rect 3427 21155 3483 21211
rect 3569 21155 3625 21211
rect 3711 21155 3767 21211
rect 3853 21155 3909 21211
rect 3995 21155 4051 21211
rect 4137 21155 4193 21211
rect 4279 21155 4335 21211
rect 4421 21155 4477 21211
rect 4563 21155 4619 21211
rect 4705 21155 4761 21211
rect 4847 21155 4903 21211
rect 4989 21155 5045 21211
rect 5131 21155 5187 21211
rect 5273 21155 5329 21211
rect 5415 21155 5471 21211
rect 5557 21155 5613 21211
rect 5699 21155 5755 21211
rect 5841 21155 5897 21211
rect 5983 21155 6039 21211
rect 6125 21155 6181 21211
rect 6267 21155 6323 21211
rect 6409 21155 6465 21211
rect 6551 21155 6607 21211
rect 6693 21155 6749 21211
rect 6835 21155 6891 21211
rect 6977 21155 7033 21211
rect 7119 21155 7175 21211
rect 7261 21155 7317 21211
rect 7403 21155 7459 21211
rect 7545 21155 7601 21211
rect 7687 21155 7743 21211
rect 7829 21155 7885 21211
rect 7971 21155 8027 21211
rect 8113 21155 8169 21211
rect 8255 21155 8311 21211
rect 8397 21155 8453 21211
rect 8539 21155 8595 21211
rect 8681 21155 8737 21211
rect 8823 21155 8879 21211
rect 8965 21155 9021 21211
rect 9107 21155 9163 21211
rect 9249 21155 9305 21211
rect 9391 21155 9447 21211
rect 9533 21155 9589 21211
rect 9675 21155 9731 21211
rect 9817 21155 9873 21211
rect 9959 21155 10015 21211
rect 10101 21155 10157 21211
rect 10243 21155 10299 21211
rect 10385 21155 10441 21211
rect 10527 21155 10583 21211
rect 10669 21155 10725 21211
rect 10811 21155 10867 21211
rect 10953 21155 11009 21211
rect 11095 21155 11151 21211
rect 11237 21155 11293 21211
rect 11379 21155 11435 21211
rect 11521 21155 11577 21211
rect 11663 21155 11719 21211
rect 11805 21155 11861 21211
rect 11947 21155 12003 21211
rect 12089 21155 12145 21211
rect 12231 21155 12287 21211
rect 12373 21155 12429 21211
rect 12515 21155 12571 21211
rect 12657 21155 12713 21211
rect 12799 21155 12855 21211
rect 12941 21155 12997 21211
rect 13083 21155 13139 21211
rect 13225 21155 13281 21211
rect 13367 21155 13423 21211
rect 13509 21155 13565 21211
rect 13651 21155 13707 21211
rect 13793 21155 13849 21211
rect 13935 21155 13991 21211
rect 14077 21155 14133 21211
rect 14219 21155 14275 21211
rect 14361 21155 14417 21211
rect 14503 21155 14559 21211
rect 14645 21155 14701 21211
rect 14787 21155 14843 21211
rect 161 21013 217 21069
rect 303 21013 359 21069
rect 445 21013 501 21069
rect 587 21013 643 21069
rect 729 21013 785 21069
rect 871 21013 927 21069
rect 1013 21013 1069 21069
rect 1155 21013 1211 21069
rect 1297 21013 1353 21069
rect 1439 21013 1495 21069
rect 1581 21013 1637 21069
rect 1723 21013 1779 21069
rect 1865 21013 1921 21069
rect 2007 21013 2063 21069
rect 2149 21013 2205 21069
rect 2291 21013 2347 21069
rect 2433 21013 2489 21069
rect 2575 21013 2631 21069
rect 2717 21013 2773 21069
rect 2859 21013 2915 21069
rect 3001 21013 3057 21069
rect 3143 21013 3199 21069
rect 3285 21013 3341 21069
rect 3427 21013 3483 21069
rect 3569 21013 3625 21069
rect 3711 21013 3767 21069
rect 3853 21013 3909 21069
rect 3995 21013 4051 21069
rect 4137 21013 4193 21069
rect 4279 21013 4335 21069
rect 4421 21013 4477 21069
rect 4563 21013 4619 21069
rect 4705 21013 4761 21069
rect 4847 21013 4903 21069
rect 4989 21013 5045 21069
rect 5131 21013 5187 21069
rect 5273 21013 5329 21069
rect 5415 21013 5471 21069
rect 5557 21013 5613 21069
rect 5699 21013 5755 21069
rect 5841 21013 5897 21069
rect 5983 21013 6039 21069
rect 6125 21013 6181 21069
rect 6267 21013 6323 21069
rect 6409 21013 6465 21069
rect 6551 21013 6607 21069
rect 6693 21013 6749 21069
rect 6835 21013 6891 21069
rect 6977 21013 7033 21069
rect 7119 21013 7175 21069
rect 7261 21013 7317 21069
rect 7403 21013 7459 21069
rect 7545 21013 7601 21069
rect 7687 21013 7743 21069
rect 7829 21013 7885 21069
rect 7971 21013 8027 21069
rect 8113 21013 8169 21069
rect 8255 21013 8311 21069
rect 8397 21013 8453 21069
rect 8539 21013 8595 21069
rect 8681 21013 8737 21069
rect 8823 21013 8879 21069
rect 8965 21013 9021 21069
rect 9107 21013 9163 21069
rect 9249 21013 9305 21069
rect 9391 21013 9447 21069
rect 9533 21013 9589 21069
rect 9675 21013 9731 21069
rect 9817 21013 9873 21069
rect 9959 21013 10015 21069
rect 10101 21013 10157 21069
rect 10243 21013 10299 21069
rect 10385 21013 10441 21069
rect 10527 21013 10583 21069
rect 10669 21013 10725 21069
rect 10811 21013 10867 21069
rect 10953 21013 11009 21069
rect 11095 21013 11151 21069
rect 11237 21013 11293 21069
rect 11379 21013 11435 21069
rect 11521 21013 11577 21069
rect 11663 21013 11719 21069
rect 11805 21013 11861 21069
rect 11947 21013 12003 21069
rect 12089 21013 12145 21069
rect 12231 21013 12287 21069
rect 12373 21013 12429 21069
rect 12515 21013 12571 21069
rect 12657 21013 12713 21069
rect 12799 21013 12855 21069
rect 12941 21013 12997 21069
rect 13083 21013 13139 21069
rect 13225 21013 13281 21069
rect 13367 21013 13423 21069
rect 13509 21013 13565 21069
rect 13651 21013 13707 21069
rect 13793 21013 13849 21069
rect 13935 21013 13991 21069
rect 14077 21013 14133 21069
rect 14219 21013 14275 21069
rect 14361 21013 14417 21069
rect 14503 21013 14559 21069
rect 14645 21013 14701 21069
rect 14787 21013 14843 21069
rect 161 20871 217 20927
rect 303 20871 359 20927
rect 445 20871 501 20927
rect 587 20871 643 20927
rect 729 20871 785 20927
rect 871 20871 927 20927
rect 1013 20871 1069 20927
rect 1155 20871 1211 20927
rect 1297 20871 1353 20927
rect 1439 20871 1495 20927
rect 1581 20871 1637 20927
rect 1723 20871 1779 20927
rect 1865 20871 1921 20927
rect 2007 20871 2063 20927
rect 2149 20871 2205 20927
rect 2291 20871 2347 20927
rect 2433 20871 2489 20927
rect 2575 20871 2631 20927
rect 2717 20871 2773 20927
rect 2859 20871 2915 20927
rect 3001 20871 3057 20927
rect 3143 20871 3199 20927
rect 3285 20871 3341 20927
rect 3427 20871 3483 20927
rect 3569 20871 3625 20927
rect 3711 20871 3767 20927
rect 3853 20871 3909 20927
rect 3995 20871 4051 20927
rect 4137 20871 4193 20927
rect 4279 20871 4335 20927
rect 4421 20871 4477 20927
rect 4563 20871 4619 20927
rect 4705 20871 4761 20927
rect 4847 20871 4903 20927
rect 4989 20871 5045 20927
rect 5131 20871 5187 20927
rect 5273 20871 5329 20927
rect 5415 20871 5471 20927
rect 5557 20871 5613 20927
rect 5699 20871 5755 20927
rect 5841 20871 5897 20927
rect 5983 20871 6039 20927
rect 6125 20871 6181 20927
rect 6267 20871 6323 20927
rect 6409 20871 6465 20927
rect 6551 20871 6607 20927
rect 6693 20871 6749 20927
rect 6835 20871 6891 20927
rect 6977 20871 7033 20927
rect 7119 20871 7175 20927
rect 7261 20871 7317 20927
rect 7403 20871 7459 20927
rect 7545 20871 7601 20927
rect 7687 20871 7743 20927
rect 7829 20871 7885 20927
rect 7971 20871 8027 20927
rect 8113 20871 8169 20927
rect 8255 20871 8311 20927
rect 8397 20871 8453 20927
rect 8539 20871 8595 20927
rect 8681 20871 8737 20927
rect 8823 20871 8879 20927
rect 8965 20871 9021 20927
rect 9107 20871 9163 20927
rect 9249 20871 9305 20927
rect 9391 20871 9447 20927
rect 9533 20871 9589 20927
rect 9675 20871 9731 20927
rect 9817 20871 9873 20927
rect 9959 20871 10015 20927
rect 10101 20871 10157 20927
rect 10243 20871 10299 20927
rect 10385 20871 10441 20927
rect 10527 20871 10583 20927
rect 10669 20871 10725 20927
rect 10811 20871 10867 20927
rect 10953 20871 11009 20927
rect 11095 20871 11151 20927
rect 11237 20871 11293 20927
rect 11379 20871 11435 20927
rect 11521 20871 11577 20927
rect 11663 20871 11719 20927
rect 11805 20871 11861 20927
rect 11947 20871 12003 20927
rect 12089 20871 12145 20927
rect 12231 20871 12287 20927
rect 12373 20871 12429 20927
rect 12515 20871 12571 20927
rect 12657 20871 12713 20927
rect 12799 20871 12855 20927
rect 12941 20871 12997 20927
rect 13083 20871 13139 20927
rect 13225 20871 13281 20927
rect 13367 20871 13423 20927
rect 13509 20871 13565 20927
rect 13651 20871 13707 20927
rect 13793 20871 13849 20927
rect 13935 20871 13991 20927
rect 14077 20871 14133 20927
rect 14219 20871 14275 20927
rect 14361 20871 14417 20927
rect 14503 20871 14559 20927
rect 14645 20871 14701 20927
rect 14787 20871 14843 20927
rect 161 20729 217 20785
rect 303 20729 359 20785
rect 445 20729 501 20785
rect 587 20729 643 20785
rect 729 20729 785 20785
rect 871 20729 927 20785
rect 1013 20729 1069 20785
rect 1155 20729 1211 20785
rect 1297 20729 1353 20785
rect 1439 20729 1495 20785
rect 1581 20729 1637 20785
rect 1723 20729 1779 20785
rect 1865 20729 1921 20785
rect 2007 20729 2063 20785
rect 2149 20729 2205 20785
rect 2291 20729 2347 20785
rect 2433 20729 2489 20785
rect 2575 20729 2631 20785
rect 2717 20729 2773 20785
rect 2859 20729 2915 20785
rect 3001 20729 3057 20785
rect 3143 20729 3199 20785
rect 3285 20729 3341 20785
rect 3427 20729 3483 20785
rect 3569 20729 3625 20785
rect 3711 20729 3767 20785
rect 3853 20729 3909 20785
rect 3995 20729 4051 20785
rect 4137 20729 4193 20785
rect 4279 20729 4335 20785
rect 4421 20729 4477 20785
rect 4563 20729 4619 20785
rect 4705 20729 4761 20785
rect 4847 20729 4903 20785
rect 4989 20729 5045 20785
rect 5131 20729 5187 20785
rect 5273 20729 5329 20785
rect 5415 20729 5471 20785
rect 5557 20729 5613 20785
rect 5699 20729 5755 20785
rect 5841 20729 5897 20785
rect 5983 20729 6039 20785
rect 6125 20729 6181 20785
rect 6267 20729 6323 20785
rect 6409 20729 6465 20785
rect 6551 20729 6607 20785
rect 6693 20729 6749 20785
rect 6835 20729 6891 20785
rect 6977 20729 7033 20785
rect 7119 20729 7175 20785
rect 7261 20729 7317 20785
rect 7403 20729 7459 20785
rect 7545 20729 7601 20785
rect 7687 20729 7743 20785
rect 7829 20729 7885 20785
rect 7971 20729 8027 20785
rect 8113 20729 8169 20785
rect 8255 20729 8311 20785
rect 8397 20729 8453 20785
rect 8539 20729 8595 20785
rect 8681 20729 8737 20785
rect 8823 20729 8879 20785
rect 8965 20729 9021 20785
rect 9107 20729 9163 20785
rect 9249 20729 9305 20785
rect 9391 20729 9447 20785
rect 9533 20729 9589 20785
rect 9675 20729 9731 20785
rect 9817 20729 9873 20785
rect 9959 20729 10015 20785
rect 10101 20729 10157 20785
rect 10243 20729 10299 20785
rect 10385 20729 10441 20785
rect 10527 20729 10583 20785
rect 10669 20729 10725 20785
rect 10811 20729 10867 20785
rect 10953 20729 11009 20785
rect 11095 20729 11151 20785
rect 11237 20729 11293 20785
rect 11379 20729 11435 20785
rect 11521 20729 11577 20785
rect 11663 20729 11719 20785
rect 11805 20729 11861 20785
rect 11947 20729 12003 20785
rect 12089 20729 12145 20785
rect 12231 20729 12287 20785
rect 12373 20729 12429 20785
rect 12515 20729 12571 20785
rect 12657 20729 12713 20785
rect 12799 20729 12855 20785
rect 12941 20729 12997 20785
rect 13083 20729 13139 20785
rect 13225 20729 13281 20785
rect 13367 20729 13423 20785
rect 13509 20729 13565 20785
rect 13651 20729 13707 20785
rect 13793 20729 13849 20785
rect 13935 20729 13991 20785
rect 14077 20729 14133 20785
rect 14219 20729 14275 20785
rect 14361 20729 14417 20785
rect 14503 20729 14559 20785
rect 14645 20729 14701 20785
rect 14787 20729 14843 20785
rect 161 20587 217 20643
rect 303 20587 359 20643
rect 445 20587 501 20643
rect 587 20587 643 20643
rect 729 20587 785 20643
rect 871 20587 927 20643
rect 1013 20587 1069 20643
rect 1155 20587 1211 20643
rect 1297 20587 1353 20643
rect 1439 20587 1495 20643
rect 1581 20587 1637 20643
rect 1723 20587 1779 20643
rect 1865 20587 1921 20643
rect 2007 20587 2063 20643
rect 2149 20587 2205 20643
rect 2291 20587 2347 20643
rect 2433 20587 2489 20643
rect 2575 20587 2631 20643
rect 2717 20587 2773 20643
rect 2859 20587 2915 20643
rect 3001 20587 3057 20643
rect 3143 20587 3199 20643
rect 3285 20587 3341 20643
rect 3427 20587 3483 20643
rect 3569 20587 3625 20643
rect 3711 20587 3767 20643
rect 3853 20587 3909 20643
rect 3995 20587 4051 20643
rect 4137 20587 4193 20643
rect 4279 20587 4335 20643
rect 4421 20587 4477 20643
rect 4563 20587 4619 20643
rect 4705 20587 4761 20643
rect 4847 20587 4903 20643
rect 4989 20587 5045 20643
rect 5131 20587 5187 20643
rect 5273 20587 5329 20643
rect 5415 20587 5471 20643
rect 5557 20587 5613 20643
rect 5699 20587 5755 20643
rect 5841 20587 5897 20643
rect 5983 20587 6039 20643
rect 6125 20587 6181 20643
rect 6267 20587 6323 20643
rect 6409 20587 6465 20643
rect 6551 20587 6607 20643
rect 6693 20587 6749 20643
rect 6835 20587 6891 20643
rect 6977 20587 7033 20643
rect 7119 20587 7175 20643
rect 7261 20587 7317 20643
rect 7403 20587 7459 20643
rect 7545 20587 7601 20643
rect 7687 20587 7743 20643
rect 7829 20587 7885 20643
rect 7971 20587 8027 20643
rect 8113 20587 8169 20643
rect 8255 20587 8311 20643
rect 8397 20587 8453 20643
rect 8539 20587 8595 20643
rect 8681 20587 8737 20643
rect 8823 20587 8879 20643
rect 8965 20587 9021 20643
rect 9107 20587 9163 20643
rect 9249 20587 9305 20643
rect 9391 20587 9447 20643
rect 9533 20587 9589 20643
rect 9675 20587 9731 20643
rect 9817 20587 9873 20643
rect 9959 20587 10015 20643
rect 10101 20587 10157 20643
rect 10243 20587 10299 20643
rect 10385 20587 10441 20643
rect 10527 20587 10583 20643
rect 10669 20587 10725 20643
rect 10811 20587 10867 20643
rect 10953 20587 11009 20643
rect 11095 20587 11151 20643
rect 11237 20587 11293 20643
rect 11379 20587 11435 20643
rect 11521 20587 11577 20643
rect 11663 20587 11719 20643
rect 11805 20587 11861 20643
rect 11947 20587 12003 20643
rect 12089 20587 12145 20643
rect 12231 20587 12287 20643
rect 12373 20587 12429 20643
rect 12515 20587 12571 20643
rect 12657 20587 12713 20643
rect 12799 20587 12855 20643
rect 12941 20587 12997 20643
rect 13083 20587 13139 20643
rect 13225 20587 13281 20643
rect 13367 20587 13423 20643
rect 13509 20587 13565 20643
rect 13651 20587 13707 20643
rect 13793 20587 13849 20643
rect 13935 20587 13991 20643
rect 14077 20587 14133 20643
rect 14219 20587 14275 20643
rect 14361 20587 14417 20643
rect 14503 20587 14559 20643
rect 14645 20587 14701 20643
rect 14787 20587 14843 20643
rect 161 20445 217 20501
rect 303 20445 359 20501
rect 445 20445 501 20501
rect 587 20445 643 20501
rect 729 20445 785 20501
rect 871 20445 927 20501
rect 1013 20445 1069 20501
rect 1155 20445 1211 20501
rect 1297 20445 1353 20501
rect 1439 20445 1495 20501
rect 1581 20445 1637 20501
rect 1723 20445 1779 20501
rect 1865 20445 1921 20501
rect 2007 20445 2063 20501
rect 2149 20445 2205 20501
rect 2291 20445 2347 20501
rect 2433 20445 2489 20501
rect 2575 20445 2631 20501
rect 2717 20445 2773 20501
rect 2859 20445 2915 20501
rect 3001 20445 3057 20501
rect 3143 20445 3199 20501
rect 3285 20445 3341 20501
rect 3427 20445 3483 20501
rect 3569 20445 3625 20501
rect 3711 20445 3767 20501
rect 3853 20445 3909 20501
rect 3995 20445 4051 20501
rect 4137 20445 4193 20501
rect 4279 20445 4335 20501
rect 4421 20445 4477 20501
rect 4563 20445 4619 20501
rect 4705 20445 4761 20501
rect 4847 20445 4903 20501
rect 4989 20445 5045 20501
rect 5131 20445 5187 20501
rect 5273 20445 5329 20501
rect 5415 20445 5471 20501
rect 5557 20445 5613 20501
rect 5699 20445 5755 20501
rect 5841 20445 5897 20501
rect 5983 20445 6039 20501
rect 6125 20445 6181 20501
rect 6267 20445 6323 20501
rect 6409 20445 6465 20501
rect 6551 20445 6607 20501
rect 6693 20445 6749 20501
rect 6835 20445 6891 20501
rect 6977 20445 7033 20501
rect 7119 20445 7175 20501
rect 7261 20445 7317 20501
rect 7403 20445 7459 20501
rect 7545 20445 7601 20501
rect 7687 20445 7743 20501
rect 7829 20445 7885 20501
rect 7971 20445 8027 20501
rect 8113 20445 8169 20501
rect 8255 20445 8311 20501
rect 8397 20445 8453 20501
rect 8539 20445 8595 20501
rect 8681 20445 8737 20501
rect 8823 20445 8879 20501
rect 8965 20445 9021 20501
rect 9107 20445 9163 20501
rect 9249 20445 9305 20501
rect 9391 20445 9447 20501
rect 9533 20445 9589 20501
rect 9675 20445 9731 20501
rect 9817 20445 9873 20501
rect 9959 20445 10015 20501
rect 10101 20445 10157 20501
rect 10243 20445 10299 20501
rect 10385 20445 10441 20501
rect 10527 20445 10583 20501
rect 10669 20445 10725 20501
rect 10811 20445 10867 20501
rect 10953 20445 11009 20501
rect 11095 20445 11151 20501
rect 11237 20445 11293 20501
rect 11379 20445 11435 20501
rect 11521 20445 11577 20501
rect 11663 20445 11719 20501
rect 11805 20445 11861 20501
rect 11947 20445 12003 20501
rect 12089 20445 12145 20501
rect 12231 20445 12287 20501
rect 12373 20445 12429 20501
rect 12515 20445 12571 20501
rect 12657 20445 12713 20501
rect 12799 20445 12855 20501
rect 12941 20445 12997 20501
rect 13083 20445 13139 20501
rect 13225 20445 13281 20501
rect 13367 20445 13423 20501
rect 13509 20445 13565 20501
rect 13651 20445 13707 20501
rect 13793 20445 13849 20501
rect 13935 20445 13991 20501
rect 14077 20445 14133 20501
rect 14219 20445 14275 20501
rect 14361 20445 14417 20501
rect 14503 20445 14559 20501
rect 14645 20445 14701 20501
rect 14787 20445 14843 20501
rect 161 20085 217 20141
rect 303 20085 359 20141
rect 445 20085 501 20141
rect 587 20085 643 20141
rect 729 20085 785 20141
rect 871 20085 927 20141
rect 1013 20085 1069 20141
rect 1155 20085 1211 20141
rect 1297 20085 1353 20141
rect 1439 20085 1495 20141
rect 1581 20085 1637 20141
rect 1723 20085 1779 20141
rect 1865 20085 1921 20141
rect 2007 20085 2063 20141
rect 2149 20085 2205 20141
rect 2291 20085 2347 20141
rect 2433 20085 2489 20141
rect 2575 20085 2631 20141
rect 2717 20085 2773 20141
rect 2859 20085 2915 20141
rect 3001 20085 3057 20141
rect 3143 20085 3199 20141
rect 3285 20085 3341 20141
rect 3427 20085 3483 20141
rect 3569 20085 3625 20141
rect 3711 20085 3767 20141
rect 3853 20085 3909 20141
rect 3995 20085 4051 20141
rect 4137 20085 4193 20141
rect 4279 20085 4335 20141
rect 4421 20085 4477 20141
rect 4563 20085 4619 20141
rect 4705 20085 4761 20141
rect 4847 20085 4903 20141
rect 4989 20085 5045 20141
rect 5131 20085 5187 20141
rect 5273 20085 5329 20141
rect 5415 20085 5471 20141
rect 5557 20085 5613 20141
rect 5699 20085 5755 20141
rect 5841 20085 5897 20141
rect 5983 20085 6039 20141
rect 6125 20085 6181 20141
rect 6267 20085 6323 20141
rect 6409 20085 6465 20141
rect 6551 20085 6607 20141
rect 6693 20085 6749 20141
rect 6835 20085 6891 20141
rect 6977 20085 7033 20141
rect 7119 20085 7175 20141
rect 7261 20085 7317 20141
rect 7403 20085 7459 20141
rect 7545 20085 7601 20141
rect 7687 20085 7743 20141
rect 7829 20085 7885 20141
rect 7971 20085 8027 20141
rect 8113 20085 8169 20141
rect 8255 20085 8311 20141
rect 8397 20085 8453 20141
rect 8539 20085 8595 20141
rect 8681 20085 8737 20141
rect 8823 20085 8879 20141
rect 8965 20085 9021 20141
rect 9107 20085 9163 20141
rect 9249 20085 9305 20141
rect 9391 20085 9447 20141
rect 9533 20085 9589 20141
rect 9675 20085 9731 20141
rect 9817 20085 9873 20141
rect 9959 20085 10015 20141
rect 10101 20085 10157 20141
rect 10243 20085 10299 20141
rect 10385 20085 10441 20141
rect 10527 20085 10583 20141
rect 10669 20085 10725 20141
rect 10811 20085 10867 20141
rect 10953 20085 11009 20141
rect 11095 20085 11151 20141
rect 11237 20085 11293 20141
rect 11379 20085 11435 20141
rect 11521 20085 11577 20141
rect 11663 20085 11719 20141
rect 11805 20085 11861 20141
rect 11947 20085 12003 20141
rect 12089 20085 12145 20141
rect 12231 20085 12287 20141
rect 12373 20085 12429 20141
rect 12515 20085 12571 20141
rect 12657 20085 12713 20141
rect 12799 20085 12855 20141
rect 12941 20085 12997 20141
rect 13083 20085 13139 20141
rect 13225 20085 13281 20141
rect 13367 20085 13423 20141
rect 13509 20085 13565 20141
rect 13651 20085 13707 20141
rect 13793 20085 13849 20141
rect 13935 20085 13991 20141
rect 14077 20085 14133 20141
rect 14219 20085 14275 20141
rect 14361 20085 14417 20141
rect 14503 20085 14559 20141
rect 14645 20085 14701 20141
rect 14787 20085 14843 20141
rect 161 19943 217 19999
rect 303 19943 359 19999
rect 445 19943 501 19999
rect 587 19943 643 19999
rect 729 19943 785 19999
rect 871 19943 927 19999
rect 1013 19943 1069 19999
rect 1155 19943 1211 19999
rect 1297 19943 1353 19999
rect 1439 19943 1495 19999
rect 1581 19943 1637 19999
rect 1723 19943 1779 19999
rect 1865 19943 1921 19999
rect 2007 19943 2063 19999
rect 2149 19943 2205 19999
rect 2291 19943 2347 19999
rect 2433 19943 2489 19999
rect 2575 19943 2631 19999
rect 2717 19943 2773 19999
rect 2859 19943 2915 19999
rect 3001 19943 3057 19999
rect 3143 19943 3199 19999
rect 3285 19943 3341 19999
rect 3427 19943 3483 19999
rect 3569 19943 3625 19999
rect 3711 19943 3767 19999
rect 3853 19943 3909 19999
rect 3995 19943 4051 19999
rect 4137 19943 4193 19999
rect 4279 19943 4335 19999
rect 4421 19943 4477 19999
rect 4563 19943 4619 19999
rect 4705 19943 4761 19999
rect 4847 19943 4903 19999
rect 4989 19943 5045 19999
rect 5131 19943 5187 19999
rect 5273 19943 5329 19999
rect 5415 19943 5471 19999
rect 5557 19943 5613 19999
rect 5699 19943 5755 19999
rect 5841 19943 5897 19999
rect 5983 19943 6039 19999
rect 6125 19943 6181 19999
rect 6267 19943 6323 19999
rect 6409 19943 6465 19999
rect 6551 19943 6607 19999
rect 6693 19943 6749 19999
rect 6835 19943 6891 19999
rect 6977 19943 7033 19999
rect 7119 19943 7175 19999
rect 7261 19943 7317 19999
rect 7403 19943 7459 19999
rect 7545 19943 7601 19999
rect 7687 19943 7743 19999
rect 7829 19943 7885 19999
rect 7971 19943 8027 19999
rect 8113 19943 8169 19999
rect 8255 19943 8311 19999
rect 8397 19943 8453 19999
rect 8539 19943 8595 19999
rect 8681 19943 8737 19999
rect 8823 19943 8879 19999
rect 8965 19943 9021 19999
rect 9107 19943 9163 19999
rect 9249 19943 9305 19999
rect 9391 19943 9447 19999
rect 9533 19943 9589 19999
rect 9675 19943 9731 19999
rect 9817 19943 9873 19999
rect 9959 19943 10015 19999
rect 10101 19943 10157 19999
rect 10243 19943 10299 19999
rect 10385 19943 10441 19999
rect 10527 19943 10583 19999
rect 10669 19943 10725 19999
rect 10811 19943 10867 19999
rect 10953 19943 11009 19999
rect 11095 19943 11151 19999
rect 11237 19943 11293 19999
rect 11379 19943 11435 19999
rect 11521 19943 11577 19999
rect 11663 19943 11719 19999
rect 11805 19943 11861 19999
rect 11947 19943 12003 19999
rect 12089 19943 12145 19999
rect 12231 19943 12287 19999
rect 12373 19943 12429 19999
rect 12515 19943 12571 19999
rect 12657 19943 12713 19999
rect 12799 19943 12855 19999
rect 12941 19943 12997 19999
rect 13083 19943 13139 19999
rect 13225 19943 13281 19999
rect 13367 19943 13423 19999
rect 13509 19943 13565 19999
rect 13651 19943 13707 19999
rect 13793 19943 13849 19999
rect 13935 19943 13991 19999
rect 14077 19943 14133 19999
rect 14219 19943 14275 19999
rect 14361 19943 14417 19999
rect 14503 19943 14559 19999
rect 14645 19943 14701 19999
rect 14787 19943 14843 19999
rect 161 19801 217 19857
rect 303 19801 359 19857
rect 445 19801 501 19857
rect 587 19801 643 19857
rect 729 19801 785 19857
rect 871 19801 927 19857
rect 1013 19801 1069 19857
rect 1155 19801 1211 19857
rect 1297 19801 1353 19857
rect 1439 19801 1495 19857
rect 1581 19801 1637 19857
rect 1723 19801 1779 19857
rect 1865 19801 1921 19857
rect 2007 19801 2063 19857
rect 2149 19801 2205 19857
rect 2291 19801 2347 19857
rect 2433 19801 2489 19857
rect 2575 19801 2631 19857
rect 2717 19801 2773 19857
rect 2859 19801 2915 19857
rect 3001 19801 3057 19857
rect 3143 19801 3199 19857
rect 3285 19801 3341 19857
rect 3427 19801 3483 19857
rect 3569 19801 3625 19857
rect 3711 19801 3767 19857
rect 3853 19801 3909 19857
rect 3995 19801 4051 19857
rect 4137 19801 4193 19857
rect 4279 19801 4335 19857
rect 4421 19801 4477 19857
rect 4563 19801 4619 19857
rect 4705 19801 4761 19857
rect 4847 19801 4903 19857
rect 4989 19801 5045 19857
rect 5131 19801 5187 19857
rect 5273 19801 5329 19857
rect 5415 19801 5471 19857
rect 5557 19801 5613 19857
rect 5699 19801 5755 19857
rect 5841 19801 5897 19857
rect 5983 19801 6039 19857
rect 6125 19801 6181 19857
rect 6267 19801 6323 19857
rect 6409 19801 6465 19857
rect 6551 19801 6607 19857
rect 6693 19801 6749 19857
rect 6835 19801 6891 19857
rect 6977 19801 7033 19857
rect 7119 19801 7175 19857
rect 7261 19801 7317 19857
rect 7403 19801 7459 19857
rect 7545 19801 7601 19857
rect 7687 19801 7743 19857
rect 7829 19801 7885 19857
rect 7971 19801 8027 19857
rect 8113 19801 8169 19857
rect 8255 19801 8311 19857
rect 8397 19801 8453 19857
rect 8539 19801 8595 19857
rect 8681 19801 8737 19857
rect 8823 19801 8879 19857
rect 8965 19801 9021 19857
rect 9107 19801 9163 19857
rect 9249 19801 9305 19857
rect 9391 19801 9447 19857
rect 9533 19801 9589 19857
rect 9675 19801 9731 19857
rect 9817 19801 9873 19857
rect 9959 19801 10015 19857
rect 10101 19801 10157 19857
rect 10243 19801 10299 19857
rect 10385 19801 10441 19857
rect 10527 19801 10583 19857
rect 10669 19801 10725 19857
rect 10811 19801 10867 19857
rect 10953 19801 11009 19857
rect 11095 19801 11151 19857
rect 11237 19801 11293 19857
rect 11379 19801 11435 19857
rect 11521 19801 11577 19857
rect 11663 19801 11719 19857
rect 11805 19801 11861 19857
rect 11947 19801 12003 19857
rect 12089 19801 12145 19857
rect 12231 19801 12287 19857
rect 12373 19801 12429 19857
rect 12515 19801 12571 19857
rect 12657 19801 12713 19857
rect 12799 19801 12855 19857
rect 12941 19801 12997 19857
rect 13083 19801 13139 19857
rect 13225 19801 13281 19857
rect 13367 19801 13423 19857
rect 13509 19801 13565 19857
rect 13651 19801 13707 19857
rect 13793 19801 13849 19857
rect 13935 19801 13991 19857
rect 14077 19801 14133 19857
rect 14219 19801 14275 19857
rect 14361 19801 14417 19857
rect 14503 19801 14559 19857
rect 14645 19801 14701 19857
rect 14787 19801 14843 19857
rect 161 19659 217 19715
rect 303 19659 359 19715
rect 445 19659 501 19715
rect 587 19659 643 19715
rect 729 19659 785 19715
rect 871 19659 927 19715
rect 1013 19659 1069 19715
rect 1155 19659 1211 19715
rect 1297 19659 1353 19715
rect 1439 19659 1495 19715
rect 1581 19659 1637 19715
rect 1723 19659 1779 19715
rect 1865 19659 1921 19715
rect 2007 19659 2063 19715
rect 2149 19659 2205 19715
rect 2291 19659 2347 19715
rect 2433 19659 2489 19715
rect 2575 19659 2631 19715
rect 2717 19659 2773 19715
rect 2859 19659 2915 19715
rect 3001 19659 3057 19715
rect 3143 19659 3199 19715
rect 3285 19659 3341 19715
rect 3427 19659 3483 19715
rect 3569 19659 3625 19715
rect 3711 19659 3767 19715
rect 3853 19659 3909 19715
rect 3995 19659 4051 19715
rect 4137 19659 4193 19715
rect 4279 19659 4335 19715
rect 4421 19659 4477 19715
rect 4563 19659 4619 19715
rect 4705 19659 4761 19715
rect 4847 19659 4903 19715
rect 4989 19659 5045 19715
rect 5131 19659 5187 19715
rect 5273 19659 5329 19715
rect 5415 19659 5471 19715
rect 5557 19659 5613 19715
rect 5699 19659 5755 19715
rect 5841 19659 5897 19715
rect 5983 19659 6039 19715
rect 6125 19659 6181 19715
rect 6267 19659 6323 19715
rect 6409 19659 6465 19715
rect 6551 19659 6607 19715
rect 6693 19659 6749 19715
rect 6835 19659 6891 19715
rect 6977 19659 7033 19715
rect 7119 19659 7175 19715
rect 7261 19659 7317 19715
rect 7403 19659 7459 19715
rect 7545 19659 7601 19715
rect 7687 19659 7743 19715
rect 7829 19659 7885 19715
rect 7971 19659 8027 19715
rect 8113 19659 8169 19715
rect 8255 19659 8311 19715
rect 8397 19659 8453 19715
rect 8539 19659 8595 19715
rect 8681 19659 8737 19715
rect 8823 19659 8879 19715
rect 8965 19659 9021 19715
rect 9107 19659 9163 19715
rect 9249 19659 9305 19715
rect 9391 19659 9447 19715
rect 9533 19659 9589 19715
rect 9675 19659 9731 19715
rect 9817 19659 9873 19715
rect 9959 19659 10015 19715
rect 10101 19659 10157 19715
rect 10243 19659 10299 19715
rect 10385 19659 10441 19715
rect 10527 19659 10583 19715
rect 10669 19659 10725 19715
rect 10811 19659 10867 19715
rect 10953 19659 11009 19715
rect 11095 19659 11151 19715
rect 11237 19659 11293 19715
rect 11379 19659 11435 19715
rect 11521 19659 11577 19715
rect 11663 19659 11719 19715
rect 11805 19659 11861 19715
rect 11947 19659 12003 19715
rect 12089 19659 12145 19715
rect 12231 19659 12287 19715
rect 12373 19659 12429 19715
rect 12515 19659 12571 19715
rect 12657 19659 12713 19715
rect 12799 19659 12855 19715
rect 12941 19659 12997 19715
rect 13083 19659 13139 19715
rect 13225 19659 13281 19715
rect 13367 19659 13423 19715
rect 13509 19659 13565 19715
rect 13651 19659 13707 19715
rect 13793 19659 13849 19715
rect 13935 19659 13991 19715
rect 14077 19659 14133 19715
rect 14219 19659 14275 19715
rect 14361 19659 14417 19715
rect 14503 19659 14559 19715
rect 14645 19659 14701 19715
rect 14787 19659 14843 19715
rect 161 19517 217 19573
rect 303 19517 359 19573
rect 445 19517 501 19573
rect 587 19517 643 19573
rect 729 19517 785 19573
rect 871 19517 927 19573
rect 1013 19517 1069 19573
rect 1155 19517 1211 19573
rect 1297 19517 1353 19573
rect 1439 19517 1495 19573
rect 1581 19517 1637 19573
rect 1723 19517 1779 19573
rect 1865 19517 1921 19573
rect 2007 19517 2063 19573
rect 2149 19517 2205 19573
rect 2291 19517 2347 19573
rect 2433 19517 2489 19573
rect 2575 19517 2631 19573
rect 2717 19517 2773 19573
rect 2859 19517 2915 19573
rect 3001 19517 3057 19573
rect 3143 19517 3199 19573
rect 3285 19517 3341 19573
rect 3427 19517 3483 19573
rect 3569 19517 3625 19573
rect 3711 19517 3767 19573
rect 3853 19517 3909 19573
rect 3995 19517 4051 19573
rect 4137 19517 4193 19573
rect 4279 19517 4335 19573
rect 4421 19517 4477 19573
rect 4563 19517 4619 19573
rect 4705 19517 4761 19573
rect 4847 19517 4903 19573
rect 4989 19517 5045 19573
rect 5131 19517 5187 19573
rect 5273 19517 5329 19573
rect 5415 19517 5471 19573
rect 5557 19517 5613 19573
rect 5699 19517 5755 19573
rect 5841 19517 5897 19573
rect 5983 19517 6039 19573
rect 6125 19517 6181 19573
rect 6267 19517 6323 19573
rect 6409 19517 6465 19573
rect 6551 19517 6607 19573
rect 6693 19517 6749 19573
rect 6835 19517 6891 19573
rect 6977 19517 7033 19573
rect 7119 19517 7175 19573
rect 7261 19517 7317 19573
rect 7403 19517 7459 19573
rect 7545 19517 7601 19573
rect 7687 19517 7743 19573
rect 7829 19517 7885 19573
rect 7971 19517 8027 19573
rect 8113 19517 8169 19573
rect 8255 19517 8311 19573
rect 8397 19517 8453 19573
rect 8539 19517 8595 19573
rect 8681 19517 8737 19573
rect 8823 19517 8879 19573
rect 8965 19517 9021 19573
rect 9107 19517 9163 19573
rect 9249 19517 9305 19573
rect 9391 19517 9447 19573
rect 9533 19517 9589 19573
rect 9675 19517 9731 19573
rect 9817 19517 9873 19573
rect 9959 19517 10015 19573
rect 10101 19517 10157 19573
rect 10243 19517 10299 19573
rect 10385 19517 10441 19573
rect 10527 19517 10583 19573
rect 10669 19517 10725 19573
rect 10811 19517 10867 19573
rect 10953 19517 11009 19573
rect 11095 19517 11151 19573
rect 11237 19517 11293 19573
rect 11379 19517 11435 19573
rect 11521 19517 11577 19573
rect 11663 19517 11719 19573
rect 11805 19517 11861 19573
rect 11947 19517 12003 19573
rect 12089 19517 12145 19573
rect 12231 19517 12287 19573
rect 12373 19517 12429 19573
rect 12515 19517 12571 19573
rect 12657 19517 12713 19573
rect 12799 19517 12855 19573
rect 12941 19517 12997 19573
rect 13083 19517 13139 19573
rect 13225 19517 13281 19573
rect 13367 19517 13423 19573
rect 13509 19517 13565 19573
rect 13651 19517 13707 19573
rect 13793 19517 13849 19573
rect 13935 19517 13991 19573
rect 14077 19517 14133 19573
rect 14219 19517 14275 19573
rect 14361 19517 14417 19573
rect 14503 19517 14559 19573
rect 14645 19517 14701 19573
rect 14787 19517 14843 19573
rect 161 19375 217 19431
rect 303 19375 359 19431
rect 445 19375 501 19431
rect 587 19375 643 19431
rect 729 19375 785 19431
rect 871 19375 927 19431
rect 1013 19375 1069 19431
rect 1155 19375 1211 19431
rect 1297 19375 1353 19431
rect 1439 19375 1495 19431
rect 1581 19375 1637 19431
rect 1723 19375 1779 19431
rect 1865 19375 1921 19431
rect 2007 19375 2063 19431
rect 2149 19375 2205 19431
rect 2291 19375 2347 19431
rect 2433 19375 2489 19431
rect 2575 19375 2631 19431
rect 2717 19375 2773 19431
rect 2859 19375 2915 19431
rect 3001 19375 3057 19431
rect 3143 19375 3199 19431
rect 3285 19375 3341 19431
rect 3427 19375 3483 19431
rect 3569 19375 3625 19431
rect 3711 19375 3767 19431
rect 3853 19375 3909 19431
rect 3995 19375 4051 19431
rect 4137 19375 4193 19431
rect 4279 19375 4335 19431
rect 4421 19375 4477 19431
rect 4563 19375 4619 19431
rect 4705 19375 4761 19431
rect 4847 19375 4903 19431
rect 4989 19375 5045 19431
rect 5131 19375 5187 19431
rect 5273 19375 5329 19431
rect 5415 19375 5471 19431
rect 5557 19375 5613 19431
rect 5699 19375 5755 19431
rect 5841 19375 5897 19431
rect 5983 19375 6039 19431
rect 6125 19375 6181 19431
rect 6267 19375 6323 19431
rect 6409 19375 6465 19431
rect 6551 19375 6607 19431
rect 6693 19375 6749 19431
rect 6835 19375 6891 19431
rect 6977 19375 7033 19431
rect 7119 19375 7175 19431
rect 7261 19375 7317 19431
rect 7403 19375 7459 19431
rect 7545 19375 7601 19431
rect 7687 19375 7743 19431
rect 7829 19375 7885 19431
rect 7971 19375 8027 19431
rect 8113 19375 8169 19431
rect 8255 19375 8311 19431
rect 8397 19375 8453 19431
rect 8539 19375 8595 19431
rect 8681 19375 8737 19431
rect 8823 19375 8879 19431
rect 8965 19375 9021 19431
rect 9107 19375 9163 19431
rect 9249 19375 9305 19431
rect 9391 19375 9447 19431
rect 9533 19375 9589 19431
rect 9675 19375 9731 19431
rect 9817 19375 9873 19431
rect 9959 19375 10015 19431
rect 10101 19375 10157 19431
rect 10243 19375 10299 19431
rect 10385 19375 10441 19431
rect 10527 19375 10583 19431
rect 10669 19375 10725 19431
rect 10811 19375 10867 19431
rect 10953 19375 11009 19431
rect 11095 19375 11151 19431
rect 11237 19375 11293 19431
rect 11379 19375 11435 19431
rect 11521 19375 11577 19431
rect 11663 19375 11719 19431
rect 11805 19375 11861 19431
rect 11947 19375 12003 19431
rect 12089 19375 12145 19431
rect 12231 19375 12287 19431
rect 12373 19375 12429 19431
rect 12515 19375 12571 19431
rect 12657 19375 12713 19431
rect 12799 19375 12855 19431
rect 12941 19375 12997 19431
rect 13083 19375 13139 19431
rect 13225 19375 13281 19431
rect 13367 19375 13423 19431
rect 13509 19375 13565 19431
rect 13651 19375 13707 19431
rect 13793 19375 13849 19431
rect 13935 19375 13991 19431
rect 14077 19375 14133 19431
rect 14219 19375 14275 19431
rect 14361 19375 14417 19431
rect 14503 19375 14559 19431
rect 14645 19375 14701 19431
rect 14787 19375 14843 19431
rect 161 19233 217 19289
rect 303 19233 359 19289
rect 445 19233 501 19289
rect 587 19233 643 19289
rect 729 19233 785 19289
rect 871 19233 927 19289
rect 1013 19233 1069 19289
rect 1155 19233 1211 19289
rect 1297 19233 1353 19289
rect 1439 19233 1495 19289
rect 1581 19233 1637 19289
rect 1723 19233 1779 19289
rect 1865 19233 1921 19289
rect 2007 19233 2063 19289
rect 2149 19233 2205 19289
rect 2291 19233 2347 19289
rect 2433 19233 2489 19289
rect 2575 19233 2631 19289
rect 2717 19233 2773 19289
rect 2859 19233 2915 19289
rect 3001 19233 3057 19289
rect 3143 19233 3199 19289
rect 3285 19233 3341 19289
rect 3427 19233 3483 19289
rect 3569 19233 3625 19289
rect 3711 19233 3767 19289
rect 3853 19233 3909 19289
rect 3995 19233 4051 19289
rect 4137 19233 4193 19289
rect 4279 19233 4335 19289
rect 4421 19233 4477 19289
rect 4563 19233 4619 19289
rect 4705 19233 4761 19289
rect 4847 19233 4903 19289
rect 4989 19233 5045 19289
rect 5131 19233 5187 19289
rect 5273 19233 5329 19289
rect 5415 19233 5471 19289
rect 5557 19233 5613 19289
rect 5699 19233 5755 19289
rect 5841 19233 5897 19289
rect 5983 19233 6039 19289
rect 6125 19233 6181 19289
rect 6267 19233 6323 19289
rect 6409 19233 6465 19289
rect 6551 19233 6607 19289
rect 6693 19233 6749 19289
rect 6835 19233 6891 19289
rect 6977 19233 7033 19289
rect 7119 19233 7175 19289
rect 7261 19233 7317 19289
rect 7403 19233 7459 19289
rect 7545 19233 7601 19289
rect 7687 19233 7743 19289
rect 7829 19233 7885 19289
rect 7971 19233 8027 19289
rect 8113 19233 8169 19289
rect 8255 19233 8311 19289
rect 8397 19233 8453 19289
rect 8539 19233 8595 19289
rect 8681 19233 8737 19289
rect 8823 19233 8879 19289
rect 8965 19233 9021 19289
rect 9107 19233 9163 19289
rect 9249 19233 9305 19289
rect 9391 19233 9447 19289
rect 9533 19233 9589 19289
rect 9675 19233 9731 19289
rect 9817 19233 9873 19289
rect 9959 19233 10015 19289
rect 10101 19233 10157 19289
rect 10243 19233 10299 19289
rect 10385 19233 10441 19289
rect 10527 19233 10583 19289
rect 10669 19233 10725 19289
rect 10811 19233 10867 19289
rect 10953 19233 11009 19289
rect 11095 19233 11151 19289
rect 11237 19233 11293 19289
rect 11379 19233 11435 19289
rect 11521 19233 11577 19289
rect 11663 19233 11719 19289
rect 11805 19233 11861 19289
rect 11947 19233 12003 19289
rect 12089 19233 12145 19289
rect 12231 19233 12287 19289
rect 12373 19233 12429 19289
rect 12515 19233 12571 19289
rect 12657 19233 12713 19289
rect 12799 19233 12855 19289
rect 12941 19233 12997 19289
rect 13083 19233 13139 19289
rect 13225 19233 13281 19289
rect 13367 19233 13423 19289
rect 13509 19233 13565 19289
rect 13651 19233 13707 19289
rect 13793 19233 13849 19289
rect 13935 19233 13991 19289
rect 14077 19233 14133 19289
rect 14219 19233 14275 19289
rect 14361 19233 14417 19289
rect 14503 19233 14559 19289
rect 14645 19233 14701 19289
rect 14787 19233 14843 19289
rect 161 19091 217 19147
rect 303 19091 359 19147
rect 445 19091 501 19147
rect 587 19091 643 19147
rect 729 19091 785 19147
rect 871 19091 927 19147
rect 1013 19091 1069 19147
rect 1155 19091 1211 19147
rect 1297 19091 1353 19147
rect 1439 19091 1495 19147
rect 1581 19091 1637 19147
rect 1723 19091 1779 19147
rect 1865 19091 1921 19147
rect 2007 19091 2063 19147
rect 2149 19091 2205 19147
rect 2291 19091 2347 19147
rect 2433 19091 2489 19147
rect 2575 19091 2631 19147
rect 2717 19091 2773 19147
rect 2859 19091 2915 19147
rect 3001 19091 3057 19147
rect 3143 19091 3199 19147
rect 3285 19091 3341 19147
rect 3427 19091 3483 19147
rect 3569 19091 3625 19147
rect 3711 19091 3767 19147
rect 3853 19091 3909 19147
rect 3995 19091 4051 19147
rect 4137 19091 4193 19147
rect 4279 19091 4335 19147
rect 4421 19091 4477 19147
rect 4563 19091 4619 19147
rect 4705 19091 4761 19147
rect 4847 19091 4903 19147
rect 4989 19091 5045 19147
rect 5131 19091 5187 19147
rect 5273 19091 5329 19147
rect 5415 19091 5471 19147
rect 5557 19091 5613 19147
rect 5699 19091 5755 19147
rect 5841 19091 5897 19147
rect 5983 19091 6039 19147
rect 6125 19091 6181 19147
rect 6267 19091 6323 19147
rect 6409 19091 6465 19147
rect 6551 19091 6607 19147
rect 6693 19091 6749 19147
rect 6835 19091 6891 19147
rect 6977 19091 7033 19147
rect 7119 19091 7175 19147
rect 7261 19091 7317 19147
rect 7403 19091 7459 19147
rect 7545 19091 7601 19147
rect 7687 19091 7743 19147
rect 7829 19091 7885 19147
rect 7971 19091 8027 19147
rect 8113 19091 8169 19147
rect 8255 19091 8311 19147
rect 8397 19091 8453 19147
rect 8539 19091 8595 19147
rect 8681 19091 8737 19147
rect 8823 19091 8879 19147
rect 8965 19091 9021 19147
rect 9107 19091 9163 19147
rect 9249 19091 9305 19147
rect 9391 19091 9447 19147
rect 9533 19091 9589 19147
rect 9675 19091 9731 19147
rect 9817 19091 9873 19147
rect 9959 19091 10015 19147
rect 10101 19091 10157 19147
rect 10243 19091 10299 19147
rect 10385 19091 10441 19147
rect 10527 19091 10583 19147
rect 10669 19091 10725 19147
rect 10811 19091 10867 19147
rect 10953 19091 11009 19147
rect 11095 19091 11151 19147
rect 11237 19091 11293 19147
rect 11379 19091 11435 19147
rect 11521 19091 11577 19147
rect 11663 19091 11719 19147
rect 11805 19091 11861 19147
rect 11947 19091 12003 19147
rect 12089 19091 12145 19147
rect 12231 19091 12287 19147
rect 12373 19091 12429 19147
rect 12515 19091 12571 19147
rect 12657 19091 12713 19147
rect 12799 19091 12855 19147
rect 12941 19091 12997 19147
rect 13083 19091 13139 19147
rect 13225 19091 13281 19147
rect 13367 19091 13423 19147
rect 13509 19091 13565 19147
rect 13651 19091 13707 19147
rect 13793 19091 13849 19147
rect 13935 19091 13991 19147
rect 14077 19091 14133 19147
rect 14219 19091 14275 19147
rect 14361 19091 14417 19147
rect 14503 19091 14559 19147
rect 14645 19091 14701 19147
rect 14787 19091 14843 19147
rect 161 18949 217 19005
rect 303 18949 359 19005
rect 445 18949 501 19005
rect 587 18949 643 19005
rect 729 18949 785 19005
rect 871 18949 927 19005
rect 1013 18949 1069 19005
rect 1155 18949 1211 19005
rect 1297 18949 1353 19005
rect 1439 18949 1495 19005
rect 1581 18949 1637 19005
rect 1723 18949 1779 19005
rect 1865 18949 1921 19005
rect 2007 18949 2063 19005
rect 2149 18949 2205 19005
rect 2291 18949 2347 19005
rect 2433 18949 2489 19005
rect 2575 18949 2631 19005
rect 2717 18949 2773 19005
rect 2859 18949 2915 19005
rect 3001 18949 3057 19005
rect 3143 18949 3199 19005
rect 3285 18949 3341 19005
rect 3427 18949 3483 19005
rect 3569 18949 3625 19005
rect 3711 18949 3767 19005
rect 3853 18949 3909 19005
rect 3995 18949 4051 19005
rect 4137 18949 4193 19005
rect 4279 18949 4335 19005
rect 4421 18949 4477 19005
rect 4563 18949 4619 19005
rect 4705 18949 4761 19005
rect 4847 18949 4903 19005
rect 4989 18949 5045 19005
rect 5131 18949 5187 19005
rect 5273 18949 5329 19005
rect 5415 18949 5471 19005
rect 5557 18949 5613 19005
rect 5699 18949 5755 19005
rect 5841 18949 5897 19005
rect 5983 18949 6039 19005
rect 6125 18949 6181 19005
rect 6267 18949 6323 19005
rect 6409 18949 6465 19005
rect 6551 18949 6607 19005
rect 6693 18949 6749 19005
rect 6835 18949 6891 19005
rect 6977 18949 7033 19005
rect 7119 18949 7175 19005
rect 7261 18949 7317 19005
rect 7403 18949 7459 19005
rect 7545 18949 7601 19005
rect 7687 18949 7743 19005
rect 7829 18949 7885 19005
rect 7971 18949 8027 19005
rect 8113 18949 8169 19005
rect 8255 18949 8311 19005
rect 8397 18949 8453 19005
rect 8539 18949 8595 19005
rect 8681 18949 8737 19005
rect 8823 18949 8879 19005
rect 8965 18949 9021 19005
rect 9107 18949 9163 19005
rect 9249 18949 9305 19005
rect 9391 18949 9447 19005
rect 9533 18949 9589 19005
rect 9675 18949 9731 19005
rect 9817 18949 9873 19005
rect 9959 18949 10015 19005
rect 10101 18949 10157 19005
rect 10243 18949 10299 19005
rect 10385 18949 10441 19005
rect 10527 18949 10583 19005
rect 10669 18949 10725 19005
rect 10811 18949 10867 19005
rect 10953 18949 11009 19005
rect 11095 18949 11151 19005
rect 11237 18949 11293 19005
rect 11379 18949 11435 19005
rect 11521 18949 11577 19005
rect 11663 18949 11719 19005
rect 11805 18949 11861 19005
rect 11947 18949 12003 19005
rect 12089 18949 12145 19005
rect 12231 18949 12287 19005
rect 12373 18949 12429 19005
rect 12515 18949 12571 19005
rect 12657 18949 12713 19005
rect 12799 18949 12855 19005
rect 12941 18949 12997 19005
rect 13083 18949 13139 19005
rect 13225 18949 13281 19005
rect 13367 18949 13423 19005
rect 13509 18949 13565 19005
rect 13651 18949 13707 19005
rect 13793 18949 13849 19005
rect 13935 18949 13991 19005
rect 14077 18949 14133 19005
rect 14219 18949 14275 19005
rect 14361 18949 14417 19005
rect 14503 18949 14559 19005
rect 14645 18949 14701 19005
rect 14787 18949 14843 19005
rect 161 18807 217 18863
rect 303 18807 359 18863
rect 445 18807 501 18863
rect 587 18807 643 18863
rect 729 18807 785 18863
rect 871 18807 927 18863
rect 1013 18807 1069 18863
rect 1155 18807 1211 18863
rect 1297 18807 1353 18863
rect 1439 18807 1495 18863
rect 1581 18807 1637 18863
rect 1723 18807 1779 18863
rect 1865 18807 1921 18863
rect 2007 18807 2063 18863
rect 2149 18807 2205 18863
rect 2291 18807 2347 18863
rect 2433 18807 2489 18863
rect 2575 18807 2631 18863
rect 2717 18807 2773 18863
rect 2859 18807 2915 18863
rect 3001 18807 3057 18863
rect 3143 18807 3199 18863
rect 3285 18807 3341 18863
rect 3427 18807 3483 18863
rect 3569 18807 3625 18863
rect 3711 18807 3767 18863
rect 3853 18807 3909 18863
rect 3995 18807 4051 18863
rect 4137 18807 4193 18863
rect 4279 18807 4335 18863
rect 4421 18807 4477 18863
rect 4563 18807 4619 18863
rect 4705 18807 4761 18863
rect 4847 18807 4903 18863
rect 4989 18807 5045 18863
rect 5131 18807 5187 18863
rect 5273 18807 5329 18863
rect 5415 18807 5471 18863
rect 5557 18807 5613 18863
rect 5699 18807 5755 18863
rect 5841 18807 5897 18863
rect 5983 18807 6039 18863
rect 6125 18807 6181 18863
rect 6267 18807 6323 18863
rect 6409 18807 6465 18863
rect 6551 18807 6607 18863
rect 6693 18807 6749 18863
rect 6835 18807 6891 18863
rect 6977 18807 7033 18863
rect 7119 18807 7175 18863
rect 7261 18807 7317 18863
rect 7403 18807 7459 18863
rect 7545 18807 7601 18863
rect 7687 18807 7743 18863
rect 7829 18807 7885 18863
rect 7971 18807 8027 18863
rect 8113 18807 8169 18863
rect 8255 18807 8311 18863
rect 8397 18807 8453 18863
rect 8539 18807 8595 18863
rect 8681 18807 8737 18863
rect 8823 18807 8879 18863
rect 8965 18807 9021 18863
rect 9107 18807 9163 18863
rect 9249 18807 9305 18863
rect 9391 18807 9447 18863
rect 9533 18807 9589 18863
rect 9675 18807 9731 18863
rect 9817 18807 9873 18863
rect 9959 18807 10015 18863
rect 10101 18807 10157 18863
rect 10243 18807 10299 18863
rect 10385 18807 10441 18863
rect 10527 18807 10583 18863
rect 10669 18807 10725 18863
rect 10811 18807 10867 18863
rect 10953 18807 11009 18863
rect 11095 18807 11151 18863
rect 11237 18807 11293 18863
rect 11379 18807 11435 18863
rect 11521 18807 11577 18863
rect 11663 18807 11719 18863
rect 11805 18807 11861 18863
rect 11947 18807 12003 18863
rect 12089 18807 12145 18863
rect 12231 18807 12287 18863
rect 12373 18807 12429 18863
rect 12515 18807 12571 18863
rect 12657 18807 12713 18863
rect 12799 18807 12855 18863
rect 12941 18807 12997 18863
rect 13083 18807 13139 18863
rect 13225 18807 13281 18863
rect 13367 18807 13423 18863
rect 13509 18807 13565 18863
rect 13651 18807 13707 18863
rect 13793 18807 13849 18863
rect 13935 18807 13991 18863
rect 14077 18807 14133 18863
rect 14219 18807 14275 18863
rect 14361 18807 14417 18863
rect 14503 18807 14559 18863
rect 14645 18807 14701 18863
rect 14787 18807 14843 18863
rect 161 18665 217 18721
rect 303 18665 359 18721
rect 445 18665 501 18721
rect 587 18665 643 18721
rect 729 18665 785 18721
rect 871 18665 927 18721
rect 1013 18665 1069 18721
rect 1155 18665 1211 18721
rect 1297 18665 1353 18721
rect 1439 18665 1495 18721
rect 1581 18665 1637 18721
rect 1723 18665 1779 18721
rect 1865 18665 1921 18721
rect 2007 18665 2063 18721
rect 2149 18665 2205 18721
rect 2291 18665 2347 18721
rect 2433 18665 2489 18721
rect 2575 18665 2631 18721
rect 2717 18665 2773 18721
rect 2859 18665 2915 18721
rect 3001 18665 3057 18721
rect 3143 18665 3199 18721
rect 3285 18665 3341 18721
rect 3427 18665 3483 18721
rect 3569 18665 3625 18721
rect 3711 18665 3767 18721
rect 3853 18665 3909 18721
rect 3995 18665 4051 18721
rect 4137 18665 4193 18721
rect 4279 18665 4335 18721
rect 4421 18665 4477 18721
rect 4563 18665 4619 18721
rect 4705 18665 4761 18721
rect 4847 18665 4903 18721
rect 4989 18665 5045 18721
rect 5131 18665 5187 18721
rect 5273 18665 5329 18721
rect 5415 18665 5471 18721
rect 5557 18665 5613 18721
rect 5699 18665 5755 18721
rect 5841 18665 5897 18721
rect 5983 18665 6039 18721
rect 6125 18665 6181 18721
rect 6267 18665 6323 18721
rect 6409 18665 6465 18721
rect 6551 18665 6607 18721
rect 6693 18665 6749 18721
rect 6835 18665 6891 18721
rect 6977 18665 7033 18721
rect 7119 18665 7175 18721
rect 7261 18665 7317 18721
rect 7403 18665 7459 18721
rect 7545 18665 7601 18721
rect 7687 18665 7743 18721
rect 7829 18665 7885 18721
rect 7971 18665 8027 18721
rect 8113 18665 8169 18721
rect 8255 18665 8311 18721
rect 8397 18665 8453 18721
rect 8539 18665 8595 18721
rect 8681 18665 8737 18721
rect 8823 18665 8879 18721
rect 8965 18665 9021 18721
rect 9107 18665 9163 18721
rect 9249 18665 9305 18721
rect 9391 18665 9447 18721
rect 9533 18665 9589 18721
rect 9675 18665 9731 18721
rect 9817 18665 9873 18721
rect 9959 18665 10015 18721
rect 10101 18665 10157 18721
rect 10243 18665 10299 18721
rect 10385 18665 10441 18721
rect 10527 18665 10583 18721
rect 10669 18665 10725 18721
rect 10811 18665 10867 18721
rect 10953 18665 11009 18721
rect 11095 18665 11151 18721
rect 11237 18665 11293 18721
rect 11379 18665 11435 18721
rect 11521 18665 11577 18721
rect 11663 18665 11719 18721
rect 11805 18665 11861 18721
rect 11947 18665 12003 18721
rect 12089 18665 12145 18721
rect 12231 18665 12287 18721
rect 12373 18665 12429 18721
rect 12515 18665 12571 18721
rect 12657 18665 12713 18721
rect 12799 18665 12855 18721
rect 12941 18665 12997 18721
rect 13083 18665 13139 18721
rect 13225 18665 13281 18721
rect 13367 18665 13423 18721
rect 13509 18665 13565 18721
rect 13651 18665 13707 18721
rect 13793 18665 13849 18721
rect 13935 18665 13991 18721
rect 14077 18665 14133 18721
rect 14219 18665 14275 18721
rect 14361 18665 14417 18721
rect 14503 18665 14559 18721
rect 14645 18665 14701 18721
rect 14787 18665 14843 18721
rect 161 18523 217 18579
rect 303 18523 359 18579
rect 445 18523 501 18579
rect 587 18523 643 18579
rect 729 18523 785 18579
rect 871 18523 927 18579
rect 1013 18523 1069 18579
rect 1155 18523 1211 18579
rect 1297 18523 1353 18579
rect 1439 18523 1495 18579
rect 1581 18523 1637 18579
rect 1723 18523 1779 18579
rect 1865 18523 1921 18579
rect 2007 18523 2063 18579
rect 2149 18523 2205 18579
rect 2291 18523 2347 18579
rect 2433 18523 2489 18579
rect 2575 18523 2631 18579
rect 2717 18523 2773 18579
rect 2859 18523 2915 18579
rect 3001 18523 3057 18579
rect 3143 18523 3199 18579
rect 3285 18523 3341 18579
rect 3427 18523 3483 18579
rect 3569 18523 3625 18579
rect 3711 18523 3767 18579
rect 3853 18523 3909 18579
rect 3995 18523 4051 18579
rect 4137 18523 4193 18579
rect 4279 18523 4335 18579
rect 4421 18523 4477 18579
rect 4563 18523 4619 18579
rect 4705 18523 4761 18579
rect 4847 18523 4903 18579
rect 4989 18523 5045 18579
rect 5131 18523 5187 18579
rect 5273 18523 5329 18579
rect 5415 18523 5471 18579
rect 5557 18523 5613 18579
rect 5699 18523 5755 18579
rect 5841 18523 5897 18579
rect 5983 18523 6039 18579
rect 6125 18523 6181 18579
rect 6267 18523 6323 18579
rect 6409 18523 6465 18579
rect 6551 18523 6607 18579
rect 6693 18523 6749 18579
rect 6835 18523 6891 18579
rect 6977 18523 7033 18579
rect 7119 18523 7175 18579
rect 7261 18523 7317 18579
rect 7403 18523 7459 18579
rect 7545 18523 7601 18579
rect 7687 18523 7743 18579
rect 7829 18523 7885 18579
rect 7971 18523 8027 18579
rect 8113 18523 8169 18579
rect 8255 18523 8311 18579
rect 8397 18523 8453 18579
rect 8539 18523 8595 18579
rect 8681 18523 8737 18579
rect 8823 18523 8879 18579
rect 8965 18523 9021 18579
rect 9107 18523 9163 18579
rect 9249 18523 9305 18579
rect 9391 18523 9447 18579
rect 9533 18523 9589 18579
rect 9675 18523 9731 18579
rect 9817 18523 9873 18579
rect 9959 18523 10015 18579
rect 10101 18523 10157 18579
rect 10243 18523 10299 18579
rect 10385 18523 10441 18579
rect 10527 18523 10583 18579
rect 10669 18523 10725 18579
rect 10811 18523 10867 18579
rect 10953 18523 11009 18579
rect 11095 18523 11151 18579
rect 11237 18523 11293 18579
rect 11379 18523 11435 18579
rect 11521 18523 11577 18579
rect 11663 18523 11719 18579
rect 11805 18523 11861 18579
rect 11947 18523 12003 18579
rect 12089 18523 12145 18579
rect 12231 18523 12287 18579
rect 12373 18523 12429 18579
rect 12515 18523 12571 18579
rect 12657 18523 12713 18579
rect 12799 18523 12855 18579
rect 12941 18523 12997 18579
rect 13083 18523 13139 18579
rect 13225 18523 13281 18579
rect 13367 18523 13423 18579
rect 13509 18523 13565 18579
rect 13651 18523 13707 18579
rect 13793 18523 13849 18579
rect 13935 18523 13991 18579
rect 14077 18523 14133 18579
rect 14219 18523 14275 18579
rect 14361 18523 14417 18579
rect 14503 18523 14559 18579
rect 14645 18523 14701 18579
rect 14787 18523 14843 18579
rect 161 18381 217 18437
rect 303 18381 359 18437
rect 445 18381 501 18437
rect 587 18381 643 18437
rect 729 18381 785 18437
rect 871 18381 927 18437
rect 1013 18381 1069 18437
rect 1155 18381 1211 18437
rect 1297 18381 1353 18437
rect 1439 18381 1495 18437
rect 1581 18381 1637 18437
rect 1723 18381 1779 18437
rect 1865 18381 1921 18437
rect 2007 18381 2063 18437
rect 2149 18381 2205 18437
rect 2291 18381 2347 18437
rect 2433 18381 2489 18437
rect 2575 18381 2631 18437
rect 2717 18381 2773 18437
rect 2859 18381 2915 18437
rect 3001 18381 3057 18437
rect 3143 18381 3199 18437
rect 3285 18381 3341 18437
rect 3427 18381 3483 18437
rect 3569 18381 3625 18437
rect 3711 18381 3767 18437
rect 3853 18381 3909 18437
rect 3995 18381 4051 18437
rect 4137 18381 4193 18437
rect 4279 18381 4335 18437
rect 4421 18381 4477 18437
rect 4563 18381 4619 18437
rect 4705 18381 4761 18437
rect 4847 18381 4903 18437
rect 4989 18381 5045 18437
rect 5131 18381 5187 18437
rect 5273 18381 5329 18437
rect 5415 18381 5471 18437
rect 5557 18381 5613 18437
rect 5699 18381 5755 18437
rect 5841 18381 5897 18437
rect 5983 18381 6039 18437
rect 6125 18381 6181 18437
rect 6267 18381 6323 18437
rect 6409 18381 6465 18437
rect 6551 18381 6607 18437
rect 6693 18381 6749 18437
rect 6835 18381 6891 18437
rect 6977 18381 7033 18437
rect 7119 18381 7175 18437
rect 7261 18381 7317 18437
rect 7403 18381 7459 18437
rect 7545 18381 7601 18437
rect 7687 18381 7743 18437
rect 7829 18381 7885 18437
rect 7971 18381 8027 18437
rect 8113 18381 8169 18437
rect 8255 18381 8311 18437
rect 8397 18381 8453 18437
rect 8539 18381 8595 18437
rect 8681 18381 8737 18437
rect 8823 18381 8879 18437
rect 8965 18381 9021 18437
rect 9107 18381 9163 18437
rect 9249 18381 9305 18437
rect 9391 18381 9447 18437
rect 9533 18381 9589 18437
rect 9675 18381 9731 18437
rect 9817 18381 9873 18437
rect 9959 18381 10015 18437
rect 10101 18381 10157 18437
rect 10243 18381 10299 18437
rect 10385 18381 10441 18437
rect 10527 18381 10583 18437
rect 10669 18381 10725 18437
rect 10811 18381 10867 18437
rect 10953 18381 11009 18437
rect 11095 18381 11151 18437
rect 11237 18381 11293 18437
rect 11379 18381 11435 18437
rect 11521 18381 11577 18437
rect 11663 18381 11719 18437
rect 11805 18381 11861 18437
rect 11947 18381 12003 18437
rect 12089 18381 12145 18437
rect 12231 18381 12287 18437
rect 12373 18381 12429 18437
rect 12515 18381 12571 18437
rect 12657 18381 12713 18437
rect 12799 18381 12855 18437
rect 12941 18381 12997 18437
rect 13083 18381 13139 18437
rect 13225 18381 13281 18437
rect 13367 18381 13423 18437
rect 13509 18381 13565 18437
rect 13651 18381 13707 18437
rect 13793 18381 13849 18437
rect 13935 18381 13991 18437
rect 14077 18381 14133 18437
rect 14219 18381 14275 18437
rect 14361 18381 14417 18437
rect 14503 18381 14559 18437
rect 14645 18381 14701 18437
rect 14787 18381 14843 18437
rect 161 18239 217 18295
rect 303 18239 359 18295
rect 445 18239 501 18295
rect 587 18239 643 18295
rect 729 18239 785 18295
rect 871 18239 927 18295
rect 1013 18239 1069 18295
rect 1155 18239 1211 18295
rect 1297 18239 1353 18295
rect 1439 18239 1495 18295
rect 1581 18239 1637 18295
rect 1723 18239 1779 18295
rect 1865 18239 1921 18295
rect 2007 18239 2063 18295
rect 2149 18239 2205 18295
rect 2291 18239 2347 18295
rect 2433 18239 2489 18295
rect 2575 18239 2631 18295
rect 2717 18239 2773 18295
rect 2859 18239 2915 18295
rect 3001 18239 3057 18295
rect 3143 18239 3199 18295
rect 3285 18239 3341 18295
rect 3427 18239 3483 18295
rect 3569 18239 3625 18295
rect 3711 18239 3767 18295
rect 3853 18239 3909 18295
rect 3995 18239 4051 18295
rect 4137 18239 4193 18295
rect 4279 18239 4335 18295
rect 4421 18239 4477 18295
rect 4563 18239 4619 18295
rect 4705 18239 4761 18295
rect 4847 18239 4903 18295
rect 4989 18239 5045 18295
rect 5131 18239 5187 18295
rect 5273 18239 5329 18295
rect 5415 18239 5471 18295
rect 5557 18239 5613 18295
rect 5699 18239 5755 18295
rect 5841 18239 5897 18295
rect 5983 18239 6039 18295
rect 6125 18239 6181 18295
rect 6267 18239 6323 18295
rect 6409 18239 6465 18295
rect 6551 18239 6607 18295
rect 6693 18239 6749 18295
rect 6835 18239 6891 18295
rect 6977 18239 7033 18295
rect 7119 18239 7175 18295
rect 7261 18239 7317 18295
rect 7403 18239 7459 18295
rect 7545 18239 7601 18295
rect 7687 18239 7743 18295
rect 7829 18239 7885 18295
rect 7971 18239 8027 18295
rect 8113 18239 8169 18295
rect 8255 18239 8311 18295
rect 8397 18239 8453 18295
rect 8539 18239 8595 18295
rect 8681 18239 8737 18295
rect 8823 18239 8879 18295
rect 8965 18239 9021 18295
rect 9107 18239 9163 18295
rect 9249 18239 9305 18295
rect 9391 18239 9447 18295
rect 9533 18239 9589 18295
rect 9675 18239 9731 18295
rect 9817 18239 9873 18295
rect 9959 18239 10015 18295
rect 10101 18239 10157 18295
rect 10243 18239 10299 18295
rect 10385 18239 10441 18295
rect 10527 18239 10583 18295
rect 10669 18239 10725 18295
rect 10811 18239 10867 18295
rect 10953 18239 11009 18295
rect 11095 18239 11151 18295
rect 11237 18239 11293 18295
rect 11379 18239 11435 18295
rect 11521 18239 11577 18295
rect 11663 18239 11719 18295
rect 11805 18239 11861 18295
rect 11947 18239 12003 18295
rect 12089 18239 12145 18295
rect 12231 18239 12287 18295
rect 12373 18239 12429 18295
rect 12515 18239 12571 18295
rect 12657 18239 12713 18295
rect 12799 18239 12855 18295
rect 12941 18239 12997 18295
rect 13083 18239 13139 18295
rect 13225 18239 13281 18295
rect 13367 18239 13423 18295
rect 13509 18239 13565 18295
rect 13651 18239 13707 18295
rect 13793 18239 13849 18295
rect 13935 18239 13991 18295
rect 14077 18239 14133 18295
rect 14219 18239 14275 18295
rect 14361 18239 14417 18295
rect 14503 18239 14559 18295
rect 14645 18239 14701 18295
rect 14787 18239 14843 18295
rect 161 18097 217 18153
rect 303 18097 359 18153
rect 445 18097 501 18153
rect 587 18097 643 18153
rect 729 18097 785 18153
rect 871 18097 927 18153
rect 1013 18097 1069 18153
rect 1155 18097 1211 18153
rect 1297 18097 1353 18153
rect 1439 18097 1495 18153
rect 1581 18097 1637 18153
rect 1723 18097 1779 18153
rect 1865 18097 1921 18153
rect 2007 18097 2063 18153
rect 2149 18097 2205 18153
rect 2291 18097 2347 18153
rect 2433 18097 2489 18153
rect 2575 18097 2631 18153
rect 2717 18097 2773 18153
rect 2859 18097 2915 18153
rect 3001 18097 3057 18153
rect 3143 18097 3199 18153
rect 3285 18097 3341 18153
rect 3427 18097 3483 18153
rect 3569 18097 3625 18153
rect 3711 18097 3767 18153
rect 3853 18097 3909 18153
rect 3995 18097 4051 18153
rect 4137 18097 4193 18153
rect 4279 18097 4335 18153
rect 4421 18097 4477 18153
rect 4563 18097 4619 18153
rect 4705 18097 4761 18153
rect 4847 18097 4903 18153
rect 4989 18097 5045 18153
rect 5131 18097 5187 18153
rect 5273 18097 5329 18153
rect 5415 18097 5471 18153
rect 5557 18097 5613 18153
rect 5699 18097 5755 18153
rect 5841 18097 5897 18153
rect 5983 18097 6039 18153
rect 6125 18097 6181 18153
rect 6267 18097 6323 18153
rect 6409 18097 6465 18153
rect 6551 18097 6607 18153
rect 6693 18097 6749 18153
rect 6835 18097 6891 18153
rect 6977 18097 7033 18153
rect 7119 18097 7175 18153
rect 7261 18097 7317 18153
rect 7403 18097 7459 18153
rect 7545 18097 7601 18153
rect 7687 18097 7743 18153
rect 7829 18097 7885 18153
rect 7971 18097 8027 18153
rect 8113 18097 8169 18153
rect 8255 18097 8311 18153
rect 8397 18097 8453 18153
rect 8539 18097 8595 18153
rect 8681 18097 8737 18153
rect 8823 18097 8879 18153
rect 8965 18097 9021 18153
rect 9107 18097 9163 18153
rect 9249 18097 9305 18153
rect 9391 18097 9447 18153
rect 9533 18097 9589 18153
rect 9675 18097 9731 18153
rect 9817 18097 9873 18153
rect 9959 18097 10015 18153
rect 10101 18097 10157 18153
rect 10243 18097 10299 18153
rect 10385 18097 10441 18153
rect 10527 18097 10583 18153
rect 10669 18097 10725 18153
rect 10811 18097 10867 18153
rect 10953 18097 11009 18153
rect 11095 18097 11151 18153
rect 11237 18097 11293 18153
rect 11379 18097 11435 18153
rect 11521 18097 11577 18153
rect 11663 18097 11719 18153
rect 11805 18097 11861 18153
rect 11947 18097 12003 18153
rect 12089 18097 12145 18153
rect 12231 18097 12287 18153
rect 12373 18097 12429 18153
rect 12515 18097 12571 18153
rect 12657 18097 12713 18153
rect 12799 18097 12855 18153
rect 12941 18097 12997 18153
rect 13083 18097 13139 18153
rect 13225 18097 13281 18153
rect 13367 18097 13423 18153
rect 13509 18097 13565 18153
rect 13651 18097 13707 18153
rect 13793 18097 13849 18153
rect 13935 18097 13991 18153
rect 14077 18097 14133 18153
rect 14219 18097 14275 18153
rect 14361 18097 14417 18153
rect 14503 18097 14559 18153
rect 14645 18097 14701 18153
rect 14787 18097 14843 18153
rect 161 17955 217 18011
rect 303 17955 359 18011
rect 445 17955 501 18011
rect 587 17955 643 18011
rect 729 17955 785 18011
rect 871 17955 927 18011
rect 1013 17955 1069 18011
rect 1155 17955 1211 18011
rect 1297 17955 1353 18011
rect 1439 17955 1495 18011
rect 1581 17955 1637 18011
rect 1723 17955 1779 18011
rect 1865 17955 1921 18011
rect 2007 17955 2063 18011
rect 2149 17955 2205 18011
rect 2291 17955 2347 18011
rect 2433 17955 2489 18011
rect 2575 17955 2631 18011
rect 2717 17955 2773 18011
rect 2859 17955 2915 18011
rect 3001 17955 3057 18011
rect 3143 17955 3199 18011
rect 3285 17955 3341 18011
rect 3427 17955 3483 18011
rect 3569 17955 3625 18011
rect 3711 17955 3767 18011
rect 3853 17955 3909 18011
rect 3995 17955 4051 18011
rect 4137 17955 4193 18011
rect 4279 17955 4335 18011
rect 4421 17955 4477 18011
rect 4563 17955 4619 18011
rect 4705 17955 4761 18011
rect 4847 17955 4903 18011
rect 4989 17955 5045 18011
rect 5131 17955 5187 18011
rect 5273 17955 5329 18011
rect 5415 17955 5471 18011
rect 5557 17955 5613 18011
rect 5699 17955 5755 18011
rect 5841 17955 5897 18011
rect 5983 17955 6039 18011
rect 6125 17955 6181 18011
rect 6267 17955 6323 18011
rect 6409 17955 6465 18011
rect 6551 17955 6607 18011
rect 6693 17955 6749 18011
rect 6835 17955 6891 18011
rect 6977 17955 7033 18011
rect 7119 17955 7175 18011
rect 7261 17955 7317 18011
rect 7403 17955 7459 18011
rect 7545 17955 7601 18011
rect 7687 17955 7743 18011
rect 7829 17955 7885 18011
rect 7971 17955 8027 18011
rect 8113 17955 8169 18011
rect 8255 17955 8311 18011
rect 8397 17955 8453 18011
rect 8539 17955 8595 18011
rect 8681 17955 8737 18011
rect 8823 17955 8879 18011
rect 8965 17955 9021 18011
rect 9107 17955 9163 18011
rect 9249 17955 9305 18011
rect 9391 17955 9447 18011
rect 9533 17955 9589 18011
rect 9675 17955 9731 18011
rect 9817 17955 9873 18011
rect 9959 17955 10015 18011
rect 10101 17955 10157 18011
rect 10243 17955 10299 18011
rect 10385 17955 10441 18011
rect 10527 17955 10583 18011
rect 10669 17955 10725 18011
rect 10811 17955 10867 18011
rect 10953 17955 11009 18011
rect 11095 17955 11151 18011
rect 11237 17955 11293 18011
rect 11379 17955 11435 18011
rect 11521 17955 11577 18011
rect 11663 17955 11719 18011
rect 11805 17955 11861 18011
rect 11947 17955 12003 18011
rect 12089 17955 12145 18011
rect 12231 17955 12287 18011
rect 12373 17955 12429 18011
rect 12515 17955 12571 18011
rect 12657 17955 12713 18011
rect 12799 17955 12855 18011
rect 12941 17955 12997 18011
rect 13083 17955 13139 18011
rect 13225 17955 13281 18011
rect 13367 17955 13423 18011
rect 13509 17955 13565 18011
rect 13651 17955 13707 18011
rect 13793 17955 13849 18011
rect 13935 17955 13991 18011
rect 14077 17955 14133 18011
rect 14219 17955 14275 18011
rect 14361 17955 14417 18011
rect 14503 17955 14559 18011
rect 14645 17955 14701 18011
rect 14787 17955 14843 18011
rect 161 17813 217 17869
rect 303 17813 359 17869
rect 445 17813 501 17869
rect 587 17813 643 17869
rect 729 17813 785 17869
rect 871 17813 927 17869
rect 1013 17813 1069 17869
rect 1155 17813 1211 17869
rect 1297 17813 1353 17869
rect 1439 17813 1495 17869
rect 1581 17813 1637 17869
rect 1723 17813 1779 17869
rect 1865 17813 1921 17869
rect 2007 17813 2063 17869
rect 2149 17813 2205 17869
rect 2291 17813 2347 17869
rect 2433 17813 2489 17869
rect 2575 17813 2631 17869
rect 2717 17813 2773 17869
rect 2859 17813 2915 17869
rect 3001 17813 3057 17869
rect 3143 17813 3199 17869
rect 3285 17813 3341 17869
rect 3427 17813 3483 17869
rect 3569 17813 3625 17869
rect 3711 17813 3767 17869
rect 3853 17813 3909 17869
rect 3995 17813 4051 17869
rect 4137 17813 4193 17869
rect 4279 17813 4335 17869
rect 4421 17813 4477 17869
rect 4563 17813 4619 17869
rect 4705 17813 4761 17869
rect 4847 17813 4903 17869
rect 4989 17813 5045 17869
rect 5131 17813 5187 17869
rect 5273 17813 5329 17869
rect 5415 17813 5471 17869
rect 5557 17813 5613 17869
rect 5699 17813 5755 17869
rect 5841 17813 5897 17869
rect 5983 17813 6039 17869
rect 6125 17813 6181 17869
rect 6267 17813 6323 17869
rect 6409 17813 6465 17869
rect 6551 17813 6607 17869
rect 6693 17813 6749 17869
rect 6835 17813 6891 17869
rect 6977 17813 7033 17869
rect 7119 17813 7175 17869
rect 7261 17813 7317 17869
rect 7403 17813 7459 17869
rect 7545 17813 7601 17869
rect 7687 17813 7743 17869
rect 7829 17813 7885 17869
rect 7971 17813 8027 17869
rect 8113 17813 8169 17869
rect 8255 17813 8311 17869
rect 8397 17813 8453 17869
rect 8539 17813 8595 17869
rect 8681 17813 8737 17869
rect 8823 17813 8879 17869
rect 8965 17813 9021 17869
rect 9107 17813 9163 17869
rect 9249 17813 9305 17869
rect 9391 17813 9447 17869
rect 9533 17813 9589 17869
rect 9675 17813 9731 17869
rect 9817 17813 9873 17869
rect 9959 17813 10015 17869
rect 10101 17813 10157 17869
rect 10243 17813 10299 17869
rect 10385 17813 10441 17869
rect 10527 17813 10583 17869
rect 10669 17813 10725 17869
rect 10811 17813 10867 17869
rect 10953 17813 11009 17869
rect 11095 17813 11151 17869
rect 11237 17813 11293 17869
rect 11379 17813 11435 17869
rect 11521 17813 11577 17869
rect 11663 17813 11719 17869
rect 11805 17813 11861 17869
rect 11947 17813 12003 17869
rect 12089 17813 12145 17869
rect 12231 17813 12287 17869
rect 12373 17813 12429 17869
rect 12515 17813 12571 17869
rect 12657 17813 12713 17869
rect 12799 17813 12855 17869
rect 12941 17813 12997 17869
rect 13083 17813 13139 17869
rect 13225 17813 13281 17869
rect 13367 17813 13423 17869
rect 13509 17813 13565 17869
rect 13651 17813 13707 17869
rect 13793 17813 13849 17869
rect 13935 17813 13991 17869
rect 14077 17813 14133 17869
rect 14219 17813 14275 17869
rect 14361 17813 14417 17869
rect 14503 17813 14559 17869
rect 14645 17813 14701 17869
rect 14787 17813 14843 17869
rect 161 17671 217 17727
rect 303 17671 359 17727
rect 445 17671 501 17727
rect 587 17671 643 17727
rect 729 17671 785 17727
rect 871 17671 927 17727
rect 1013 17671 1069 17727
rect 1155 17671 1211 17727
rect 1297 17671 1353 17727
rect 1439 17671 1495 17727
rect 1581 17671 1637 17727
rect 1723 17671 1779 17727
rect 1865 17671 1921 17727
rect 2007 17671 2063 17727
rect 2149 17671 2205 17727
rect 2291 17671 2347 17727
rect 2433 17671 2489 17727
rect 2575 17671 2631 17727
rect 2717 17671 2773 17727
rect 2859 17671 2915 17727
rect 3001 17671 3057 17727
rect 3143 17671 3199 17727
rect 3285 17671 3341 17727
rect 3427 17671 3483 17727
rect 3569 17671 3625 17727
rect 3711 17671 3767 17727
rect 3853 17671 3909 17727
rect 3995 17671 4051 17727
rect 4137 17671 4193 17727
rect 4279 17671 4335 17727
rect 4421 17671 4477 17727
rect 4563 17671 4619 17727
rect 4705 17671 4761 17727
rect 4847 17671 4903 17727
rect 4989 17671 5045 17727
rect 5131 17671 5187 17727
rect 5273 17671 5329 17727
rect 5415 17671 5471 17727
rect 5557 17671 5613 17727
rect 5699 17671 5755 17727
rect 5841 17671 5897 17727
rect 5983 17671 6039 17727
rect 6125 17671 6181 17727
rect 6267 17671 6323 17727
rect 6409 17671 6465 17727
rect 6551 17671 6607 17727
rect 6693 17671 6749 17727
rect 6835 17671 6891 17727
rect 6977 17671 7033 17727
rect 7119 17671 7175 17727
rect 7261 17671 7317 17727
rect 7403 17671 7459 17727
rect 7545 17671 7601 17727
rect 7687 17671 7743 17727
rect 7829 17671 7885 17727
rect 7971 17671 8027 17727
rect 8113 17671 8169 17727
rect 8255 17671 8311 17727
rect 8397 17671 8453 17727
rect 8539 17671 8595 17727
rect 8681 17671 8737 17727
rect 8823 17671 8879 17727
rect 8965 17671 9021 17727
rect 9107 17671 9163 17727
rect 9249 17671 9305 17727
rect 9391 17671 9447 17727
rect 9533 17671 9589 17727
rect 9675 17671 9731 17727
rect 9817 17671 9873 17727
rect 9959 17671 10015 17727
rect 10101 17671 10157 17727
rect 10243 17671 10299 17727
rect 10385 17671 10441 17727
rect 10527 17671 10583 17727
rect 10669 17671 10725 17727
rect 10811 17671 10867 17727
rect 10953 17671 11009 17727
rect 11095 17671 11151 17727
rect 11237 17671 11293 17727
rect 11379 17671 11435 17727
rect 11521 17671 11577 17727
rect 11663 17671 11719 17727
rect 11805 17671 11861 17727
rect 11947 17671 12003 17727
rect 12089 17671 12145 17727
rect 12231 17671 12287 17727
rect 12373 17671 12429 17727
rect 12515 17671 12571 17727
rect 12657 17671 12713 17727
rect 12799 17671 12855 17727
rect 12941 17671 12997 17727
rect 13083 17671 13139 17727
rect 13225 17671 13281 17727
rect 13367 17671 13423 17727
rect 13509 17671 13565 17727
rect 13651 17671 13707 17727
rect 13793 17671 13849 17727
rect 13935 17671 13991 17727
rect 14077 17671 14133 17727
rect 14219 17671 14275 17727
rect 14361 17671 14417 17727
rect 14503 17671 14559 17727
rect 14645 17671 14701 17727
rect 14787 17671 14843 17727
rect 161 17529 217 17585
rect 303 17529 359 17585
rect 445 17529 501 17585
rect 587 17529 643 17585
rect 729 17529 785 17585
rect 871 17529 927 17585
rect 1013 17529 1069 17585
rect 1155 17529 1211 17585
rect 1297 17529 1353 17585
rect 1439 17529 1495 17585
rect 1581 17529 1637 17585
rect 1723 17529 1779 17585
rect 1865 17529 1921 17585
rect 2007 17529 2063 17585
rect 2149 17529 2205 17585
rect 2291 17529 2347 17585
rect 2433 17529 2489 17585
rect 2575 17529 2631 17585
rect 2717 17529 2773 17585
rect 2859 17529 2915 17585
rect 3001 17529 3057 17585
rect 3143 17529 3199 17585
rect 3285 17529 3341 17585
rect 3427 17529 3483 17585
rect 3569 17529 3625 17585
rect 3711 17529 3767 17585
rect 3853 17529 3909 17585
rect 3995 17529 4051 17585
rect 4137 17529 4193 17585
rect 4279 17529 4335 17585
rect 4421 17529 4477 17585
rect 4563 17529 4619 17585
rect 4705 17529 4761 17585
rect 4847 17529 4903 17585
rect 4989 17529 5045 17585
rect 5131 17529 5187 17585
rect 5273 17529 5329 17585
rect 5415 17529 5471 17585
rect 5557 17529 5613 17585
rect 5699 17529 5755 17585
rect 5841 17529 5897 17585
rect 5983 17529 6039 17585
rect 6125 17529 6181 17585
rect 6267 17529 6323 17585
rect 6409 17529 6465 17585
rect 6551 17529 6607 17585
rect 6693 17529 6749 17585
rect 6835 17529 6891 17585
rect 6977 17529 7033 17585
rect 7119 17529 7175 17585
rect 7261 17529 7317 17585
rect 7403 17529 7459 17585
rect 7545 17529 7601 17585
rect 7687 17529 7743 17585
rect 7829 17529 7885 17585
rect 7971 17529 8027 17585
rect 8113 17529 8169 17585
rect 8255 17529 8311 17585
rect 8397 17529 8453 17585
rect 8539 17529 8595 17585
rect 8681 17529 8737 17585
rect 8823 17529 8879 17585
rect 8965 17529 9021 17585
rect 9107 17529 9163 17585
rect 9249 17529 9305 17585
rect 9391 17529 9447 17585
rect 9533 17529 9589 17585
rect 9675 17529 9731 17585
rect 9817 17529 9873 17585
rect 9959 17529 10015 17585
rect 10101 17529 10157 17585
rect 10243 17529 10299 17585
rect 10385 17529 10441 17585
rect 10527 17529 10583 17585
rect 10669 17529 10725 17585
rect 10811 17529 10867 17585
rect 10953 17529 11009 17585
rect 11095 17529 11151 17585
rect 11237 17529 11293 17585
rect 11379 17529 11435 17585
rect 11521 17529 11577 17585
rect 11663 17529 11719 17585
rect 11805 17529 11861 17585
rect 11947 17529 12003 17585
rect 12089 17529 12145 17585
rect 12231 17529 12287 17585
rect 12373 17529 12429 17585
rect 12515 17529 12571 17585
rect 12657 17529 12713 17585
rect 12799 17529 12855 17585
rect 12941 17529 12997 17585
rect 13083 17529 13139 17585
rect 13225 17529 13281 17585
rect 13367 17529 13423 17585
rect 13509 17529 13565 17585
rect 13651 17529 13707 17585
rect 13793 17529 13849 17585
rect 13935 17529 13991 17585
rect 14077 17529 14133 17585
rect 14219 17529 14275 17585
rect 14361 17529 14417 17585
rect 14503 17529 14559 17585
rect 14645 17529 14701 17585
rect 14787 17529 14843 17585
rect 161 17387 217 17443
rect 303 17387 359 17443
rect 445 17387 501 17443
rect 587 17387 643 17443
rect 729 17387 785 17443
rect 871 17387 927 17443
rect 1013 17387 1069 17443
rect 1155 17387 1211 17443
rect 1297 17387 1353 17443
rect 1439 17387 1495 17443
rect 1581 17387 1637 17443
rect 1723 17387 1779 17443
rect 1865 17387 1921 17443
rect 2007 17387 2063 17443
rect 2149 17387 2205 17443
rect 2291 17387 2347 17443
rect 2433 17387 2489 17443
rect 2575 17387 2631 17443
rect 2717 17387 2773 17443
rect 2859 17387 2915 17443
rect 3001 17387 3057 17443
rect 3143 17387 3199 17443
rect 3285 17387 3341 17443
rect 3427 17387 3483 17443
rect 3569 17387 3625 17443
rect 3711 17387 3767 17443
rect 3853 17387 3909 17443
rect 3995 17387 4051 17443
rect 4137 17387 4193 17443
rect 4279 17387 4335 17443
rect 4421 17387 4477 17443
rect 4563 17387 4619 17443
rect 4705 17387 4761 17443
rect 4847 17387 4903 17443
rect 4989 17387 5045 17443
rect 5131 17387 5187 17443
rect 5273 17387 5329 17443
rect 5415 17387 5471 17443
rect 5557 17387 5613 17443
rect 5699 17387 5755 17443
rect 5841 17387 5897 17443
rect 5983 17387 6039 17443
rect 6125 17387 6181 17443
rect 6267 17387 6323 17443
rect 6409 17387 6465 17443
rect 6551 17387 6607 17443
rect 6693 17387 6749 17443
rect 6835 17387 6891 17443
rect 6977 17387 7033 17443
rect 7119 17387 7175 17443
rect 7261 17387 7317 17443
rect 7403 17387 7459 17443
rect 7545 17387 7601 17443
rect 7687 17387 7743 17443
rect 7829 17387 7885 17443
rect 7971 17387 8027 17443
rect 8113 17387 8169 17443
rect 8255 17387 8311 17443
rect 8397 17387 8453 17443
rect 8539 17387 8595 17443
rect 8681 17387 8737 17443
rect 8823 17387 8879 17443
rect 8965 17387 9021 17443
rect 9107 17387 9163 17443
rect 9249 17387 9305 17443
rect 9391 17387 9447 17443
rect 9533 17387 9589 17443
rect 9675 17387 9731 17443
rect 9817 17387 9873 17443
rect 9959 17387 10015 17443
rect 10101 17387 10157 17443
rect 10243 17387 10299 17443
rect 10385 17387 10441 17443
rect 10527 17387 10583 17443
rect 10669 17387 10725 17443
rect 10811 17387 10867 17443
rect 10953 17387 11009 17443
rect 11095 17387 11151 17443
rect 11237 17387 11293 17443
rect 11379 17387 11435 17443
rect 11521 17387 11577 17443
rect 11663 17387 11719 17443
rect 11805 17387 11861 17443
rect 11947 17387 12003 17443
rect 12089 17387 12145 17443
rect 12231 17387 12287 17443
rect 12373 17387 12429 17443
rect 12515 17387 12571 17443
rect 12657 17387 12713 17443
rect 12799 17387 12855 17443
rect 12941 17387 12997 17443
rect 13083 17387 13139 17443
rect 13225 17387 13281 17443
rect 13367 17387 13423 17443
rect 13509 17387 13565 17443
rect 13651 17387 13707 17443
rect 13793 17387 13849 17443
rect 13935 17387 13991 17443
rect 14077 17387 14133 17443
rect 14219 17387 14275 17443
rect 14361 17387 14417 17443
rect 14503 17387 14559 17443
rect 14645 17387 14701 17443
rect 14787 17387 14843 17443
rect 161 17245 217 17301
rect 303 17245 359 17301
rect 445 17245 501 17301
rect 587 17245 643 17301
rect 729 17245 785 17301
rect 871 17245 927 17301
rect 1013 17245 1069 17301
rect 1155 17245 1211 17301
rect 1297 17245 1353 17301
rect 1439 17245 1495 17301
rect 1581 17245 1637 17301
rect 1723 17245 1779 17301
rect 1865 17245 1921 17301
rect 2007 17245 2063 17301
rect 2149 17245 2205 17301
rect 2291 17245 2347 17301
rect 2433 17245 2489 17301
rect 2575 17245 2631 17301
rect 2717 17245 2773 17301
rect 2859 17245 2915 17301
rect 3001 17245 3057 17301
rect 3143 17245 3199 17301
rect 3285 17245 3341 17301
rect 3427 17245 3483 17301
rect 3569 17245 3625 17301
rect 3711 17245 3767 17301
rect 3853 17245 3909 17301
rect 3995 17245 4051 17301
rect 4137 17245 4193 17301
rect 4279 17245 4335 17301
rect 4421 17245 4477 17301
rect 4563 17245 4619 17301
rect 4705 17245 4761 17301
rect 4847 17245 4903 17301
rect 4989 17245 5045 17301
rect 5131 17245 5187 17301
rect 5273 17245 5329 17301
rect 5415 17245 5471 17301
rect 5557 17245 5613 17301
rect 5699 17245 5755 17301
rect 5841 17245 5897 17301
rect 5983 17245 6039 17301
rect 6125 17245 6181 17301
rect 6267 17245 6323 17301
rect 6409 17245 6465 17301
rect 6551 17245 6607 17301
rect 6693 17245 6749 17301
rect 6835 17245 6891 17301
rect 6977 17245 7033 17301
rect 7119 17245 7175 17301
rect 7261 17245 7317 17301
rect 7403 17245 7459 17301
rect 7545 17245 7601 17301
rect 7687 17245 7743 17301
rect 7829 17245 7885 17301
rect 7971 17245 8027 17301
rect 8113 17245 8169 17301
rect 8255 17245 8311 17301
rect 8397 17245 8453 17301
rect 8539 17245 8595 17301
rect 8681 17245 8737 17301
rect 8823 17245 8879 17301
rect 8965 17245 9021 17301
rect 9107 17245 9163 17301
rect 9249 17245 9305 17301
rect 9391 17245 9447 17301
rect 9533 17245 9589 17301
rect 9675 17245 9731 17301
rect 9817 17245 9873 17301
rect 9959 17245 10015 17301
rect 10101 17245 10157 17301
rect 10243 17245 10299 17301
rect 10385 17245 10441 17301
rect 10527 17245 10583 17301
rect 10669 17245 10725 17301
rect 10811 17245 10867 17301
rect 10953 17245 11009 17301
rect 11095 17245 11151 17301
rect 11237 17245 11293 17301
rect 11379 17245 11435 17301
rect 11521 17245 11577 17301
rect 11663 17245 11719 17301
rect 11805 17245 11861 17301
rect 11947 17245 12003 17301
rect 12089 17245 12145 17301
rect 12231 17245 12287 17301
rect 12373 17245 12429 17301
rect 12515 17245 12571 17301
rect 12657 17245 12713 17301
rect 12799 17245 12855 17301
rect 12941 17245 12997 17301
rect 13083 17245 13139 17301
rect 13225 17245 13281 17301
rect 13367 17245 13423 17301
rect 13509 17245 13565 17301
rect 13651 17245 13707 17301
rect 13793 17245 13849 17301
rect 13935 17245 13991 17301
rect 14077 17245 14133 17301
rect 14219 17245 14275 17301
rect 14361 17245 14417 17301
rect 14503 17245 14559 17301
rect 14645 17245 14701 17301
rect 14787 17245 14843 17301
rect 161 16885 217 16941
rect 303 16885 359 16941
rect 445 16885 501 16941
rect 587 16885 643 16941
rect 729 16885 785 16941
rect 871 16885 927 16941
rect 1013 16885 1069 16941
rect 1155 16885 1211 16941
rect 1297 16885 1353 16941
rect 1439 16885 1495 16941
rect 1581 16885 1637 16941
rect 1723 16885 1779 16941
rect 1865 16885 1921 16941
rect 2007 16885 2063 16941
rect 2149 16885 2205 16941
rect 2291 16885 2347 16941
rect 2433 16885 2489 16941
rect 2575 16885 2631 16941
rect 2717 16885 2773 16941
rect 2859 16885 2915 16941
rect 3001 16885 3057 16941
rect 3143 16885 3199 16941
rect 3285 16885 3341 16941
rect 3427 16885 3483 16941
rect 3569 16885 3625 16941
rect 3711 16885 3767 16941
rect 3853 16885 3909 16941
rect 3995 16885 4051 16941
rect 4137 16885 4193 16941
rect 4279 16885 4335 16941
rect 4421 16885 4477 16941
rect 4563 16885 4619 16941
rect 4705 16885 4761 16941
rect 4847 16885 4903 16941
rect 4989 16885 5045 16941
rect 5131 16885 5187 16941
rect 5273 16885 5329 16941
rect 5415 16885 5471 16941
rect 5557 16885 5613 16941
rect 5699 16885 5755 16941
rect 5841 16885 5897 16941
rect 5983 16885 6039 16941
rect 6125 16885 6181 16941
rect 6267 16885 6323 16941
rect 6409 16885 6465 16941
rect 6551 16885 6607 16941
rect 6693 16885 6749 16941
rect 6835 16885 6891 16941
rect 6977 16885 7033 16941
rect 7119 16885 7175 16941
rect 7261 16885 7317 16941
rect 7403 16885 7459 16941
rect 7545 16885 7601 16941
rect 7687 16885 7743 16941
rect 7829 16885 7885 16941
rect 7971 16885 8027 16941
rect 8113 16885 8169 16941
rect 8255 16885 8311 16941
rect 8397 16885 8453 16941
rect 8539 16885 8595 16941
rect 8681 16885 8737 16941
rect 8823 16885 8879 16941
rect 8965 16885 9021 16941
rect 9107 16885 9163 16941
rect 9249 16885 9305 16941
rect 9391 16885 9447 16941
rect 9533 16885 9589 16941
rect 9675 16885 9731 16941
rect 9817 16885 9873 16941
rect 9959 16885 10015 16941
rect 10101 16885 10157 16941
rect 10243 16885 10299 16941
rect 10385 16885 10441 16941
rect 10527 16885 10583 16941
rect 10669 16885 10725 16941
rect 10811 16885 10867 16941
rect 10953 16885 11009 16941
rect 11095 16885 11151 16941
rect 11237 16885 11293 16941
rect 11379 16885 11435 16941
rect 11521 16885 11577 16941
rect 11663 16885 11719 16941
rect 11805 16885 11861 16941
rect 11947 16885 12003 16941
rect 12089 16885 12145 16941
rect 12231 16885 12287 16941
rect 12373 16885 12429 16941
rect 12515 16885 12571 16941
rect 12657 16885 12713 16941
rect 12799 16885 12855 16941
rect 12941 16885 12997 16941
rect 13083 16885 13139 16941
rect 13225 16885 13281 16941
rect 13367 16885 13423 16941
rect 13509 16885 13565 16941
rect 13651 16885 13707 16941
rect 13793 16885 13849 16941
rect 13935 16885 13991 16941
rect 14077 16885 14133 16941
rect 14219 16885 14275 16941
rect 14361 16885 14417 16941
rect 14503 16885 14559 16941
rect 14645 16885 14701 16941
rect 14787 16885 14843 16941
rect 161 16743 217 16799
rect 303 16743 359 16799
rect 445 16743 501 16799
rect 587 16743 643 16799
rect 729 16743 785 16799
rect 871 16743 927 16799
rect 1013 16743 1069 16799
rect 1155 16743 1211 16799
rect 1297 16743 1353 16799
rect 1439 16743 1495 16799
rect 1581 16743 1637 16799
rect 1723 16743 1779 16799
rect 1865 16743 1921 16799
rect 2007 16743 2063 16799
rect 2149 16743 2205 16799
rect 2291 16743 2347 16799
rect 2433 16743 2489 16799
rect 2575 16743 2631 16799
rect 2717 16743 2773 16799
rect 2859 16743 2915 16799
rect 3001 16743 3057 16799
rect 3143 16743 3199 16799
rect 3285 16743 3341 16799
rect 3427 16743 3483 16799
rect 3569 16743 3625 16799
rect 3711 16743 3767 16799
rect 3853 16743 3909 16799
rect 3995 16743 4051 16799
rect 4137 16743 4193 16799
rect 4279 16743 4335 16799
rect 4421 16743 4477 16799
rect 4563 16743 4619 16799
rect 4705 16743 4761 16799
rect 4847 16743 4903 16799
rect 4989 16743 5045 16799
rect 5131 16743 5187 16799
rect 5273 16743 5329 16799
rect 5415 16743 5471 16799
rect 5557 16743 5613 16799
rect 5699 16743 5755 16799
rect 5841 16743 5897 16799
rect 5983 16743 6039 16799
rect 6125 16743 6181 16799
rect 6267 16743 6323 16799
rect 6409 16743 6465 16799
rect 6551 16743 6607 16799
rect 6693 16743 6749 16799
rect 6835 16743 6891 16799
rect 6977 16743 7033 16799
rect 7119 16743 7175 16799
rect 7261 16743 7317 16799
rect 7403 16743 7459 16799
rect 7545 16743 7601 16799
rect 7687 16743 7743 16799
rect 7829 16743 7885 16799
rect 7971 16743 8027 16799
rect 8113 16743 8169 16799
rect 8255 16743 8311 16799
rect 8397 16743 8453 16799
rect 8539 16743 8595 16799
rect 8681 16743 8737 16799
rect 8823 16743 8879 16799
rect 8965 16743 9021 16799
rect 9107 16743 9163 16799
rect 9249 16743 9305 16799
rect 9391 16743 9447 16799
rect 9533 16743 9589 16799
rect 9675 16743 9731 16799
rect 9817 16743 9873 16799
rect 9959 16743 10015 16799
rect 10101 16743 10157 16799
rect 10243 16743 10299 16799
rect 10385 16743 10441 16799
rect 10527 16743 10583 16799
rect 10669 16743 10725 16799
rect 10811 16743 10867 16799
rect 10953 16743 11009 16799
rect 11095 16743 11151 16799
rect 11237 16743 11293 16799
rect 11379 16743 11435 16799
rect 11521 16743 11577 16799
rect 11663 16743 11719 16799
rect 11805 16743 11861 16799
rect 11947 16743 12003 16799
rect 12089 16743 12145 16799
rect 12231 16743 12287 16799
rect 12373 16743 12429 16799
rect 12515 16743 12571 16799
rect 12657 16743 12713 16799
rect 12799 16743 12855 16799
rect 12941 16743 12997 16799
rect 13083 16743 13139 16799
rect 13225 16743 13281 16799
rect 13367 16743 13423 16799
rect 13509 16743 13565 16799
rect 13651 16743 13707 16799
rect 13793 16743 13849 16799
rect 13935 16743 13991 16799
rect 14077 16743 14133 16799
rect 14219 16743 14275 16799
rect 14361 16743 14417 16799
rect 14503 16743 14559 16799
rect 14645 16743 14701 16799
rect 14787 16743 14843 16799
rect 161 16601 217 16657
rect 303 16601 359 16657
rect 445 16601 501 16657
rect 587 16601 643 16657
rect 729 16601 785 16657
rect 871 16601 927 16657
rect 1013 16601 1069 16657
rect 1155 16601 1211 16657
rect 1297 16601 1353 16657
rect 1439 16601 1495 16657
rect 1581 16601 1637 16657
rect 1723 16601 1779 16657
rect 1865 16601 1921 16657
rect 2007 16601 2063 16657
rect 2149 16601 2205 16657
rect 2291 16601 2347 16657
rect 2433 16601 2489 16657
rect 2575 16601 2631 16657
rect 2717 16601 2773 16657
rect 2859 16601 2915 16657
rect 3001 16601 3057 16657
rect 3143 16601 3199 16657
rect 3285 16601 3341 16657
rect 3427 16601 3483 16657
rect 3569 16601 3625 16657
rect 3711 16601 3767 16657
rect 3853 16601 3909 16657
rect 3995 16601 4051 16657
rect 4137 16601 4193 16657
rect 4279 16601 4335 16657
rect 4421 16601 4477 16657
rect 4563 16601 4619 16657
rect 4705 16601 4761 16657
rect 4847 16601 4903 16657
rect 4989 16601 5045 16657
rect 5131 16601 5187 16657
rect 5273 16601 5329 16657
rect 5415 16601 5471 16657
rect 5557 16601 5613 16657
rect 5699 16601 5755 16657
rect 5841 16601 5897 16657
rect 5983 16601 6039 16657
rect 6125 16601 6181 16657
rect 6267 16601 6323 16657
rect 6409 16601 6465 16657
rect 6551 16601 6607 16657
rect 6693 16601 6749 16657
rect 6835 16601 6891 16657
rect 6977 16601 7033 16657
rect 7119 16601 7175 16657
rect 7261 16601 7317 16657
rect 7403 16601 7459 16657
rect 7545 16601 7601 16657
rect 7687 16601 7743 16657
rect 7829 16601 7885 16657
rect 7971 16601 8027 16657
rect 8113 16601 8169 16657
rect 8255 16601 8311 16657
rect 8397 16601 8453 16657
rect 8539 16601 8595 16657
rect 8681 16601 8737 16657
rect 8823 16601 8879 16657
rect 8965 16601 9021 16657
rect 9107 16601 9163 16657
rect 9249 16601 9305 16657
rect 9391 16601 9447 16657
rect 9533 16601 9589 16657
rect 9675 16601 9731 16657
rect 9817 16601 9873 16657
rect 9959 16601 10015 16657
rect 10101 16601 10157 16657
rect 10243 16601 10299 16657
rect 10385 16601 10441 16657
rect 10527 16601 10583 16657
rect 10669 16601 10725 16657
rect 10811 16601 10867 16657
rect 10953 16601 11009 16657
rect 11095 16601 11151 16657
rect 11237 16601 11293 16657
rect 11379 16601 11435 16657
rect 11521 16601 11577 16657
rect 11663 16601 11719 16657
rect 11805 16601 11861 16657
rect 11947 16601 12003 16657
rect 12089 16601 12145 16657
rect 12231 16601 12287 16657
rect 12373 16601 12429 16657
rect 12515 16601 12571 16657
rect 12657 16601 12713 16657
rect 12799 16601 12855 16657
rect 12941 16601 12997 16657
rect 13083 16601 13139 16657
rect 13225 16601 13281 16657
rect 13367 16601 13423 16657
rect 13509 16601 13565 16657
rect 13651 16601 13707 16657
rect 13793 16601 13849 16657
rect 13935 16601 13991 16657
rect 14077 16601 14133 16657
rect 14219 16601 14275 16657
rect 14361 16601 14417 16657
rect 14503 16601 14559 16657
rect 14645 16601 14701 16657
rect 14787 16601 14843 16657
rect 161 16459 217 16515
rect 303 16459 359 16515
rect 445 16459 501 16515
rect 587 16459 643 16515
rect 729 16459 785 16515
rect 871 16459 927 16515
rect 1013 16459 1069 16515
rect 1155 16459 1211 16515
rect 1297 16459 1353 16515
rect 1439 16459 1495 16515
rect 1581 16459 1637 16515
rect 1723 16459 1779 16515
rect 1865 16459 1921 16515
rect 2007 16459 2063 16515
rect 2149 16459 2205 16515
rect 2291 16459 2347 16515
rect 2433 16459 2489 16515
rect 2575 16459 2631 16515
rect 2717 16459 2773 16515
rect 2859 16459 2915 16515
rect 3001 16459 3057 16515
rect 3143 16459 3199 16515
rect 3285 16459 3341 16515
rect 3427 16459 3483 16515
rect 3569 16459 3625 16515
rect 3711 16459 3767 16515
rect 3853 16459 3909 16515
rect 3995 16459 4051 16515
rect 4137 16459 4193 16515
rect 4279 16459 4335 16515
rect 4421 16459 4477 16515
rect 4563 16459 4619 16515
rect 4705 16459 4761 16515
rect 4847 16459 4903 16515
rect 4989 16459 5045 16515
rect 5131 16459 5187 16515
rect 5273 16459 5329 16515
rect 5415 16459 5471 16515
rect 5557 16459 5613 16515
rect 5699 16459 5755 16515
rect 5841 16459 5897 16515
rect 5983 16459 6039 16515
rect 6125 16459 6181 16515
rect 6267 16459 6323 16515
rect 6409 16459 6465 16515
rect 6551 16459 6607 16515
rect 6693 16459 6749 16515
rect 6835 16459 6891 16515
rect 6977 16459 7033 16515
rect 7119 16459 7175 16515
rect 7261 16459 7317 16515
rect 7403 16459 7459 16515
rect 7545 16459 7601 16515
rect 7687 16459 7743 16515
rect 7829 16459 7885 16515
rect 7971 16459 8027 16515
rect 8113 16459 8169 16515
rect 8255 16459 8311 16515
rect 8397 16459 8453 16515
rect 8539 16459 8595 16515
rect 8681 16459 8737 16515
rect 8823 16459 8879 16515
rect 8965 16459 9021 16515
rect 9107 16459 9163 16515
rect 9249 16459 9305 16515
rect 9391 16459 9447 16515
rect 9533 16459 9589 16515
rect 9675 16459 9731 16515
rect 9817 16459 9873 16515
rect 9959 16459 10015 16515
rect 10101 16459 10157 16515
rect 10243 16459 10299 16515
rect 10385 16459 10441 16515
rect 10527 16459 10583 16515
rect 10669 16459 10725 16515
rect 10811 16459 10867 16515
rect 10953 16459 11009 16515
rect 11095 16459 11151 16515
rect 11237 16459 11293 16515
rect 11379 16459 11435 16515
rect 11521 16459 11577 16515
rect 11663 16459 11719 16515
rect 11805 16459 11861 16515
rect 11947 16459 12003 16515
rect 12089 16459 12145 16515
rect 12231 16459 12287 16515
rect 12373 16459 12429 16515
rect 12515 16459 12571 16515
rect 12657 16459 12713 16515
rect 12799 16459 12855 16515
rect 12941 16459 12997 16515
rect 13083 16459 13139 16515
rect 13225 16459 13281 16515
rect 13367 16459 13423 16515
rect 13509 16459 13565 16515
rect 13651 16459 13707 16515
rect 13793 16459 13849 16515
rect 13935 16459 13991 16515
rect 14077 16459 14133 16515
rect 14219 16459 14275 16515
rect 14361 16459 14417 16515
rect 14503 16459 14559 16515
rect 14645 16459 14701 16515
rect 14787 16459 14843 16515
rect 161 16317 217 16373
rect 303 16317 359 16373
rect 445 16317 501 16373
rect 587 16317 643 16373
rect 729 16317 785 16373
rect 871 16317 927 16373
rect 1013 16317 1069 16373
rect 1155 16317 1211 16373
rect 1297 16317 1353 16373
rect 1439 16317 1495 16373
rect 1581 16317 1637 16373
rect 1723 16317 1779 16373
rect 1865 16317 1921 16373
rect 2007 16317 2063 16373
rect 2149 16317 2205 16373
rect 2291 16317 2347 16373
rect 2433 16317 2489 16373
rect 2575 16317 2631 16373
rect 2717 16317 2773 16373
rect 2859 16317 2915 16373
rect 3001 16317 3057 16373
rect 3143 16317 3199 16373
rect 3285 16317 3341 16373
rect 3427 16317 3483 16373
rect 3569 16317 3625 16373
rect 3711 16317 3767 16373
rect 3853 16317 3909 16373
rect 3995 16317 4051 16373
rect 4137 16317 4193 16373
rect 4279 16317 4335 16373
rect 4421 16317 4477 16373
rect 4563 16317 4619 16373
rect 4705 16317 4761 16373
rect 4847 16317 4903 16373
rect 4989 16317 5045 16373
rect 5131 16317 5187 16373
rect 5273 16317 5329 16373
rect 5415 16317 5471 16373
rect 5557 16317 5613 16373
rect 5699 16317 5755 16373
rect 5841 16317 5897 16373
rect 5983 16317 6039 16373
rect 6125 16317 6181 16373
rect 6267 16317 6323 16373
rect 6409 16317 6465 16373
rect 6551 16317 6607 16373
rect 6693 16317 6749 16373
rect 6835 16317 6891 16373
rect 6977 16317 7033 16373
rect 7119 16317 7175 16373
rect 7261 16317 7317 16373
rect 7403 16317 7459 16373
rect 7545 16317 7601 16373
rect 7687 16317 7743 16373
rect 7829 16317 7885 16373
rect 7971 16317 8027 16373
rect 8113 16317 8169 16373
rect 8255 16317 8311 16373
rect 8397 16317 8453 16373
rect 8539 16317 8595 16373
rect 8681 16317 8737 16373
rect 8823 16317 8879 16373
rect 8965 16317 9021 16373
rect 9107 16317 9163 16373
rect 9249 16317 9305 16373
rect 9391 16317 9447 16373
rect 9533 16317 9589 16373
rect 9675 16317 9731 16373
rect 9817 16317 9873 16373
rect 9959 16317 10015 16373
rect 10101 16317 10157 16373
rect 10243 16317 10299 16373
rect 10385 16317 10441 16373
rect 10527 16317 10583 16373
rect 10669 16317 10725 16373
rect 10811 16317 10867 16373
rect 10953 16317 11009 16373
rect 11095 16317 11151 16373
rect 11237 16317 11293 16373
rect 11379 16317 11435 16373
rect 11521 16317 11577 16373
rect 11663 16317 11719 16373
rect 11805 16317 11861 16373
rect 11947 16317 12003 16373
rect 12089 16317 12145 16373
rect 12231 16317 12287 16373
rect 12373 16317 12429 16373
rect 12515 16317 12571 16373
rect 12657 16317 12713 16373
rect 12799 16317 12855 16373
rect 12941 16317 12997 16373
rect 13083 16317 13139 16373
rect 13225 16317 13281 16373
rect 13367 16317 13423 16373
rect 13509 16317 13565 16373
rect 13651 16317 13707 16373
rect 13793 16317 13849 16373
rect 13935 16317 13991 16373
rect 14077 16317 14133 16373
rect 14219 16317 14275 16373
rect 14361 16317 14417 16373
rect 14503 16317 14559 16373
rect 14645 16317 14701 16373
rect 14787 16317 14843 16373
rect 161 16175 217 16231
rect 303 16175 359 16231
rect 445 16175 501 16231
rect 587 16175 643 16231
rect 729 16175 785 16231
rect 871 16175 927 16231
rect 1013 16175 1069 16231
rect 1155 16175 1211 16231
rect 1297 16175 1353 16231
rect 1439 16175 1495 16231
rect 1581 16175 1637 16231
rect 1723 16175 1779 16231
rect 1865 16175 1921 16231
rect 2007 16175 2063 16231
rect 2149 16175 2205 16231
rect 2291 16175 2347 16231
rect 2433 16175 2489 16231
rect 2575 16175 2631 16231
rect 2717 16175 2773 16231
rect 2859 16175 2915 16231
rect 3001 16175 3057 16231
rect 3143 16175 3199 16231
rect 3285 16175 3341 16231
rect 3427 16175 3483 16231
rect 3569 16175 3625 16231
rect 3711 16175 3767 16231
rect 3853 16175 3909 16231
rect 3995 16175 4051 16231
rect 4137 16175 4193 16231
rect 4279 16175 4335 16231
rect 4421 16175 4477 16231
rect 4563 16175 4619 16231
rect 4705 16175 4761 16231
rect 4847 16175 4903 16231
rect 4989 16175 5045 16231
rect 5131 16175 5187 16231
rect 5273 16175 5329 16231
rect 5415 16175 5471 16231
rect 5557 16175 5613 16231
rect 5699 16175 5755 16231
rect 5841 16175 5897 16231
rect 5983 16175 6039 16231
rect 6125 16175 6181 16231
rect 6267 16175 6323 16231
rect 6409 16175 6465 16231
rect 6551 16175 6607 16231
rect 6693 16175 6749 16231
rect 6835 16175 6891 16231
rect 6977 16175 7033 16231
rect 7119 16175 7175 16231
rect 7261 16175 7317 16231
rect 7403 16175 7459 16231
rect 7545 16175 7601 16231
rect 7687 16175 7743 16231
rect 7829 16175 7885 16231
rect 7971 16175 8027 16231
rect 8113 16175 8169 16231
rect 8255 16175 8311 16231
rect 8397 16175 8453 16231
rect 8539 16175 8595 16231
rect 8681 16175 8737 16231
rect 8823 16175 8879 16231
rect 8965 16175 9021 16231
rect 9107 16175 9163 16231
rect 9249 16175 9305 16231
rect 9391 16175 9447 16231
rect 9533 16175 9589 16231
rect 9675 16175 9731 16231
rect 9817 16175 9873 16231
rect 9959 16175 10015 16231
rect 10101 16175 10157 16231
rect 10243 16175 10299 16231
rect 10385 16175 10441 16231
rect 10527 16175 10583 16231
rect 10669 16175 10725 16231
rect 10811 16175 10867 16231
rect 10953 16175 11009 16231
rect 11095 16175 11151 16231
rect 11237 16175 11293 16231
rect 11379 16175 11435 16231
rect 11521 16175 11577 16231
rect 11663 16175 11719 16231
rect 11805 16175 11861 16231
rect 11947 16175 12003 16231
rect 12089 16175 12145 16231
rect 12231 16175 12287 16231
rect 12373 16175 12429 16231
rect 12515 16175 12571 16231
rect 12657 16175 12713 16231
rect 12799 16175 12855 16231
rect 12941 16175 12997 16231
rect 13083 16175 13139 16231
rect 13225 16175 13281 16231
rect 13367 16175 13423 16231
rect 13509 16175 13565 16231
rect 13651 16175 13707 16231
rect 13793 16175 13849 16231
rect 13935 16175 13991 16231
rect 14077 16175 14133 16231
rect 14219 16175 14275 16231
rect 14361 16175 14417 16231
rect 14503 16175 14559 16231
rect 14645 16175 14701 16231
rect 14787 16175 14843 16231
rect 161 16033 217 16089
rect 303 16033 359 16089
rect 445 16033 501 16089
rect 587 16033 643 16089
rect 729 16033 785 16089
rect 871 16033 927 16089
rect 1013 16033 1069 16089
rect 1155 16033 1211 16089
rect 1297 16033 1353 16089
rect 1439 16033 1495 16089
rect 1581 16033 1637 16089
rect 1723 16033 1779 16089
rect 1865 16033 1921 16089
rect 2007 16033 2063 16089
rect 2149 16033 2205 16089
rect 2291 16033 2347 16089
rect 2433 16033 2489 16089
rect 2575 16033 2631 16089
rect 2717 16033 2773 16089
rect 2859 16033 2915 16089
rect 3001 16033 3057 16089
rect 3143 16033 3199 16089
rect 3285 16033 3341 16089
rect 3427 16033 3483 16089
rect 3569 16033 3625 16089
rect 3711 16033 3767 16089
rect 3853 16033 3909 16089
rect 3995 16033 4051 16089
rect 4137 16033 4193 16089
rect 4279 16033 4335 16089
rect 4421 16033 4477 16089
rect 4563 16033 4619 16089
rect 4705 16033 4761 16089
rect 4847 16033 4903 16089
rect 4989 16033 5045 16089
rect 5131 16033 5187 16089
rect 5273 16033 5329 16089
rect 5415 16033 5471 16089
rect 5557 16033 5613 16089
rect 5699 16033 5755 16089
rect 5841 16033 5897 16089
rect 5983 16033 6039 16089
rect 6125 16033 6181 16089
rect 6267 16033 6323 16089
rect 6409 16033 6465 16089
rect 6551 16033 6607 16089
rect 6693 16033 6749 16089
rect 6835 16033 6891 16089
rect 6977 16033 7033 16089
rect 7119 16033 7175 16089
rect 7261 16033 7317 16089
rect 7403 16033 7459 16089
rect 7545 16033 7601 16089
rect 7687 16033 7743 16089
rect 7829 16033 7885 16089
rect 7971 16033 8027 16089
rect 8113 16033 8169 16089
rect 8255 16033 8311 16089
rect 8397 16033 8453 16089
rect 8539 16033 8595 16089
rect 8681 16033 8737 16089
rect 8823 16033 8879 16089
rect 8965 16033 9021 16089
rect 9107 16033 9163 16089
rect 9249 16033 9305 16089
rect 9391 16033 9447 16089
rect 9533 16033 9589 16089
rect 9675 16033 9731 16089
rect 9817 16033 9873 16089
rect 9959 16033 10015 16089
rect 10101 16033 10157 16089
rect 10243 16033 10299 16089
rect 10385 16033 10441 16089
rect 10527 16033 10583 16089
rect 10669 16033 10725 16089
rect 10811 16033 10867 16089
rect 10953 16033 11009 16089
rect 11095 16033 11151 16089
rect 11237 16033 11293 16089
rect 11379 16033 11435 16089
rect 11521 16033 11577 16089
rect 11663 16033 11719 16089
rect 11805 16033 11861 16089
rect 11947 16033 12003 16089
rect 12089 16033 12145 16089
rect 12231 16033 12287 16089
rect 12373 16033 12429 16089
rect 12515 16033 12571 16089
rect 12657 16033 12713 16089
rect 12799 16033 12855 16089
rect 12941 16033 12997 16089
rect 13083 16033 13139 16089
rect 13225 16033 13281 16089
rect 13367 16033 13423 16089
rect 13509 16033 13565 16089
rect 13651 16033 13707 16089
rect 13793 16033 13849 16089
rect 13935 16033 13991 16089
rect 14077 16033 14133 16089
rect 14219 16033 14275 16089
rect 14361 16033 14417 16089
rect 14503 16033 14559 16089
rect 14645 16033 14701 16089
rect 14787 16033 14843 16089
rect 161 15891 217 15947
rect 303 15891 359 15947
rect 445 15891 501 15947
rect 587 15891 643 15947
rect 729 15891 785 15947
rect 871 15891 927 15947
rect 1013 15891 1069 15947
rect 1155 15891 1211 15947
rect 1297 15891 1353 15947
rect 1439 15891 1495 15947
rect 1581 15891 1637 15947
rect 1723 15891 1779 15947
rect 1865 15891 1921 15947
rect 2007 15891 2063 15947
rect 2149 15891 2205 15947
rect 2291 15891 2347 15947
rect 2433 15891 2489 15947
rect 2575 15891 2631 15947
rect 2717 15891 2773 15947
rect 2859 15891 2915 15947
rect 3001 15891 3057 15947
rect 3143 15891 3199 15947
rect 3285 15891 3341 15947
rect 3427 15891 3483 15947
rect 3569 15891 3625 15947
rect 3711 15891 3767 15947
rect 3853 15891 3909 15947
rect 3995 15891 4051 15947
rect 4137 15891 4193 15947
rect 4279 15891 4335 15947
rect 4421 15891 4477 15947
rect 4563 15891 4619 15947
rect 4705 15891 4761 15947
rect 4847 15891 4903 15947
rect 4989 15891 5045 15947
rect 5131 15891 5187 15947
rect 5273 15891 5329 15947
rect 5415 15891 5471 15947
rect 5557 15891 5613 15947
rect 5699 15891 5755 15947
rect 5841 15891 5897 15947
rect 5983 15891 6039 15947
rect 6125 15891 6181 15947
rect 6267 15891 6323 15947
rect 6409 15891 6465 15947
rect 6551 15891 6607 15947
rect 6693 15891 6749 15947
rect 6835 15891 6891 15947
rect 6977 15891 7033 15947
rect 7119 15891 7175 15947
rect 7261 15891 7317 15947
rect 7403 15891 7459 15947
rect 7545 15891 7601 15947
rect 7687 15891 7743 15947
rect 7829 15891 7885 15947
rect 7971 15891 8027 15947
rect 8113 15891 8169 15947
rect 8255 15891 8311 15947
rect 8397 15891 8453 15947
rect 8539 15891 8595 15947
rect 8681 15891 8737 15947
rect 8823 15891 8879 15947
rect 8965 15891 9021 15947
rect 9107 15891 9163 15947
rect 9249 15891 9305 15947
rect 9391 15891 9447 15947
rect 9533 15891 9589 15947
rect 9675 15891 9731 15947
rect 9817 15891 9873 15947
rect 9959 15891 10015 15947
rect 10101 15891 10157 15947
rect 10243 15891 10299 15947
rect 10385 15891 10441 15947
rect 10527 15891 10583 15947
rect 10669 15891 10725 15947
rect 10811 15891 10867 15947
rect 10953 15891 11009 15947
rect 11095 15891 11151 15947
rect 11237 15891 11293 15947
rect 11379 15891 11435 15947
rect 11521 15891 11577 15947
rect 11663 15891 11719 15947
rect 11805 15891 11861 15947
rect 11947 15891 12003 15947
rect 12089 15891 12145 15947
rect 12231 15891 12287 15947
rect 12373 15891 12429 15947
rect 12515 15891 12571 15947
rect 12657 15891 12713 15947
rect 12799 15891 12855 15947
rect 12941 15891 12997 15947
rect 13083 15891 13139 15947
rect 13225 15891 13281 15947
rect 13367 15891 13423 15947
rect 13509 15891 13565 15947
rect 13651 15891 13707 15947
rect 13793 15891 13849 15947
rect 13935 15891 13991 15947
rect 14077 15891 14133 15947
rect 14219 15891 14275 15947
rect 14361 15891 14417 15947
rect 14503 15891 14559 15947
rect 14645 15891 14701 15947
rect 14787 15891 14843 15947
rect 161 15749 217 15805
rect 303 15749 359 15805
rect 445 15749 501 15805
rect 587 15749 643 15805
rect 729 15749 785 15805
rect 871 15749 927 15805
rect 1013 15749 1069 15805
rect 1155 15749 1211 15805
rect 1297 15749 1353 15805
rect 1439 15749 1495 15805
rect 1581 15749 1637 15805
rect 1723 15749 1779 15805
rect 1865 15749 1921 15805
rect 2007 15749 2063 15805
rect 2149 15749 2205 15805
rect 2291 15749 2347 15805
rect 2433 15749 2489 15805
rect 2575 15749 2631 15805
rect 2717 15749 2773 15805
rect 2859 15749 2915 15805
rect 3001 15749 3057 15805
rect 3143 15749 3199 15805
rect 3285 15749 3341 15805
rect 3427 15749 3483 15805
rect 3569 15749 3625 15805
rect 3711 15749 3767 15805
rect 3853 15749 3909 15805
rect 3995 15749 4051 15805
rect 4137 15749 4193 15805
rect 4279 15749 4335 15805
rect 4421 15749 4477 15805
rect 4563 15749 4619 15805
rect 4705 15749 4761 15805
rect 4847 15749 4903 15805
rect 4989 15749 5045 15805
rect 5131 15749 5187 15805
rect 5273 15749 5329 15805
rect 5415 15749 5471 15805
rect 5557 15749 5613 15805
rect 5699 15749 5755 15805
rect 5841 15749 5897 15805
rect 5983 15749 6039 15805
rect 6125 15749 6181 15805
rect 6267 15749 6323 15805
rect 6409 15749 6465 15805
rect 6551 15749 6607 15805
rect 6693 15749 6749 15805
rect 6835 15749 6891 15805
rect 6977 15749 7033 15805
rect 7119 15749 7175 15805
rect 7261 15749 7317 15805
rect 7403 15749 7459 15805
rect 7545 15749 7601 15805
rect 7687 15749 7743 15805
rect 7829 15749 7885 15805
rect 7971 15749 8027 15805
rect 8113 15749 8169 15805
rect 8255 15749 8311 15805
rect 8397 15749 8453 15805
rect 8539 15749 8595 15805
rect 8681 15749 8737 15805
rect 8823 15749 8879 15805
rect 8965 15749 9021 15805
rect 9107 15749 9163 15805
rect 9249 15749 9305 15805
rect 9391 15749 9447 15805
rect 9533 15749 9589 15805
rect 9675 15749 9731 15805
rect 9817 15749 9873 15805
rect 9959 15749 10015 15805
rect 10101 15749 10157 15805
rect 10243 15749 10299 15805
rect 10385 15749 10441 15805
rect 10527 15749 10583 15805
rect 10669 15749 10725 15805
rect 10811 15749 10867 15805
rect 10953 15749 11009 15805
rect 11095 15749 11151 15805
rect 11237 15749 11293 15805
rect 11379 15749 11435 15805
rect 11521 15749 11577 15805
rect 11663 15749 11719 15805
rect 11805 15749 11861 15805
rect 11947 15749 12003 15805
rect 12089 15749 12145 15805
rect 12231 15749 12287 15805
rect 12373 15749 12429 15805
rect 12515 15749 12571 15805
rect 12657 15749 12713 15805
rect 12799 15749 12855 15805
rect 12941 15749 12997 15805
rect 13083 15749 13139 15805
rect 13225 15749 13281 15805
rect 13367 15749 13423 15805
rect 13509 15749 13565 15805
rect 13651 15749 13707 15805
rect 13793 15749 13849 15805
rect 13935 15749 13991 15805
rect 14077 15749 14133 15805
rect 14219 15749 14275 15805
rect 14361 15749 14417 15805
rect 14503 15749 14559 15805
rect 14645 15749 14701 15805
rect 14787 15749 14843 15805
rect 161 15607 217 15663
rect 303 15607 359 15663
rect 445 15607 501 15663
rect 587 15607 643 15663
rect 729 15607 785 15663
rect 871 15607 927 15663
rect 1013 15607 1069 15663
rect 1155 15607 1211 15663
rect 1297 15607 1353 15663
rect 1439 15607 1495 15663
rect 1581 15607 1637 15663
rect 1723 15607 1779 15663
rect 1865 15607 1921 15663
rect 2007 15607 2063 15663
rect 2149 15607 2205 15663
rect 2291 15607 2347 15663
rect 2433 15607 2489 15663
rect 2575 15607 2631 15663
rect 2717 15607 2773 15663
rect 2859 15607 2915 15663
rect 3001 15607 3057 15663
rect 3143 15607 3199 15663
rect 3285 15607 3341 15663
rect 3427 15607 3483 15663
rect 3569 15607 3625 15663
rect 3711 15607 3767 15663
rect 3853 15607 3909 15663
rect 3995 15607 4051 15663
rect 4137 15607 4193 15663
rect 4279 15607 4335 15663
rect 4421 15607 4477 15663
rect 4563 15607 4619 15663
rect 4705 15607 4761 15663
rect 4847 15607 4903 15663
rect 4989 15607 5045 15663
rect 5131 15607 5187 15663
rect 5273 15607 5329 15663
rect 5415 15607 5471 15663
rect 5557 15607 5613 15663
rect 5699 15607 5755 15663
rect 5841 15607 5897 15663
rect 5983 15607 6039 15663
rect 6125 15607 6181 15663
rect 6267 15607 6323 15663
rect 6409 15607 6465 15663
rect 6551 15607 6607 15663
rect 6693 15607 6749 15663
rect 6835 15607 6891 15663
rect 6977 15607 7033 15663
rect 7119 15607 7175 15663
rect 7261 15607 7317 15663
rect 7403 15607 7459 15663
rect 7545 15607 7601 15663
rect 7687 15607 7743 15663
rect 7829 15607 7885 15663
rect 7971 15607 8027 15663
rect 8113 15607 8169 15663
rect 8255 15607 8311 15663
rect 8397 15607 8453 15663
rect 8539 15607 8595 15663
rect 8681 15607 8737 15663
rect 8823 15607 8879 15663
rect 8965 15607 9021 15663
rect 9107 15607 9163 15663
rect 9249 15607 9305 15663
rect 9391 15607 9447 15663
rect 9533 15607 9589 15663
rect 9675 15607 9731 15663
rect 9817 15607 9873 15663
rect 9959 15607 10015 15663
rect 10101 15607 10157 15663
rect 10243 15607 10299 15663
rect 10385 15607 10441 15663
rect 10527 15607 10583 15663
rect 10669 15607 10725 15663
rect 10811 15607 10867 15663
rect 10953 15607 11009 15663
rect 11095 15607 11151 15663
rect 11237 15607 11293 15663
rect 11379 15607 11435 15663
rect 11521 15607 11577 15663
rect 11663 15607 11719 15663
rect 11805 15607 11861 15663
rect 11947 15607 12003 15663
rect 12089 15607 12145 15663
rect 12231 15607 12287 15663
rect 12373 15607 12429 15663
rect 12515 15607 12571 15663
rect 12657 15607 12713 15663
rect 12799 15607 12855 15663
rect 12941 15607 12997 15663
rect 13083 15607 13139 15663
rect 13225 15607 13281 15663
rect 13367 15607 13423 15663
rect 13509 15607 13565 15663
rect 13651 15607 13707 15663
rect 13793 15607 13849 15663
rect 13935 15607 13991 15663
rect 14077 15607 14133 15663
rect 14219 15607 14275 15663
rect 14361 15607 14417 15663
rect 14503 15607 14559 15663
rect 14645 15607 14701 15663
rect 14787 15607 14843 15663
rect 161 15465 217 15521
rect 303 15465 359 15521
rect 445 15465 501 15521
rect 587 15465 643 15521
rect 729 15465 785 15521
rect 871 15465 927 15521
rect 1013 15465 1069 15521
rect 1155 15465 1211 15521
rect 1297 15465 1353 15521
rect 1439 15465 1495 15521
rect 1581 15465 1637 15521
rect 1723 15465 1779 15521
rect 1865 15465 1921 15521
rect 2007 15465 2063 15521
rect 2149 15465 2205 15521
rect 2291 15465 2347 15521
rect 2433 15465 2489 15521
rect 2575 15465 2631 15521
rect 2717 15465 2773 15521
rect 2859 15465 2915 15521
rect 3001 15465 3057 15521
rect 3143 15465 3199 15521
rect 3285 15465 3341 15521
rect 3427 15465 3483 15521
rect 3569 15465 3625 15521
rect 3711 15465 3767 15521
rect 3853 15465 3909 15521
rect 3995 15465 4051 15521
rect 4137 15465 4193 15521
rect 4279 15465 4335 15521
rect 4421 15465 4477 15521
rect 4563 15465 4619 15521
rect 4705 15465 4761 15521
rect 4847 15465 4903 15521
rect 4989 15465 5045 15521
rect 5131 15465 5187 15521
rect 5273 15465 5329 15521
rect 5415 15465 5471 15521
rect 5557 15465 5613 15521
rect 5699 15465 5755 15521
rect 5841 15465 5897 15521
rect 5983 15465 6039 15521
rect 6125 15465 6181 15521
rect 6267 15465 6323 15521
rect 6409 15465 6465 15521
rect 6551 15465 6607 15521
rect 6693 15465 6749 15521
rect 6835 15465 6891 15521
rect 6977 15465 7033 15521
rect 7119 15465 7175 15521
rect 7261 15465 7317 15521
rect 7403 15465 7459 15521
rect 7545 15465 7601 15521
rect 7687 15465 7743 15521
rect 7829 15465 7885 15521
rect 7971 15465 8027 15521
rect 8113 15465 8169 15521
rect 8255 15465 8311 15521
rect 8397 15465 8453 15521
rect 8539 15465 8595 15521
rect 8681 15465 8737 15521
rect 8823 15465 8879 15521
rect 8965 15465 9021 15521
rect 9107 15465 9163 15521
rect 9249 15465 9305 15521
rect 9391 15465 9447 15521
rect 9533 15465 9589 15521
rect 9675 15465 9731 15521
rect 9817 15465 9873 15521
rect 9959 15465 10015 15521
rect 10101 15465 10157 15521
rect 10243 15465 10299 15521
rect 10385 15465 10441 15521
rect 10527 15465 10583 15521
rect 10669 15465 10725 15521
rect 10811 15465 10867 15521
rect 10953 15465 11009 15521
rect 11095 15465 11151 15521
rect 11237 15465 11293 15521
rect 11379 15465 11435 15521
rect 11521 15465 11577 15521
rect 11663 15465 11719 15521
rect 11805 15465 11861 15521
rect 11947 15465 12003 15521
rect 12089 15465 12145 15521
rect 12231 15465 12287 15521
rect 12373 15465 12429 15521
rect 12515 15465 12571 15521
rect 12657 15465 12713 15521
rect 12799 15465 12855 15521
rect 12941 15465 12997 15521
rect 13083 15465 13139 15521
rect 13225 15465 13281 15521
rect 13367 15465 13423 15521
rect 13509 15465 13565 15521
rect 13651 15465 13707 15521
rect 13793 15465 13849 15521
rect 13935 15465 13991 15521
rect 14077 15465 14133 15521
rect 14219 15465 14275 15521
rect 14361 15465 14417 15521
rect 14503 15465 14559 15521
rect 14645 15465 14701 15521
rect 14787 15465 14843 15521
rect 161 15323 217 15379
rect 303 15323 359 15379
rect 445 15323 501 15379
rect 587 15323 643 15379
rect 729 15323 785 15379
rect 871 15323 927 15379
rect 1013 15323 1069 15379
rect 1155 15323 1211 15379
rect 1297 15323 1353 15379
rect 1439 15323 1495 15379
rect 1581 15323 1637 15379
rect 1723 15323 1779 15379
rect 1865 15323 1921 15379
rect 2007 15323 2063 15379
rect 2149 15323 2205 15379
rect 2291 15323 2347 15379
rect 2433 15323 2489 15379
rect 2575 15323 2631 15379
rect 2717 15323 2773 15379
rect 2859 15323 2915 15379
rect 3001 15323 3057 15379
rect 3143 15323 3199 15379
rect 3285 15323 3341 15379
rect 3427 15323 3483 15379
rect 3569 15323 3625 15379
rect 3711 15323 3767 15379
rect 3853 15323 3909 15379
rect 3995 15323 4051 15379
rect 4137 15323 4193 15379
rect 4279 15323 4335 15379
rect 4421 15323 4477 15379
rect 4563 15323 4619 15379
rect 4705 15323 4761 15379
rect 4847 15323 4903 15379
rect 4989 15323 5045 15379
rect 5131 15323 5187 15379
rect 5273 15323 5329 15379
rect 5415 15323 5471 15379
rect 5557 15323 5613 15379
rect 5699 15323 5755 15379
rect 5841 15323 5897 15379
rect 5983 15323 6039 15379
rect 6125 15323 6181 15379
rect 6267 15323 6323 15379
rect 6409 15323 6465 15379
rect 6551 15323 6607 15379
rect 6693 15323 6749 15379
rect 6835 15323 6891 15379
rect 6977 15323 7033 15379
rect 7119 15323 7175 15379
rect 7261 15323 7317 15379
rect 7403 15323 7459 15379
rect 7545 15323 7601 15379
rect 7687 15323 7743 15379
rect 7829 15323 7885 15379
rect 7971 15323 8027 15379
rect 8113 15323 8169 15379
rect 8255 15323 8311 15379
rect 8397 15323 8453 15379
rect 8539 15323 8595 15379
rect 8681 15323 8737 15379
rect 8823 15323 8879 15379
rect 8965 15323 9021 15379
rect 9107 15323 9163 15379
rect 9249 15323 9305 15379
rect 9391 15323 9447 15379
rect 9533 15323 9589 15379
rect 9675 15323 9731 15379
rect 9817 15323 9873 15379
rect 9959 15323 10015 15379
rect 10101 15323 10157 15379
rect 10243 15323 10299 15379
rect 10385 15323 10441 15379
rect 10527 15323 10583 15379
rect 10669 15323 10725 15379
rect 10811 15323 10867 15379
rect 10953 15323 11009 15379
rect 11095 15323 11151 15379
rect 11237 15323 11293 15379
rect 11379 15323 11435 15379
rect 11521 15323 11577 15379
rect 11663 15323 11719 15379
rect 11805 15323 11861 15379
rect 11947 15323 12003 15379
rect 12089 15323 12145 15379
rect 12231 15323 12287 15379
rect 12373 15323 12429 15379
rect 12515 15323 12571 15379
rect 12657 15323 12713 15379
rect 12799 15323 12855 15379
rect 12941 15323 12997 15379
rect 13083 15323 13139 15379
rect 13225 15323 13281 15379
rect 13367 15323 13423 15379
rect 13509 15323 13565 15379
rect 13651 15323 13707 15379
rect 13793 15323 13849 15379
rect 13935 15323 13991 15379
rect 14077 15323 14133 15379
rect 14219 15323 14275 15379
rect 14361 15323 14417 15379
rect 14503 15323 14559 15379
rect 14645 15323 14701 15379
rect 14787 15323 14843 15379
rect 161 15181 217 15237
rect 303 15181 359 15237
rect 445 15181 501 15237
rect 587 15181 643 15237
rect 729 15181 785 15237
rect 871 15181 927 15237
rect 1013 15181 1069 15237
rect 1155 15181 1211 15237
rect 1297 15181 1353 15237
rect 1439 15181 1495 15237
rect 1581 15181 1637 15237
rect 1723 15181 1779 15237
rect 1865 15181 1921 15237
rect 2007 15181 2063 15237
rect 2149 15181 2205 15237
rect 2291 15181 2347 15237
rect 2433 15181 2489 15237
rect 2575 15181 2631 15237
rect 2717 15181 2773 15237
rect 2859 15181 2915 15237
rect 3001 15181 3057 15237
rect 3143 15181 3199 15237
rect 3285 15181 3341 15237
rect 3427 15181 3483 15237
rect 3569 15181 3625 15237
rect 3711 15181 3767 15237
rect 3853 15181 3909 15237
rect 3995 15181 4051 15237
rect 4137 15181 4193 15237
rect 4279 15181 4335 15237
rect 4421 15181 4477 15237
rect 4563 15181 4619 15237
rect 4705 15181 4761 15237
rect 4847 15181 4903 15237
rect 4989 15181 5045 15237
rect 5131 15181 5187 15237
rect 5273 15181 5329 15237
rect 5415 15181 5471 15237
rect 5557 15181 5613 15237
rect 5699 15181 5755 15237
rect 5841 15181 5897 15237
rect 5983 15181 6039 15237
rect 6125 15181 6181 15237
rect 6267 15181 6323 15237
rect 6409 15181 6465 15237
rect 6551 15181 6607 15237
rect 6693 15181 6749 15237
rect 6835 15181 6891 15237
rect 6977 15181 7033 15237
rect 7119 15181 7175 15237
rect 7261 15181 7317 15237
rect 7403 15181 7459 15237
rect 7545 15181 7601 15237
rect 7687 15181 7743 15237
rect 7829 15181 7885 15237
rect 7971 15181 8027 15237
rect 8113 15181 8169 15237
rect 8255 15181 8311 15237
rect 8397 15181 8453 15237
rect 8539 15181 8595 15237
rect 8681 15181 8737 15237
rect 8823 15181 8879 15237
rect 8965 15181 9021 15237
rect 9107 15181 9163 15237
rect 9249 15181 9305 15237
rect 9391 15181 9447 15237
rect 9533 15181 9589 15237
rect 9675 15181 9731 15237
rect 9817 15181 9873 15237
rect 9959 15181 10015 15237
rect 10101 15181 10157 15237
rect 10243 15181 10299 15237
rect 10385 15181 10441 15237
rect 10527 15181 10583 15237
rect 10669 15181 10725 15237
rect 10811 15181 10867 15237
rect 10953 15181 11009 15237
rect 11095 15181 11151 15237
rect 11237 15181 11293 15237
rect 11379 15181 11435 15237
rect 11521 15181 11577 15237
rect 11663 15181 11719 15237
rect 11805 15181 11861 15237
rect 11947 15181 12003 15237
rect 12089 15181 12145 15237
rect 12231 15181 12287 15237
rect 12373 15181 12429 15237
rect 12515 15181 12571 15237
rect 12657 15181 12713 15237
rect 12799 15181 12855 15237
rect 12941 15181 12997 15237
rect 13083 15181 13139 15237
rect 13225 15181 13281 15237
rect 13367 15181 13423 15237
rect 13509 15181 13565 15237
rect 13651 15181 13707 15237
rect 13793 15181 13849 15237
rect 13935 15181 13991 15237
rect 14077 15181 14133 15237
rect 14219 15181 14275 15237
rect 14361 15181 14417 15237
rect 14503 15181 14559 15237
rect 14645 15181 14701 15237
rect 14787 15181 14843 15237
rect 161 15039 217 15095
rect 303 15039 359 15095
rect 445 15039 501 15095
rect 587 15039 643 15095
rect 729 15039 785 15095
rect 871 15039 927 15095
rect 1013 15039 1069 15095
rect 1155 15039 1211 15095
rect 1297 15039 1353 15095
rect 1439 15039 1495 15095
rect 1581 15039 1637 15095
rect 1723 15039 1779 15095
rect 1865 15039 1921 15095
rect 2007 15039 2063 15095
rect 2149 15039 2205 15095
rect 2291 15039 2347 15095
rect 2433 15039 2489 15095
rect 2575 15039 2631 15095
rect 2717 15039 2773 15095
rect 2859 15039 2915 15095
rect 3001 15039 3057 15095
rect 3143 15039 3199 15095
rect 3285 15039 3341 15095
rect 3427 15039 3483 15095
rect 3569 15039 3625 15095
rect 3711 15039 3767 15095
rect 3853 15039 3909 15095
rect 3995 15039 4051 15095
rect 4137 15039 4193 15095
rect 4279 15039 4335 15095
rect 4421 15039 4477 15095
rect 4563 15039 4619 15095
rect 4705 15039 4761 15095
rect 4847 15039 4903 15095
rect 4989 15039 5045 15095
rect 5131 15039 5187 15095
rect 5273 15039 5329 15095
rect 5415 15039 5471 15095
rect 5557 15039 5613 15095
rect 5699 15039 5755 15095
rect 5841 15039 5897 15095
rect 5983 15039 6039 15095
rect 6125 15039 6181 15095
rect 6267 15039 6323 15095
rect 6409 15039 6465 15095
rect 6551 15039 6607 15095
rect 6693 15039 6749 15095
rect 6835 15039 6891 15095
rect 6977 15039 7033 15095
rect 7119 15039 7175 15095
rect 7261 15039 7317 15095
rect 7403 15039 7459 15095
rect 7545 15039 7601 15095
rect 7687 15039 7743 15095
rect 7829 15039 7885 15095
rect 7971 15039 8027 15095
rect 8113 15039 8169 15095
rect 8255 15039 8311 15095
rect 8397 15039 8453 15095
rect 8539 15039 8595 15095
rect 8681 15039 8737 15095
rect 8823 15039 8879 15095
rect 8965 15039 9021 15095
rect 9107 15039 9163 15095
rect 9249 15039 9305 15095
rect 9391 15039 9447 15095
rect 9533 15039 9589 15095
rect 9675 15039 9731 15095
rect 9817 15039 9873 15095
rect 9959 15039 10015 15095
rect 10101 15039 10157 15095
rect 10243 15039 10299 15095
rect 10385 15039 10441 15095
rect 10527 15039 10583 15095
rect 10669 15039 10725 15095
rect 10811 15039 10867 15095
rect 10953 15039 11009 15095
rect 11095 15039 11151 15095
rect 11237 15039 11293 15095
rect 11379 15039 11435 15095
rect 11521 15039 11577 15095
rect 11663 15039 11719 15095
rect 11805 15039 11861 15095
rect 11947 15039 12003 15095
rect 12089 15039 12145 15095
rect 12231 15039 12287 15095
rect 12373 15039 12429 15095
rect 12515 15039 12571 15095
rect 12657 15039 12713 15095
rect 12799 15039 12855 15095
rect 12941 15039 12997 15095
rect 13083 15039 13139 15095
rect 13225 15039 13281 15095
rect 13367 15039 13423 15095
rect 13509 15039 13565 15095
rect 13651 15039 13707 15095
rect 13793 15039 13849 15095
rect 13935 15039 13991 15095
rect 14077 15039 14133 15095
rect 14219 15039 14275 15095
rect 14361 15039 14417 15095
rect 14503 15039 14559 15095
rect 14645 15039 14701 15095
rect 14787 15039 14843 15095
rect 161 14897 217 14953
rect 303 14897 359 14953
rect 445 14897 501 14953
rect 587 14897 643 14953
rect 729 14897 785 14953
rect 871 14897 927 14953
rect 1013 14897 1069 14953
rect 1155 14897 1211 14953
rect 1297 14897 1353 14953
rect 1439 14897 1495 14953
rect 1581 14897 1637 14953
rect 1723 14897 1779 14953
rect 1865 14897 1921 14953
rect 2007 14897 2063 14953
rect 2149 14897 2205 14953
rect 2291 14897 2347 14953
rect 2433 14897 2489 14953
rect 2575 14897 2631 14953
rect 2717 14897 2773 14953
rect 2859 14897 2915 14953
rect 3001 14897 3057 14953
rect 3143 14897 3199 14953
rect 3285 14897 3341 14953
rect 3427 14897 3483 14953
rect 3569 14897 3625 14953
rect 3711 14897 3767 14953
rect 3853 14897 3909 14953
rect 3995 14897 4051 14953
rect 4137 14897 4193 14953
rect 4279 14897 4335 14953
rect 4421 14897 4477 14953
rect 4563 14897 4619 14953
rect 4705 14897 4761 14953
rect 4847 14897 4903 14953
rect 4989 14897 5045 14953
rect 5131 14897 5187 14953
rect 5273 14897 5329 14953
rect 5415 14897 5471 14953
rect 5557 14897 5613 14953
rect 5699 14897 5755 14953
rect 5841 14897 5897 14953
rect 5983 14897 6039 14953
rect 6125 14897 6181 14953
rect 6267 14897 6323 14953
rect 6409 14897 6465 14953
rect 6551 14897 6607 14953
rect 6693 14897 6749 14953
rect 6835 14897 6891 14953
rect 6977 14897 7033 14953
rect 7119 14897 7175 14953
rect 7261 14897 7317 14953
rect 7403 14897 7459 14953
rect 7545 14897 7601 14953
rect 7687 14897 7743 14953
rect 7829 14897 7885 14953
rect 7971 14897 8027 14953
rect 8113 14897 8169 14953
rect 8255 14897 8311 14953
rect 8397 14897 8453 14953
rect 8539 14897 8595 14953
rect 8681 14897 8737 14953
rect 8823 14897 8879 14953
rect 8965 14897 9021 14953
rect 9107 14897 9163 14953
rect 9249 14897 9305 14953
rect 9391 14897 9447 14953
rect 9533 14897 9589 14953
rect 9675 14897 9731 14953
rect 9817 14897 9873 14953
rect 9959 14897 10015 14953
rect 10101 14897 10157 14953
rect 10243 14897 10299 14953
rect 10385 14897 10441 14953
rect 10527 14897 10583 14953
rect 10669 14897 10725 14953
rect 10811 14897 10867 14953
rect 10953 14897 11009 14953
rect 11095 14897 11151 14953
rect 11237 14897 11293 14953
rect 11379 14897 11435 14953
rect 11521 14897 11577 14953
rect 11663 14897 11719 14953
rect 11805 14897 11861 14953
rect 11947 14897 12003 14953
rect 12089 14897 12145 14953
rect 12231 14897 12287 14953
rect 12373 14897 12429 14953
rect 12515 14897 12571 14953
rect 12657 14897 12713 14953
rect 12799 14897 12855 14953
rect 12941 14897 12997 14953
rect 13083 14897 13139 14953
rect 13225 14897 13281 14953
rect 13367 14897 13423 14953
rect 13509 14897 13565 14953
rect 13651 14897 13707 14953
rect 13793 14897 13849 14953
rect 13935 14897 13991 14953
rect 14077 14897 14133 14953
rect 14219 14897 14275 14953
rect 14361 14897 14417 14953
rect 14503 14897 14559 14953
rect 14645 14897 14701 14953
rect 14787 14897 14843 14953
rect 161 14755 217 14811
rect 303 14755 359 14811
rect 445 14755 501 14811
rect 587 14755 643 14811
rect 729 14755 785 14811
rect 871 14755 927 14811
rect 1013 14755 1069 14811
rect 1155 14755 1211 14811
rect 1297 14755 1353 14811
rect 1439 14755 1495 14811
rect 1581 14755 1637 14811
rect 1723 14755 1779 14811
rect 1865 14755 1921 14811
rect 2007 14755 2063 14811
rect 2149 14755 2205 14811
rect 2291 14755 2347 14811
rect 2433 14755 2489 14811
rect 2575 14755 2631 14811
rect 2717 14755 2773 14811
rect 2859 14755 2915 14811
rect 3001 14755 3057 14811
rect 3143 14755 3199 14811
rect 3285 14755 3341 14811
rect 3427 14755 3483 14811
rect 3569 14755 3625 14811
rect 3711 14755 3767 14811
rect 3853 14755 3909 14811
rect 3995 14755 4051 14811
rect 4137 14755 4193 14811
rect 4279 14755 4335 14811
rect 4421 14755 4477 14811
rect 4563 14755 4619 14811
rect 4705 14755 4761 14811
rect 4847 14755 4903 14811
rect 4989 14755 5045 14811
rect 5131 14755 5187 14811
rect 5273 14755 5329 14811
rect 5415 14755 5471 14811
rect 5557 14755 5613 14811
rect 5699 14755 5755 14811
rect 5841 14755 5897 14811
rect 5983 14755 6039 14811
rect 6125 14755 6181 14811
rect 6267 14755 6323 14811
rect 6409 14755 6465 14811
rect 6551 14755 6607 14811
rect 6693 14755 6749 14811
rect 6835 14755 6891 14811
rect 6977 14755 7033 14811
rect 7119 14755 7175 14811
rect 7261 14755 7317 14811
rect 7403 14755 7459 14811
rect 7545 14755 7601 14811
rect 7687 14755 7743 14811
rect 7829 14755 7885 14811
rect 7971 14755 8027 14811
rect 8113 14755 8169 14811
rect 8255 14755 8311 14811
rect 8397 14755 8453 14811
rect 8539 14755 8595 14811
rect 8681 14755 8737 14811
rect 8823 14755 8879 14811
rect 8965 14755 9021 14811
rect 9107 14755 9163 14811
rect 9249 14755 9305 14811
rect 9391 14755 9447 14811
rect 9533 14755 9589 14811
rect 9675 14755 9731 14811
rect 9817 14755 9873 14811
rect 9959 14755 10015 14811
rect 10101 14755 10157 14811
rect 10243 14755 10299 14811
rect 10385 14755 10441 14811
rect 10527 14755 10583 14811
rect 10669 14755 10725 14811
rect 10811 14755 10867 14811
rect 10953 14755 11009 14811
rect 11095 14755 11151 14811
rect 11237 14755 11293 14811
rect 11379 14755 11435 14811
rect 11521 14755 11577 14811
rect 11663 14755 11719 14811
rect 11805 14755 11861 14811
rect 11947 14755 12003 14811
rect 12089 14755 12145 14811
rect 12231 14755 12287 14811
rect 12373 14755 12429 14811
rect 12515 14755 12571 14811
rect 12657 14755 12713 14811
rect 12799 14755 12855 14811
rect 12941 14755 12997 14811
rect 13083 14755 13139 14811
rect 13225 14755 13281 14811
rect 13367 14755 13423 14811
rect 13509 14755 13565 14811
rect 13651 14755 13707 14811
rect 13793 14755 13849 14811
rect 13935 14755 13991 14811
rect 14077 14755 14133 14811
rect 14219 14755 14275 14811
rect 14361 14755 14417 14811
rect 14503 14755 14559 14811
rect 14645 14755 14701 14811
rect 14787 14755 14843 14811
rect 161 14613 217 14669
rect 303 14613 359 14669
rect 445 14613 501 14669
rect 587 14613 643 14669
rect 729 14613 785 14669
rect 871 14613 927 14669
rect 1013 14613 1069 14669
rect 1155 14613 1211 14669
rect 1297 14613 1353 14669
rect 1439 14613 1495 14669
rect 1581 14613 1637 14669
rect 1723 14613 1779 14669
rect 1865 14613 1921 14669
rect 2007 14613 2063 14669
rect 2149 14613 2205 14669
rect 2291 14613 2347 14669
rect 2433 14613 2489 14669
rect 2575 14613 2631 14669
rect 2717 14613 2773 14669
rect 2859 14613 2915 14669
rect 3001 14613 3057 14669
rect 3143 14613 3199 14669
rect 3285 14613 3341 14669
rect 3427 14613 3483 14669
rect 3569 14613 3625 14669
rect 3711 14613 3767 14669
rect 3853 14613 3909 14669
rect 3995 14613 4051 14669
rect 4137 14613 4193 14669
rect 4279 14613 4335 14669
rect 4421 14613 4477 14669
rect 4563 14613 4619 14669
rect 4705 14613 4761 14669
rect 4847 14613 4903 14669
rect 4989 14613 5045 14669
rect 5131 14613 5187 14669
rect 5273 14613 5329 14669
rect 5415 14613 5471 14669
rect 5557 14613 5613 14669
rect 5699 14613 5755 14669
rect 5841 14613 5897 14669
rect 5983 14613 6039 14669
rect 6125 14613 6181 14669
rect 6267 14613 6323 14669
rect 6409 14613 6465 14669
rect 6551 14613 6607 14669
rect 6693 14613 6749 14669
rect 6835 14613 6891 14669
rect 6977 14613 7033 14669
rect 7119 14613 7175 14669
rect 7261 14613 7317 14669
rect 7403 14613 7459 14669
rect 7545 14613 7601 14669
rect 7687 14613 7743 14669
rect 7829 14613 7885 14669
rect 7971 14613 8027 14669
rect 8113 14613 8169 14669
rect 8255 14613 8311 14669
rect 8397 14613 8453 14669
rect 8539 14613 8595 14669
rect 8681 14613 8737 14669
rect 8823 14613 8879 14669
rect 8965 14613 9021 14669
rect 9107 14613 9163 14669
rect 9249 14613 9305 14669
rect 9391 14613 9447 14669
rect 9533 14613 9589 14669
rect 9675 14613 9731 14669
rect 9817 14613 9873 14669
rect 9959 14613 10015 14669
rect 10101 14613 10157 14669
rect 10243 14613 10299 14669
rect 10385 14613 10441 14669
rect 10527 14613 10583 14669
rect 10669 14613 10725 14669
rect 10811 14613 10867 14669
rect 10953 14613 11009 14669
rect 11095 14613 11151 14669
rect 11237 14613 11293 14669
rect 11379 14613 11435 14669
rect 11521 14613 11577 14669
rect 11663 14613 11719 14669
rect 11805 14613 11861 14669
rect 11947 14613 12003 14669
rect 12089 14613 12145 14669
rect 12231 14613 12287 14669
rect 12373 14613 12429 14669
rect 12515 14613 12571 14669
rect 12657 14613 12713 14669
rect 12799 14613 12855 14669
rect 12941 14613 12997 14669
rect 13083 14613 13139 14669
rect 13225 14613 13281 14669
rect 13367 14613 13423 14669
rect 13509 14613 13565 14669
rect 13651 14613 13707 14669
rect 13793 14613 13849 14669
rect 13935 14613 13991 14669
rect 14077 14613 14133 14669
rect 14219 14613 14275 14669
rect 14361 14613 14417 14669
rect 14503 14613 14559 14669
rect 14645 14613 14701 14669
rect 14787 14613 14843 14669
rect 161 14471 217 14527
rect 303 14471 359 14527
rect 445 14471 501 14527
rect 587 14471 643 14527
rect 729 14471 785 14527
rect 871 14471 927 14527
rect 1013 14471 1069 14527
rect 1155 14471 1211 14527
rect 1297 14471 1353 14527
rect 1439 14471 1495 14527
rect 1581 14471 1637 14527
rect 1723 14471 1779 14527
rect 1865 14471 1921 14527
rect 2007 14471 2063 14527
rect 2149 14471 2205 14527
rect 2291 14471 2347 14527
rect 2433 14471 2489 14527
rect 2575 14471 2631 14527
rect 2717 14471 2773 14527
rect 2859 14471 2915 14527
rect 3001 14471 3057 14527
rect 3143 14471 3199 14527
rect 3285 14471 3341 14527
rect 3427 14471 3483 14527
rect 3569 14471 3625 14527
rect 3711 14471 3767 14527
rect 3853 14471 3909 14527
rect 3995 14471 4051 14527
rect 4137 14471 4193 14527
rect 4279 14471 4335 14527
rect 4421 14471 4477 14527
rect 4563 14471 4619 14527
rect 4705 14471 4761 14527
rect 4847 14471 4903 14527
rect 4989 14471 5045 14527
rect 5131 14471 5187 14527
rect 5273 14471 5329 14527
rect 5415 14471 5471 14527
rect 5557 14471 5613 14527
rect 5699 14471 5755 14527
rect 5841 14471 5897 14527
rect 5983 14471 6039 14527
rect 6125 14471 6181 14527
rect 6267 14471 6323 14527
rect 6409 14471 6465 14527
rect 6551 14471 6607 14527
rect 6693 14471 6749 14527
rect 6835 14471 6891 14527
rect 6977 14471 7033 14527
rect 7119 14471 7175 14527
rect 7261 14471 7317 14527
rect 7403 14471 7459 14527
rect 7545 14471 7601 14527
rect 7687 14471 7743 14527
rect 7829 14471 7885 14527
rect 7971 14471 8027 14527
rect 8113 14471 8169 14527
rect 8255 14471 8311 14527
rect 8397 14471 8453 14527
rect 8539 14471 8595 14527
rect 8681 14471 8737 14527
rect 8823 14471 8879 14527
rect 8965 14471 9021 14527
rect 9107 14471 9163 14527
rect 9249 14471 9305 14527
rect 9391 14471 9447 14527
rect 9533 14471 9589 14527
rect 9675 14471 9731 14527
rect 9817 14471 9873 14527
rect 9959 14471 10015 14527
rect 10101 14471 10157 14527
rect 10243 14471 10299 14527
rect 10385 14471 10441 14527
rect 10527 14471 10583 14527
rect 10669 14471 10725 14527
rect 10811 14471 10867 14527
rect 10953 14471 11009 14527
rect 11095 14471 11151 14527
rect 11237 14471 11293 14527
rect 11379 14471 11435 14527
rect 11521 14471 11577 14527
rect 11663 14471 11719 14527
rect 11805 14471 11861 14527
rect 11947 14471 12003 14527
rect 12089 14471 12145 14527
rect 12231 14471 12287 14527
rect 12373 14471 12429 14527
rect 12515 14471 12571 14527
rect 12657 14471 12713 14527
rect 12799 14471 12855 14527
rect 12941 14471 12997 14527
rect 13083 14471 13139 14527
rect 13225 14471 13281 14527
rect 13367 14471 13423 14527
rect 13509 14471 13565 14527
rect 13651 14471 13707 14527
rect 13793 14471 13849 14527
rect 13935 14471 13991 14527
rect 14077 14471 14133 14527
rect 14219 14471 14275 14527
rect 14361 14471 14417 14527
rect 14503 14471 14559 14527
rect 14645 14471 14701 14527
rect 14787 14471 14843 14527
rect 161 14329 217 14385
rect 303 14329 359 14385
rect 445 14329 501 14385
rect 587 14329 643 14385
rect 729 14329 785 14385
rect 871 14329 927 14385
rect 1013 14329 1069 14385
rect 1155 14329 1211 14385
rect 1297 14329 1353 14385
rect 1439 14329 1495 14385
rect 1581 14329 1637 14385
rect 1723 14329 1779 14385
rect 1865 14329 1921 14385
rect 2007 14329 2063 14385
rect 2149 14329 2205 14385
rect 2291 14329 2347 14385
rect 2433 14329 2489 14385
rect 2575 14329 2631 14385
rect 2717 14329 2773 14385
rect 2859 14329 2915 14385
rect 3001 14329 3057 14385
rect 3143 14329 3199 14385
rect 3285 14329 3341 14385
rect 3427 14329 3483 14385
rect 3569 14329 3625 14385
rect 3711 14329 3767 14385
rect 3853 14329 3909 14385
rect 3995 14329 4051 14385
rect 4137 14329 4193 14385
rect 4279 14329 4335 14385
rect 4421 14329 4477 14385
rect 4563 14329 4619 14385
rect 4705 14329 4761 14385
rect 4847 14329 4903 14385
rect 4989 14329 5045 14385
rect 5131 14329 5187 14385
rect 5273 14329 5329 14385
rect 5415 14329 5471 14385
rect 5557 14329 5613 14385
rect 5699 14329 5755 14385
rect 5841 14329 5897 14385
rect 5983 14329 6039 14385
rect 6125 14329 6181 14385
rect 6267 14329 6323 14385
rect 6409 14329 6465 14385
rect 6551 14329 6607 14385
rect 6693 14329 6749 14385
rect 6835 14329 6891 14385
rect 6977 14329 7033 14385
rect 7119 14329 7175 14385
rect 7261 14329 7317 14385
rect 7403 14329 7459 14385
rect 7545 14329 7601 14385
rect 7687 14329 7743 14385
rect 7829 14329 7885 14385
rect 7971 14329 8027 14385
rect 8113 14329 8169 14385
rect 8255 14329 8311 14385
rect 8397 14329 8453 14385
rect 8539 14329 8595 14385
rect 8681 14329 8737 14385
rect 8823 14329 8879 14385
rect 8965 14329 9021 14385
rect 9107 14329 9163 14385
rect 9249 14329 9305 14385
rect 9391 14329 9447 14385
rect 9533 14329 9589 14385
rect 9675 14329 9731 14385
rect 9817 14329 9873 14385
rect 9959 14329 10015 14385
rect 10101 14329 10157 14385
rect 10243 14329 10299 14385
rect 10385 14329 10441 14385
rect 10527 14329 10583 14385
rect 10669 14329 10725 14385
rect 10811 14329 10867 14385
rect 10953 14329 11009 14385
rect 11095 14329 11151 14385
rect 11237 14329 11293 14385
rect 11379 14329 11435 14385
rect 11521 14329 11577 14385
rect 11663 14329 11719 14385
rect 11805 14329 11861 14385
rect 11947 14329 12003 14385
rect 12089 14329 12145 14385
rect 12231 14329 12287 14385
rect 12373 14329 12429 14385
rect 12515 14329 12571 14385
rect 12657 14329 12713 14385
rect 12799 14329 12855 14385
rect 12941 14329 12997 14385
rect 13083 14329 13139 14385
rect 13225 14329 13281 14385
rect 13367 14329 13423 14385
rect 13509 14329 13565 14385
rect 13651 14329 13707 14385
rect 13793 14329 13849 14385
rect 13935 14329 13991 14385
rect 14077 14329 14133 14385
rect 14219 14329 14275 14385
rect 14361 14329 14417 14385
rect 14503 14329 14559 14385
rect 14645 14329 14701 14385
rect 14787 14329 14843 14385
rect 161 14187 217 14243
rect 303 14187 359 14243
rect 445 14187 501 14243
rect 587 14187 643 14243
rect 729 14187 785 14243
rect 871 14187 927 14243
rect 1013 14187 1069 14243
rect 1155 14187 1211 14243
rect 1297 14187 1353 14243
rect 1439 14187 1495 14243
rect 1581 14187 1637 14243
rect 1723 14187 1779 14243
rect 1865 14187 1921 14243
rect 2007 14187 2063 14243
rect 2149 14187 2205 14243
rect 2291 14187 2347 14243
rect 2433 14187 2489 14243
rect 2575 14187 2631 14243
rect 2717 14187 2773 14243
rect 2859 14187 2915 14243
rect 3001 14187 3057 14243
rect 3143 14187 3199 14243
rect 3285 14187 3341 14243
rect 3427 14187 3483 14243
rect 3569 14187 3625 14243
rect 3711 14187 3767 14243
rect 3853 14187 3909 14243
rect 3995 14187 4051 14243
rect 4137 14187 4193 14243
rect 4279 14187 4335 14243
rect 4421 14187 4477 14243
rect 4563 14187 4619 14243
rect 4705 14187 4761 14243
rect 4847 14187 4903 14243
rect 4989 14187 5045 14243
rect 5131 14187 5187 14243
rect 5273 14187 5329 14243
rect 5415 14187 5471 14243
rect 5557 14187 5613 14243
rect 5699 14187 5755 14243
rect 5841 14187 5897 14243
rect 5983 14187 6039 14243
rect 6125 14187 6181 14243
rect 6267 14187 6323 14243
rect 6409 14187 6465 14243
rect 6551 14187 6607 14243
rect 6693 14187 6749 14243
rect 6835 14187 6891 14243
rect 6977 14187 7033 14243
rect 7119 14187 7175 14243
rect 7261 14187 7317 14243
rect 7403 14187 7459 14243
rect 7545 14187 7601 14243
rect 7687 14187 7743 14243
rect 7829 14187 7885 14243
rect 7971 14187 8027 14243
rect 8113 14187 8169 14243
rect 8255 14187 8311 14243
rect 8397 14187 8453 14243
rect 8539 14187 8595 14243
rect 8681 14187 8737 14243
rect 8823 14187 8879 14243
rect 8965 14187 9021 14243
rect 9107 14187 9163 14243
rect 9249 14187 9305 14243
rect 9391 14187 9447 14243
rect 9533 14187 9589 14243
rect 9675 14187 9731 14243
rect 9817 14187 9873 14243
rect 9959 14187 10015 14243
rect 10101 14187 10157 14243
rect 10243 14187 10299 14243
rect 10385 14187 10441 14243
rect 10527 14187 10583 14243
rect 10669 14187 10725 14243
rect 10811 14187 10867 14243
rect 10953 14187 11009 14243
rect 11095 14187 11151 14243
rect 11237 14187 11293 14243
rect 11379 14187 11435 14243
rect 11521 14187 11577 14243
rect 11663 14187 11719 14243
rect 11805 14187 11861 14243
rect 11947 14187 12003 14243
rect 12089 14187 12145 14243
rect 12231 14187 12287 14243
rect 12373 14187 12429 14243
rect 12515 14187 12571 14243
rect 12657 14187 12713 14243
rect 12799 14187 12855 14243
rect 12941 14187 12997 14243
rect 13083 14187 13139 14243
rect 13225 14187 13281 14243
rect 13367 14187 13423 14243
rect 13509 14187 13565 14243
rect 13651 14187 13707 14243
rect 13793 14187 13849 14243
rect 13935 14187 13991 14243
rect 14077 14187 14133 14243
rect 14219 14187 14275 14243
rect 14361 14187 14417 14243
rect 14503 14187 14559 14243
rect 14645 14187 14701 14243
rect 14787 14187 14843 14243
rect 161 14045 217 14101
rect 303 14045 359 14101
rect 445 14045 501 14101
rect 587 14045 643 14101
rect 729 14045 785 14101
rect 871 14045 927 14101
rect 1013 14045 1069 14101
rect 1155 14045 1211 14101
rect 1297 14045 1353 14101
rect 1439 14045 1495 14101
rect 1581 14045 1637 14101
rect 1723 14045 1779 14101
rect 1865 14045 1921 14101
rect 2007 14045 2063 14101
rect 2149 14045 2205 14101
rect 2291 14045 2347 14101
rect 2433 14045 2489 14101
rect 2575 14045 2631 14101
rect 2717 14045 2773 14101
rect 2859 14045 2915 14101
rect 3001 14045 3057 14101
rect 3143 14045 3199 14101
rect 3285 14045 3341 14101
rect 3427 14045 3483 14101
rect 3569 14045 3625 14101
rect 3711 14045 3767 14101
rect 3853 14045 3909 14101
rect 3995 14045 4051 14101
rect 4137 14045 4193 14101
rect 4279 14045 4335 14101
rect 4421 14045 4477 14101
rect 4563 14045 4619 14101
rect 4705 14045 4761 14101
rect 4847 14045 4903 14101
rect 4989 14045 5045 14101
rect 5131 14045 5187 14101
rect 5273 14045 5329 14101
rect 5415 14045 5471 14101
rect 5557 14045 5613 14101
rect 5699 14045 5755 14101
rect 5841 14045 5897 14101
rect 5983 14045 6039 14101
rect 6125 14045 6181 14101
rect 6267 14045 6323 14101
rect 6409 14045 6465 14101
rect 6551 14045 6607 14101
rect 6693 14045 6749 14101
rect 6835 14045 6891 14101
rect 6977 14045 7033 14101
rect 7119 14045 7175 14101
rect 7261 14045 7317 14101
rect 7403 14045 7459 14101
rect 7545 14045 7601 14101
rect 7687 14045 7743 14101
rect 7829 14045 7885 14101
rect 7971 14045 8027 14101
rect 8113 14045 8169 14101
rect 8255 14045 8311 14101
rect 8397 14045 8453 14101
rect 8539 14045 8595 14101
rect 8681 14045 8737 14101
rect 8823 14045 8879 14101
rect 8965 14045 9021 14101
rect 9107 14045 9163 14101
rect 9249 14045 9305 14101
rect 9391 14045 9447 14101
rect 9533 14045 9589 14101
rect 9675 14045 9731 14101
rect 9817 14045 9873 14101
rect 9959 14045 10015 14101
rect 10101 14045 10157 14101
rect 10243 14045 10299 14101
rect 10385 14045 10441 14101
rect 10527 14045 10583 14101
rect 10669 14045 10725 14101
rect 10811 14045 10867 14101
rect 10953 14045 11009 14101
rect 11095 14045 11151 14101
rect 11237 14045 11293 14101
rect 11379 14045 11435 14101
rect 11521 14045 11577 14101
rect 11663 14045 11719 14101
rect 11805 14045 11861 14101
rect 11947 14045 12003 14101
rect 12089 14045 12145 14101
rect 12231 14045 12287 14101
rect 12373 14045 12429 14101
rect 12515 14045 12571 14101
rect 12657 14045 12713 14101
rect 12799 14045 12855 14101
rect 12941 14045 12997 14101
rect 13083 14045 13139 14101
rect 13225 14045 13281 14101
rect 13367 14045 13423 14101
rect 13509 14045 13565 14101
rect 13651 14045 13707 14101
rect 13793 14045 13849 14101
rect 13935 14045 13991 14101
rect 14077 14045 14133 14101
rect 14219 14045 14275 14101
rect 14361 14045 14417 14101
rect 14503 14045 14559 14101
rect 14645 14045 14701 14101
rect 14787 14045 14843 14101
<< metal4 >>
rect 0 69637 15000 69678
rect 0 69581 161 69637
rect 217 69581 303 69637
rect 359 69581 445 69637
rect 501 69581 587 69637
rect 643 69581 729 69637
rect 785 69581 871 69637
rect 927 69581 1013 69637
rect 1069 69581 1155 69637
rect 1211 69581 1297 69637
rect 1353 69581 1439 69637
rect 1495 69581 1581 69637
rect 1637 69581 1723 69637
rect 1779 69581 1865 69637
rect 1921 69581 2007 69637
rect 2063 69581 2149 69637
rect 2205 69581 2291 69637
rect 2347 69581 2433 69637
rect 2489 69581 2575 69637
rect 2631 69581 2717 69637
rect 2773 69581 2859 69637
rect 2915 69581 3001 69637
rect 3057 69581 3143 69637
rect 3199 69581 3285 69637
rect 3341 69581 3427 69637
rect 3483 69581 3569 69637
rect 3625 69581 3711 69637
rect 3767 69581 3853 69637
rect 3909 69581 3995 69637
rect 4051 69581 4137 69637
rect 4193 69581 4279 69637
rect 4335 69581 4421 69637
rect 4477 69581 4563 69637
rect 4619 69581 4705 69637
rect 4761 69581 4847 69637
rect 4903 69581 4989 69637
rect 5045 69581 5131 69637
rect 5187 69581 5273 69637
rect 5329 69581 5415 69637
rect 5471 69581 5557 69637
rect 5613 69581 5699 69637
rect 5755 69581 5841 69637
rect 5897 69581 5983 69637
rect 6039 69581 6125 69637
rect 6181 69581 6267 69637
rect 6323 69581 6409 69637
rect 6465 69581 6551 69637
rect 6607 69581 6693 69637
rect 6749 69581 6835 69637
rect 6891 69581 6977 69637
rect 7033 69581 7119 69637
rect 7175 69581 7261 69637
rect 7317 69581 7403 69637
rect 7459 69581 7545 69637
rect 7601 69581 7687 69637
rect 7743 69581 7829 69637
rect 7885 69581 7971 69637
rect 8027 69581 8113 69637
rect 8169 69581 8255 69637
rect 8311 69581 8397 69637
rect 8453 69581 8539 69637
rect 8595 69581 8681 69637
rect 8737 69581 8823 69637
rect 8879 69581 8965 69637
rect 9021 69581 9107 69637
rect 9163 69581 9249 69637
rect 9305 69581 9391 69637
rect 9447 69581 9533 69637
rect 9589 69581 9675 69637
rect 9731 69581 9817 69637
rect 9873 69581 9959 69637
rect 10015 69581 10101 69637
rect 10157 69581 10243 69637
rect 10299 69581 10385 69637
rect 10441 69581 10527 69637
rect 10583 69581 10669 69637
rect 10725 69581 10811 69637
rect 10867 69581 10953 69637
rect 11009 69581 11095 69637
rect 11151 69581 11237 69637
rect 11293 69581 11379 69637
rect 11435 69581 11521 69637
rect 11577 69581 11663 69637
rect 11719 69581 11805 69637
rect 11861 69581 11947 69637
rect 12003 69581 12089 69637
rect 12145 69581 12231 69637
rect 12287 69581 12373 69637
rect 12429 69581 12515 69637
rect 12571 69581 12657 69637
rect 12713 69581 12799 69637
rect 12855 69581 12941 69637
rect 12997 69581 13083 69637
rect 13139 69581 13225 69637
rect 13281 69581 13367 69637
rect 13423 69581 13509 69637
rect 13565 69581 13651 69637
rect 13707 69581 13793 69637
rect 13849 69581 13935 69637
rect 13991 69581 14077 69637
rect 14133 69581 14219 69637
rect 14275 69581 14361 69637
rect 14417 69581 14503 69637
rect 14559 69581 14645 69637
rect 14701 69581 14787 69637
rect 14843 69581 15000 69637
rect 0 69495 15000 69581
rect 0 69439 161 69495
rect 217 69439 303 69495
rect 359 69439 445 69495
rect 501 69439 587 69495
rect 643 69439 729 69495
rect 785 69439 871 69495
rect 927 69439 1013 69495
rect 1069 69439 1155 69495
rect 1211 69439 1297 69495
rect 1353 69439 1439 69495
rect 1495 69439 1581 69495
rect 1637 69439 1723 69495
rect 1779 69439 1865 69495
rect 1921 69439 2007 69495
rect 2063 69439 2149 69495
rect 2205 69439 2291 69495
rect 2347 69439 2433 69495
rect 2489 69439 2575 69495
rect 2631 69439 2717 69495
rect 2773 69439 2859 69495
rect 2915 69439 3001 69495
rect 3057 69439 3143 69495
rect 3199 69439 3285 69495
rect 3341 69439 3427 69495
rect 3483 69439 3569 69495
rect 3625 69439 3711 69495
rect 3767 69439 3853 69495
rect 3909 69439 3995 69495
rect 4051 69439 4137 69495
rect 4193 69439 4279 69495
rect 4335 69439 4421 69495
rect 4477 69439 4563 69495
rect 4619 69439 4705 69495
rect 4761 69439 4847 69495
rect 4903 69439 4989 69495
rect 5045 69439 5131 69495
rect 5187 69439 5273 69495
rect 5329 69439 5415 69495
rect 5471 69439 5557 69495
rect 5613 69439 5699 69495
rect 5755 69439 5841 69495
rect 5897 69439 5983 69495
rect 6039 69439 6125 69495
rect 6181 69439 6267 69495
rect 6323 69439 6409 69495
rect 6465 69439 6551 69495
rect 6607 69439 6693 69495
rect 6749 69439 6835 69495
rect 6891 69439 6977 69495
rect 7033 69439 7119 69495
rect 7175 69439 7261 69495
rect 7317 69439 7403 69495
rect 7459 69439 7545 69495
rect 7601 69439 7687 69495
rect 7743 69439 7829 69495
rect 7885 69439 7971 69495
rect 8027 69439 8113 69495
rect 8169 69439 8255 69495
rect 8311 69439 8397 69495
rect 8453 69439 8539 69495
rect 8595 69439 8681 69495
rect 8737 69439 8823 69495
rect 8879 69439 8965 69495
rect 9021 69439 9107 69495
rect 9163 69439 9249 69495
rect 9305 69439 9391 69495
rect 9447 69439 9533 69495
rect 9589 69439 9675 69495
rect 9731 69439 9817 69495
rect 9873 69439 9959 69495
rect 10015 69439 10101 69495
rect 10157 69439 10243 69495
rect 10299 69439 10385 69495
rect 10441 69439 10527 69495
rect 10583 69439 10669 69495
rect 10725 69439 10811 69495
rect 10867 69439 10953 69495
rect 11009 69439 11095 69495
rect 11151 69439 11237 69495
rect 11293 69439 11379 69495
rect 11435 69439 11521 69495
rect 11577 69439 11663 69495
rect 11719 69439 11805 69495
rect 11861 69439 11947 69495
rect 12003 69439 12089 69495
rect 12145 69439 12231 69495
rect 12287 69439 12373 69495
rect 12429 69439 12515 69495
rect 12571 69439 12657 69495
rect 12713 69439 12799 69495
rect 12855 69439 12941 69495
rect 12997 69439 13083 69495
rect 13139 69439 13225 69495
rect 13281 69439 13367 69495
rect 13423 69439 13509 69495
rect 13565 69439 13651 69495
rect 13707 69439 13793 69495
rect 13849 69439 13935 69495
rect 13991 69439 14077 69495
rect 14133 69439 14219 69495
rect 14275 69439 14361 69495
rect 14417 69439 14503 69495
rect 14559 69439 14645 69495
rect 14701 69439 14787 69495
rect 14843 69439 15000 69495
rect 0 69353 15000 69439
rect 0 69297 161 69353
rect 217 69297 303 69353
rect 359 69297 445 69353
rect 501 69297 587 69353
rect 643 69297 729 69353
rect 785 69297 871 69353
rect 927 69297 1013 69353
rect 1069 69297 1155 69353
rect 1211 69297 1297 69353
rect 1353 69297 1439 69353
rect 1495 69297 1581 69353
rect 1637 69297 1723 69353
rect 1779 69297 1865 69353
rect 1921 69297 2007 69353
rect 2063 69297 2149 69353
rect 2205 69297 2291 69353
rect 2347 69297 2433 69353
rect 2489 69297 2575 69353
rect 2631 69297 2717 69353
rect 2773 69297 2859 69353
rect 2915 69297 3001 69353
rect 3057 69297 3143 69353
rect 3199 69297 3285 69353
rect 3341 69297 3427 69353
rect 3483 69297 3569 69353
rect 3625 69297 3711 69353
rect 3767 69297 3853 69353
rect 3909 69297 3995 69353
rect 4051 69297 4137 69353
rect 4193 69297 4279 69353
rect 4335 69297 4421 69353
rect 4477 69297 4563 69353
rect 4619 69297 4705 69353
rect 4761 69297 4847 69353
rect 4903 69297 4989 69353
rect 5045 69297 5131 69353
rect 5187 69297 5273 69353
rect 5329 69297 5415 69353
rect 5471 69297 5557 69353
rect 5613 69297 5699 69353
rect 5755 69297 5841 69353
rect 5897 69297 5983 69353
rect 6039 69297 6125 69353
rect 6181 69297 6267 69353
rect 6323 69297 6409 69353
rect 6465 69297 6551 69353
rect 6607 69297 6693 69353
rect 6749 69297 6835 69353
rect 6891 69297 6977 69353
rect 7033 69297 7119 69353
rect 7175 69297 7261 69353
rect 7317 69297 7403 69353
rect 7459 69297 7545 69353
rect 7601 69297 7687 69353
rect 7743 69297 7829 69353
rect 7885 69297 7971 69353
rect 8027 69297 8113 69353
rect 8169 69297 8255 69353
rect 8311 69297 8397 69353
rect 8453 69297 8539 69353
rect 8595 69297 8681 69353
rect 8737 69297 8823 69353
rect 8879 69297 8965 69353
rect 9021 69297 9107 69353
rect 9163 69297 9249 69353
rect 9305 69297 9391 69353
rect 9447 69297 9533 69353
rect 9589 69297 9675 69353
rect 9731 69297 9817 69353
rect 9873 69297 9959 69353
rect 10015 69297 10101 69353
rect 10157 69297 10243 69353
rect 10299 69297 10385 69353
rect 10441 69297 10527 69353
rect 10583 69297 10669 69353
rect 10725 69297 10811 69353
rect 10867 69297 10953 69353
rect 11009 69297 11095 69353
rect 11151 69297 11237 69353
rect 11293 69297 11379 69353
rect 11435 69297 11521 69353
rect 11577 69297 11663 69353
rect 11719 69297 11805 69353
rect 11861 69297 11947 69353
rect 12003 69297 12089 69353
rect 12145 69297 12231 69353
rect 12287 69297 12373 69353
rect 12429 69297 12515 69353
rect 12571 69297 12657 69353
rect 12713 69297 12799 69353
rect 12855 69297 12941 69353
rect 12997 69297 13083 69353
rect 13139 69297 13225 69353
rect 13281 69297 13367 69353
rect 13423 69297 13509 69353
rect 13565 69297 13651 69353
rect 13707 69297 13793 69353
rect 13849 69297 13935 69353
rect 13991 69297 14077 69353
rect 14133 69297 14219 69353
rect 14275 69297 14361 69353
rect 14417 69297 14503 69353
rect 14559 69297 14645 69353
rect 14701 69297 14787 69353
rect 14843 69297 15000 69353
rect 0 69211 15000 69297
rect 0 69155 161 69211
rect 217 69155 303 69211
rect 359 69155 445 69211
rect 501 69155 587 69211
rect 643 69155 729 69211
rect 785 69155 871 69211
rect 927 69155 1013 69211
rect 1069 69155 1155 69211
rect 1211 69155 1297 69211
rect 1353 69155 1439 69211
rect 1495 69155 1581 69211
rect 1637 69155 1723 69211
rect 1779 69155 1865 69211
rect 1921 69155 2007 69211
rect 2063 69155 2149 69211
rect 2205 69155 2291 69211
rect 2347 69155 2433 69211
rect 2489 69155 2575 69211
rect 2631 69155 2717 69211
rect 2773 69155 2859 69211
rect 2915 69155 3001 69211
rect 3057 69155 3143 69211
rect 3199 69155 3285 69211
rect 3341 69155 3427 69211
rect 3483 69155 3569 69211
rect 3625 69155 3711 69211
rect 3767 69155 3853 69211
rect 3909 69155 3995 69211
rect 4051 69155 4137 69211
rect 4193 69155 4279 69211
rect 4335 69155 4421 69211
rect 4477 69155 4563 69211
rect 4619 69155 4705 69211
rect 4761 69155 4847 69211
rect 4903 69155 4989 69211
rect 5045 69155 5131 69211
rect 5187 69155 5273 69211
rect 5329 69155 5415 69211
rect 5471 69155 5557 69211
rect 5613 69155 5699 69211
rect 5755 69155 5841 69211
rect 5897 69155 5983 69211
rect 6039 69155 6125 69211
rect 6181 69155 6267 69211
rect 6323 69155 6409 69211
rect 6465 69155 6551 69211
rect 6607 69155 6693 69211
rect 6749 69155 6835 69211
rect 6891 69155 6977 69211
rect 7033 69155 7119 69211
rect 7175 69155 7261 69211
rect 7317 69155 7403 69211
rect 7459 69155 7545 69211
rect 7601 69155 7687 69211
rect 7743 69155 7829 69211
rect 7885 69155 7971 69211
rect 8027 69155 8113 69211
rect 8169 69155 8255 69211
rect 8311 69155 8397 69211
rect 8453 69155 8539 69211
rect 8595 69155 8681 69211
rect 8737 69155 8823 69211
rect 8879 69155 8965 69211
rect 9021 69155 9107 69211
rect 9163 69155 9249 69211
rect 9305 69155 9391 69211
rect 9447 69155 9533 69211
rect 9589 69155 9675 69211
rect 9731 69155 9817 69211
rect 9873 69155 9959 69211
rect 10015 69155 10101 69211
rect 10157 69155 10243 69211
rect 10299 69155 10385 69211
rect 10441 69155 10527 69211
rect 10583 69155 10669 69211
rect 10725 69155 10811 69211
rect 10867 69155 10953 69211
rect 11009 69155 11095 69211
rect 11151 69155 11237 69211
rect 11293 69155 11379 69211
rect 11435 69155 11521 69211
rect 11577 69155 11663 69211
rect 11719 69155 11805 69211
rect 11861 69155 11947 69211
rect 12003 69155 12089 69211
rect 12145 69155 12231 69211
rect 12287 69155 12373 69211
rect 12429 69155 12515 69211
rect 12571 69155 12657 69211
rect 12713 69155 12799 69211
rect 12855 69155 12941 69211
rect 12997 69155 13083 69211
rect 13139 69155 13225 69211
rect 13281 69155 13367 69211
rect 13423 69155 13509 69211
rect 13565 69155 13651 69211
rect 13707 69155 13793 69211
rect 13849 69155 13935 69211
rect 13991 69155 14077 69211
rect 14133 69155 14219 69211
rect 14275 69155 14361 69211
rect 14417 69155 14503 69211
rect 14559 69155 14645 69211
rect 14701 69155 14787 69211
rect 14843 69155 15000 69211
rect 0 69069 15000 69155
rect 0 69013 161 69069
rect 217 69013 303 69069
rect 359 69013 445 69069
rect 501 69013 587 69069
rect 643 69013 729 69069
rect 785 69013 871 69069
rect 927 69013 1013 69069
rect 1069 69013 1155 69069
rect 1211 69013 1297 69069
rect 1353 69013 1439 69069
rect 1495 69013 1581 69069
rect 1637 69013 1723 69069
rect 1779 69013 1865 69069
rect 1921 69013 2007 69069
rect 2063 69013 2149 69069
rect 2205 69013 2291 69069
rect 2347 69013 2433 69069
rect 2489 69013 2575 69069
rect 2631 69013 2717 69069
rect 2773 69013 2859 69069
rect 2915 69013 3001 69069
rect 3057 69013 3143 69069
rect 3199 69013 3285 69069
rect 3341 69013 3427 69069
rect 3483 69013 3569 69069
rect 3625 69013 3711 69069
rect 3767 69013 3853 69069
rect 3909 69013 3995 69069
rect 4051 69013 4137 69069
rect 4193 69013 4279 69069
rect 4335 69013 4421 69069
rect 4477 69013 4563 69069
rect 4619 69013 4705 69069
rect 4761 69013 4847 69069
rect 4903 69013 4989 69069
rect 5045 69013 5131 69069
rect 5187 69013 5273 69069
rect 5329 69013 5415 69069
rect 5471 69013 5557 69069
rect 5613 69013 5699 69069
rect 5755 69013 5841 69069
rect 5897 69013 5983 69069
rect 6039 69013 6125 69069
rect 6181 69013 6267 69069
rect 6323 69013 6409 69069
rect 6465 69013 6551 69069
rect 6607 69013 6693 69069
rect 6749 69013 6835 69069
rect 6891 69013 6977 69069
rect 7033 69013 7119 69069
rect 7175 69013 7261 69069
rect 7317 69013 7403 69069
rect 7459 69013 7545 69069
rect 7601 69013 7687 69069
rect 7743 69013 7829 69069
rect 7885 69013 7971 69069
rect 8027 69013 8113 69069
rect 8169 69013 8255 69069
rect 8311 69013 8397 69069
rect 8453 69013 8539 69069
rect 8595 69013 8681 69069
rect 8737 69013 8823 69069
rect 8879 69013 8965 69069
rect 9021 69013 9107 69069
rect 9163 69013 9249 69069
rect 9305 69013 9391 69069
rect 9447 69013 9533 69069
rect 9589 69013 9675 69069
rect 9731 69013 9817 69069
rect 9873 69013 9959 69069
rect 10015 69013 10101 69069
rect 10157 69013 10243 69069
rect 10299 69013 10385 69069
rect 10441 69013 10527 69069
rect 10583 69013 10669 69069
rect 10725 69013 10811 69069
rect 10867 69013 10953 69069
rect 11009 69013 11095 69069
rect 11151 69013 11237 69069
rect 11293 69013 11379 69069
rect 11435 69013 11521 69069
rect 11577 69013 11663 69069
rect 11719 69013 11805 69069
rect 11861 69013 11947 69069
rect 12003 69013 12089 69069
rect 12145 69013 12231 69069
rect 12287 69013 12373 69069
rect 12429 69013 12515 69069
rect 12571 69013 12657 69069
rect 12713 69013 12799 69069
rect 12855 69013 12941 69069
rect 12997 69013 13083 69069
rect 13139 69013 13225 69069
rect 13281 69013 13367 69069
rect 13423 69013 13509 69069
rect 13565 69013 13651 69069
rect 13707 69013 13793 69069
rect 13849 69013 13935 69069
rect 13991 69013 14077 69069
rect 14133 69013 14219 69069
rect 14275 69013 14361 69069
rect 14417 69013 14503 69069
rect 14559 69013 14645 69069
rect 14701 69013 14787 69069
rect 14843 69013 15000 69069
rect 0 68927 15000 69013
rect 0 68871 161 68927
rect 217 68871 303 68927
rect 359 68871 445 68927
rect 501 68871 587 68927
rect 643 68871 729 68927
rect 785 68871 871 68927
rect 927 68871 1013 68927
rect 1069 68871 1155 68927
rect 1211 68871 1297 68927
rect 1353 68871 1439 68927
rect 1495 68871 1581 68927
rect 1637 68871 1723 68927
rect 1779 68871 1865 68927
rect 1921 68871 2007 68927
rect 2063 68871 2149 68927
rect 2205 68871 2291 68927
rect 2347 68871 2433 68927
rect 2489 68871 2575 68927
rect 2631 68871 2717 68927
rect 2773 68871 2859 68927
rect 2915 68871 3001 68927
rect 3057 68871 3143 68927
rect 3199 68871 3285 68927
rect 3341 68871 3427 68927
rect 3483 68871 3569 68927
rect 3625 68871 3711 68927
rect 3767 68871 3853 68927
rect 3909 68871 3995 68927
rect 4051 68871 4137 68927
rect 4193 68871 4279 68927
rect 4335 68871 4421 68927
rect 4477 68871 4563 68927
rect 4619 68871 4705 68927
rect 4761 68871 4847 68927
rect 4903 68871 4989 68927
rect 5045 68871 5131 68927
rect 5187 68871 5273 68927
rect 5329 68871 5415 68927
rect 5471 68871 5557 68927
rect 5613 68871 5699 68927
rect 5755 68871 5841 68927
rect 5897 68871 5983 68927
rect 6039 68871 6125 68927
rect 6181 68871 6267 68927
rect 6323 68871 6409 68927
rect 6465 68871 6551 68927
rect 6607 68871 6693 68927
rect 6749 68871 6835 68927
rect 6891 68871 6977 68927
rect 7033 68871 7119 68927
rect 7175 68871 7261 68927
rect 7317 68871 7403 68927
rect 7459 68871 7545 68927
rect 7601 68871 7687 68927
rect 7743 68871 7829 68927
rect 7885 68871 7971 68927
rect 8027 68871 8113 68927
rect 8169 68871 8255 68927
rect 8311 68871 8397 68927
rect 8453 68871 8539 68927
rect 8595 68871 8681 68927
rect 8737 68871 8823 68927
rect 8879 68871 8965 68927
rect 9021 68871 9107 68927
rect 9163 68871 9249 68927
rect 9305 68871 9391 68927
rect 9447 68871 9533 68927
rect 9589 68871 9675 68927
rect 9731 68871 9817 68927
rect 9873 68871 9959 68927
rect 10015 68871 10101 68927
rect 10157 68871 10243 68927
rect 10299 68871 10385 68927
rect 10441 68871 10527 68927
rect 10583 68871 10669 68927
rect 10725 68871 10811 68927
rect 10867 68871 10953 68927
rect 11009 68871 11095 68927
rect 11151 68871 11237 68927
rect 11293 68871 11379 68927
rect 11435 68871 11521 68927
rect 11577 68871 11663 68927
rect 11719 68871 11805 68927
rect 11861 68871 11947 68927
rect 12003 68871 12089 68927
rect 12145 68871 12231 68927
rect 12287 68871 12373 68927
rect 12429 68871 12515 68927
rect 12571 68871 12657 68927
rect 12713 68871 12799 68927
rect 12855 68871 12941 68927
rect 12997 68871 13083 68927
rect 13139 68871 13225 68927
rect 13281 68871 13367 68927
rect 13423 68871 13509 68927
rect 13565 68871 13651 68927
rect 13707 68871 13793 68927
rect 13849 68871 13935 68927
rect 13991 68871 14077 68927
rect 14133 68871 14219 68927
rect 14275 68871 14361 68927
rect 14417 68871 14503 68927
rect 14559 68871 14645 68927
rect 14701 68871 14787 68927
rect 14843 68871 15000 68927
rect 0 68785 15000 68871
rect 0 68729 161 68785
rect 217 68729 303 68785
rect 359 68729 445 68785
rect 501 68729 587 68785
rect 643 68729 729 68785
rect 785 68729 871 68785
rect 927 68729 1013 68785
rect 1069 68729 1155 68785
rect 1211 68729 1297 68785
rect 1353 68729 1439 68785
rect 1495 68729 1581 68785
rect 1637 68729 1723 68785
rect 1779 68729 1865 68785
rect 1921 68729 2007 68785
rect 2063 68729 2149 68785
rect 2205 68729 2291 68785
rect 2347 68729 2433 68785
rect 2489 68729 2575 68785
rect 2631 68729 2717 68785
rect 2773 68729 2859 68785
rect 2915 68729 3001 68785
rect 3057 68729 3143 68785
rect 3199 68729 3285 68785
rect 3341 68729 3427 68785
rect 3483 68729 3569 68785
rect 3625 68729 3711 68785
rect 3767 68729 3853 68785
rect 3909 68729 3995 68785
rect 4051 68729 4137 68785
rect 4193 68729 4279 68785
rect 4335 68729 4421 68785
rect 4477 68729 4563 68785
rect 4619 68729 4705 68785
rect 4761 68729 4847 68785
rect 4903 68729 4989 68785
rect 5045 68729 5131 68785
rect 5187 68729 5273 68785
rect 5329 68729 5415 68785
rect 5471 68729 5557 68785
rect 5613 68729 5699 68785
rect 5755 68729 5841 68785
rect 5897 68729 5983 68785
rect 6039 68729 6125 68785
rect 6181 68729 6267 68785
rect 6323 68729 6409 68785
rect 6465 68729 6551 68785
rect 6607 68729 6693 68785
rect 6749 68729 6835 68785
rect 6891 68729 6977 68785
rect 7033 68729 7119 68785
rect 7175 68729 7261 68785
rect 7317 68729 7403 68785
rect 7459 68729 7545 68785
rect 7601 68729 7687 68785
rect 7743 68729 7829 68785
rect 7885 68729 7971 68785
rect 8027 68729 8113 68785
rect 8169 68729 8255 68785
rect 8311 68729 8397 68785
rect 8453 68729 8539 68785
rect 8595 68729 8681 68785
rect 8737 68729 8823 68785
rect 8879 68729 8965 68785
rect 9021 68729 9107 68785
rect 9163 68729 9249 68785
rect 9305 68729 9391 68785
rect 9447 68729 9533 68785
rect 9589 68729 9675 68785
rect 9731 68729 9817 68785
rect 9873 68729 9959 68785
rect 10015 68729 10101 68785
rect 10157 68729 10243 68785
rect 10299 68729 10385 68785
rect 10441 68729 10527 68785
rect 10583 68729 10669 68785
rect 10725 68729 10811 68785
rect 10867 68729 10953 68785
rect 11009 68729 11095 68785
rect 11151 68729 11237 68785
rect 11293 68729 11379 68785
rect 11435 68729 11521 68785
rect 11577 68729 11663 68785
rect 11719 68729 11805 68785
rect 11861 68729 11947 68785
rect 12003 68729 12089 68785
rect 12145 68729 12231 68785
rect 12287 68729 12373 68785
rect 12429 68729 12515 68785
rect 12571 68729 12657 68785
rect 12713 68729 12799 68785
rect 12855 68729 12941 68785
rect 12997 68729 13083 68785
rect 13139 68729 13225 68785
rect 13281 68729 13367 68785
rect 13423 68729 13509 68785
rect 13565 68729 13651 68785
rect 13707 68729 13793 68785
rect 13849 68729 13935 68785
rect 13991 68729 14077 68785
rect 14133 68729 14219 68785
rect 14275 68729 14361 68785
rect 14417 68729 14503 68785
rect 14559 68729 14645 68785
rect 14701 68729 14787 68785
rect 14843 68729 15000 68785
rect 0 68643 15000 68729
rect 0 68587 161 68643
rect 217 68587 303 68643
rect 359 68587 445 68643
rect 501 68587 587 68643
rect 643 68587 729 68643
rect 785 68587 871 68643
rect 927 68587 1013 68643
rect 1069 68587 1155 68643
rect 1211 68587 1297 68643
rect 1353 68587 1439 68643
rect 1495 68587 1581 68643
rect 1637 68587 1723 68643
rect 1779 68587 1865 68643
rect 1921 68587 2007 68643
rect 2063 68587 2149 68643
rect 2205 68587 2291 68643
rect 2347 68587 2433 68643
rect 2489 68587 2575 68643
rect 2631 68587 2717 68643
rect 2773 68587 2859 68643
rect 2915 68587 3001 68643
rect 3057 68587 3143 68643
rect 3199 68587 3285 68643
rect 3341 68587 3427 68643
rect 3483 68587 3569 68643
rect 3625 68587 3711 68643
rect 3767 68587 3853 68643
rect 3909 68587 3995 68643
rect 4051 68587 4137 68643
rect 4193 68587 4279 68643
rect 4335 68587 4421 68643
rect 4477 68587 4563 68643
rect 4619 68587 4705 68643
rect 4761 68587 4847 68643
rect 4903 68587 4989 68643
rect 5045 68587 5131 68643
rect 5187 68587 5273 68643
rect 5329 68587 5415 68643
rect 5471 68587 5557 68643
rect 5613 68587 5699 68643
rect 5755 68587 5841 68643
rect 5897 68587 5983 68643
rect 6039 68587 6125 68643
rect 6181 68587 6267 68643
rect 6323 68587 6409 68643
rect 6465 68587 6551 68643
rect 6607 68587 6693 68643
rect 6749 68587 6835 68643
rect 6891 68587 6977 68643
rect 7033 68587 7119 68643
rect 7175 68587 7261 68643
rect 7317 68587 7403 68643
rect 7459 68587 7545 68643
rect 7601 68587 7687 68643
rect 7743 68587 7829 68643
rect 7885 68587 7971 68643
rect 8027 68587 8113 68643
rect 8169 68587 8255 68643
rect 8311 68587 8397 68643
rect 8453 68587 8539 68643
rect 8595 68587 8681 68643
rect 8737 68587 8823 68643
rect 8879 68587 8965 68643
rect 9021 68587 9107 68643
rect 9163 68587 9249 68643
rect 9305 68587 9391 68643
rect 9447 68587 9533 68643
rect 9589 68587 9675 68643
rect 9731 68587 9817 68643
rect 9873 68587 9959 68643
rect 10015 68587 10101 68643
rect 10157 68587 10243 68643
rect 10299 68587 10385 68643
rect 10441 68587 10527 68643
rect 10583 68587 10669 68643
rect 10725 68587 10811 68643
rect 10867 68587 10953 68643
rect 11009 68587 11095 68643
rect 11151 68587 11237 68643
rect 11293 68587 11379 68643
rect 11435 68587 11521 68643
rect 11577 68587 11663 68643
rect 11719 68587 11805 68643
rect 11861 68587 11947 68643
rect 12003 68587 12089 68643
rect 12145 68587 12231 68643
rect 12287 68587 12373 68643
rect 12429 68587 12515 68643
rect 12571 68587 12657 68643
rect 12713 68587 12799 68643
rect 12855 68587 12941 68643
rect 12997 68587 13083 68643
rect 13139 68587 13225 68643
rect 13281 68587 13367 68643
rect 13423 68587 13509 68643
rect 13565 68587 13651 68643
rect 13707 68587 13793 68643
rect 13849 68587 13935 68643
rect 13991 68587 14077 68643
rect 14133 68587 14219 68643
rect 14275 68587 14361 68643
rect 14417 68587 14503 68643
rect 14559 68587 14645 68643
rect 14701 68587 14787 68643
rect 14843 68587 15000 68643
rect 0 68501 15000 68587
rect 0 68445 161 68501
rect 217 68445 303 68501
rect 359 68445 445 68501
rect 501 68445 587 68501
rect 643 68445 729 68501
rect 785 68445 871 68501
rect 927 68445 1013 68501
rect 1069 68445 1155 68501
rect 1211 68445 1297 68501
rect 1353 68445 1439 68501
rect 1495 68445 1581 68501
rect 1637 68445 1723 68501
rect 1779 68445 1865 68501
rect 1921 68445 2007 68501
rect 2063 68445 2149 68501
rect 2205 68445 2291 68501
rect 2347 68445 2433 68501
rect 2489 68445 2575 68501
rect 2631 68445 2717 68501
rect 2773 68445 2859 68501
rect 2915 68445 3001 68501
rect 3057 68445 3143 68501
rect 3199 68445 3285 68501
rect 3341 68445 3427 68501
rect 3483 68445 3569 68501
rect 3625 68445 3711 68501
rect 3767 68445 3853 68501
rect 3909 68445 3995 68501
rect 4051 68445 4137 68501
rect 4193 68445 4279 68501
rect 4335 68445 4421 68501
rect 4477 68445 4563 68501
rect 4619 68445 4705 68501
rect 4761 68445 4847 68501
rect 4903 68445 4989 68501
rect 5045 68445 5131 68501
rect 5187 68445 5273 68501
rect 5329 68445 5415 68501
rect 5471 68445 5557 68501
rect 5613 68445 5699 68501
rect 5755 68445 5841 68501
rect 5897 68445 5983 68501
rect 6039 68445 6125 68501
rect 6181 68445 6267 68501
rect 6323 68445 6409 68501
rect 6465 68445 6551 68501
rect 6607 68445 6693 68501
rect 6749 68445 6835 68501
rect 6891 68445 6977 68501
rect 7033 68445 7119 68501
rect 7175 68445 7261 68501
rect 7317 68445 7403 68501
rect 7459 68445 7545 68501
rect 7601 68445 7687 68501
rect 7743 68445 7829 68501
rect 7885 68445 7971 68501
rect 8027 68445 8113 68501
rect 8169 68445 8255 68501
rect 8311 68445 8397 68501
rect 8453 68445 8539 68501
rect 8595 68445 8681 68501
rect 8737 68445 8823 68501
rect 8879 68445 8965 68501
rect 9021 68445 9107 68501
rect 9163 68445 9249 68501
rect 9305 68445 9391 68501
rect 9447 68445 9533 68501
rect 9589 68445 9675 68501
rect 9731 68445 9817 68501
rect 9873 68445 9959 68501
rect 10015 68445 10101 68501
rect 10157 68445 10243 68501
rect 10299 68445 10385 68501
rect 10441 68445 10527 68501
rect 10583 68445 10669 68501
rect 10725 68445 10811 68501
rect 10867 68445 10953 68501
rect 11009 68445 11095 68501
rect 11151 68445 11237 68501
rect 11293 68445 11379 68501
rect 11435 68445 11521 68501
rect 11577 68445 11663 68501
rect 11719 68445 11805 68501
rect 11861 68445 11947 68501
rect 12003 68445 12089 68501
rect 12145 68445 12231 68501
rect 12287 68445 12373 68501
rect 12429 68445 12515 68501
rect 12571 68445 12657 68501
rect 12713 68445 12799 68501
rect 12855 68445 12941 68501
rect 12997 68445 13083 68501
rect 13139 68445 13225 68501
rect 13281 68445 13367 68501
rect 13423 68445 13509 68501
rect 13565 68445 13651 68501
rect 13707 68445 13793 68501
rect 13849 68445 13935 68501
rect 13991 68445 14077 68501
rect 14133 68445 14219 68501
rect 14275 68445 14361 68501
rect 14417 68445 14503 68501
rect 14559 68445 14645 68501
rect 14701 68445 14787 68501
rect 14843 68445 15000 68501
rect 0 68400 15000 68445
rect 0 68171 15000 68200
rect 0 68115 161 68171
rect 217 68115 303 68171
rect 359 68115 445 68171
rect 501 68115 587 68171
rect 643 68115 729 68171
rect 785 68115 871 68171
rect 927 68115 1013 68171
rect 1069 68115 1155 68171
rect 1211 68115 1297 68171
rect 1353 68115 1439 68171
rect 1495 68115 1581 68171
rect 1637 68115 1723 68171
rect 1779 68115 1865 68171
rect 1921 68115 2007 68171
rect 2063 68115 2149 68171
rect 2205 68115 2291 68171
rect 2347 68115 2433 68171
rect 2489 68115 2575 68171
rect 2631 68115 2717 68171
rect 2773 68115 2859 68171
rect 2915 68115 3001 68171
rect 3057 68115 3143 68171
rect 3199 68115 3285 68171
rect 3341 68115 3427 68171
rect 3483 68115 3569 68171
rect 3625 68115 3711 68171
rect 3767 68115 3853 68171
rect 3909 68115 3995 68171
rect 4051 68115 4137 68171
rect 4193 68115 4279 68171
rect 4335 68115 4421 68171
rect 4477 68115 4563 68171
rect 4619 68115 4705 68171
rect 4761 68115 4847 68171
rect 4903 68115 4989 68171
rect 5045 68115 5131 68171
rect 5187 68115 5273 68171
rect 5329 68115 5415 68171
rect 5471 68115 5557 68171
rect 5613 68115 5699 68171
rect 5755 68115 5841 68171
rect 5897 68115 5983 68171
rect 6039 68115 6125 68171
rect 6181 68115 6267 68171
rect 6323 68115 6409 68171
rect 6465 68115 6551 68171
rect 6607 68115 6693 68171
rect 6749 68115 6835 68171
rect 6891 68115 6977 68171
rect 7033 68115 7119 68171
rect 7175 68115 7261 68171
rect 7317 68115 7403 68171
rect 7459 68115 7545 68171
rect 7601 68115 7687 68171
rect 7743 68115 7829 68171
rect 7885 68115 7971 68171
rect 8027 68115 8113 68171
rect 8169 68115 8255 68171
rect 8311 68115 8397 68171
rect 8453 68115 8539 68171
rect 8595 68115 8681 68171
rect 8737 68115 8823 68171
rect 8879 68115 8965 68171
rect 9021 68115 9107 68171
rect 9163 68115 9249 68171
rect 9305 68115 9391 68171
rect 9447 68115 9533 68171
rect 9589 68115 9675 68171
rect 9731 68115 9817 68171
rect 9873 68115 9959 68171
rect 10015 68115 10101 68171
rect 10157 68115 10243 68171
rect 10299 68115 10385 68171
rect 10441 68115 10527 68171
rect 10583 68115 10669 68171
rect 10725 68115 10811 68171
rect 10867 68115 10953 68171
rect 11009 68115 11095 68171
rect 11151 68115 11237 68171
rect 11293 68115 11379 68171
rect 11435 68115 11521 68171
rect 11577 68115 11663 68171
rect 11719 68115 11805 68171
rect 11861 68115 11947 68171
rect 12003 68115 12089 68171
rect 12145 68115 12231 68171
rect 12287 68115 12373 68171
rect 12429 68115 12515 68171
rect 12571 68115 12657 68171
rect 12713 68115 12799 68171
rect 12855 68115 12941 68171
rect 12997 68115 13083 68171
rect 13139 68115 13225 68171
rect 13281 68115 13367 68171
rect 13423 68115 13509 68171
rect 13565 68115 13651 68171
rect 13707 68115 13793 68171
rect 13849 68115 13935 68171
rect 13991 68115 14077 68171
rect 14133 68115 14219 68171
rect 14275 68115 14361 68171
rect 14417 68115 14503 68171
rect 14559 68115 14645 68171
rect 14701 68115 14787 68171
rect 14843 68115 15000 68171
rect 0 68029 15000 68115
rect 0 67973 161 68029
rect 217 67973 303 68029
rect 359 67973 445 68029
rect 501 67973 587 68029
rect 643 67973 729 68029
rect 785 67973 871 68029
rect 927 67973 1013 68029
rect 1069 67973 1155 68029
rect 1211 67973 1297 68029
rect 1353 67973 1439 68029
rect 1495 67973 1581 68029
rect 1637 67973 1723 68029
rect 1779 67973 1865 68029
rect 1921 67973 2007 68029
rect 2063 67973 2149 68029
rect 2205 67973 2291 68029
rect 2347 67973 2433 68029
rect 2489 67973 2575 68029
rect 2631 67973 2717 68029
rect 2773 67973 2859 68029
rect 2915 67973 3001 68029
rect 3057 67973 3143 68029
rect 3199 67973 3285 68029
rect 3341 67973 3427 68029
rect 3483 67973 3569 68029
rect 3625 67973 3711 68029
rect 3767 67973 3853 68029
rect 3909 67973 3995 68029
rect 4051 67973 4137 68029
rect 4193 67973 4279 68029
rect 4335 67973 4421 68029
rect 4477 67973 4563 68029
rect 4619 67973 4705 68029
rect 4761 67973 4847 68029
rect 4903 67973 4989 68029
rect 5045 67973 5131 68029
rect 5187 67973 5273 68029
rect 5329 67973 5415 68029
rect 5471 67973 5557 68029
rect 5613 67973 5699 68029
rect 5755 67973 5841 68029
rect 5897 67973 5983 68029
rect 6039 67973 6125 68029
rect 6181 67973 6267 68029
rect 6323 67973 6409 68029
rect 6465 67973 6551 68029
rect 6607 67973 6693 68029
rect 6749 67973 6835 68029
rect 6891 67973 6977 68029
rect 7033 67973 7119 68029
rect 7175 67973 7261 68029
rect 7317 67973 7403 68029
rect 7459 67973 7545 68029
rect 7601 67973 7687 68029
rect 7743 67973 7829 68029
rect 7885 67973 7971 68029
rect 8027 67973 8113 68029
rect 8169 67973 8255 68029
rect 8311 67973 8397 68029
rect 8453 67973 8539 68029
rect 8595 67973 8681 68029
rect 8737 67973 8823 68029
rect 8879 67973 8965 68029
rect 9021 67973 9107 68029
rect 9163 67973 9249 68029
rect 9305 67973 9391 68029
rect 9447 67973 9533 68029
rect 9589 67973 9675 68029
rect 9731 67973 9817 68029
rect 9873 67973 9959 68029
rect 10015 67973 10101 68029
rect 10157 67973 10243 68029
rect 10299 67973 10385 68029
rect 10441 67973 10527 68029
rect 10583 67973 10669 68029
rect 10725 67973 10811 68029
rect 10867 67973 10953 68029
rect 11009 67973 11095 68029
rect 11151 67973 11237 68029
rect 11293 67973 11379 68029
rect 11435 67973 11521 68029
rect 11577 67973 11663 68029
rect 11719 67973 11805 68029
rect 11861 67973 11947 68029
rect 12003 67973 12089 68029
rect 12145 67973 12231 68029
rect 12287 67973 12373 68029
rect 12429 67973 12515 68029
rect 12571 67973 12657 68029
rect 12713 67973 12799 68029
rect 12855 67973 12941 68029
rect 12997 67973 13083 68029
rect 13139 67973 13225 68029
rect 13281 67973 13367 68029
rect 13423 67973 13509 68029
rect 13565 67973 13651 68029
rect 13707 67973 13793 68029
rect 13849 67973 13935 68029
rect 13991 67973 14077 68029
rect 14133 67973 14219 68029
rect 14275 67973 14361 68029
rect 14417 67973 14503 68029
rect 14559 67973 14645 68029
rect 14701 67973 14787 68029
rect 14843 67973 15000 68029
rect 0 67887 15000 67973
rect 0 67831 161 67887
rect 217 67831 303 67887
rect 359 67831 445 67887
rect 501 67831 587 67887
rect 643 67831 729 67887
rect 785 67831 871 67887
rect 927 67831 1013 67887
rect 1069 67831 1155 67887
rect 1211 67831 1297 67887
rect 1353 67831 1439 67887
rect 1495 67831 1581 67887
rect 1637 67831 1723 67887
rect 1779 67831 1865 67887
rect 1921 67831 2007 67887
rect 2063 67831 2149 67887
rect 2205 67831 2291 67887
rect 2347 67831 2433 67887
rect 2489 67831 2575 67887
rect 2631 67831 2717 67887
rect 2773 67831 2859 67887
rect 2915 67831 3001 67887
rect 3057 67831 3143 67887
rect 3199 67831 3285 67887
rect 3341 67831 3427 67887
rect 3483 67831 3569 67887
rect 3625 67831 3711 67887
rect 3767 67831 3853 67887
rect 3909 67831 3995 67887
rect 4051 67831 4137 67887
rect 4193 67831 4279 67887
rect 4335 67831 4421 67887
rect 4477 67831 4563 67887
rect 4619 67831 4705 67887
rect 4761 67831 4847 67887
rect 4903 67831 4989 67887
rect 5045 67831 5131 67887
rect 5187 67831 5273 67887
rect 5329 67831 5415 67887
rect 5471 67831 5557 67887
rect 5613 67831 5699 67887
rect 5755 67831 5841 67887
rect 5897 67831 5983 67887
rect 6039 67831 6125 67887
rect 6181 67831 6267 67887
rect 6323 67831 6409 67887
rect 6465 67831 6551 67887
rect 6607 67831 6693 67887
rect 6749 67831 6835 67887
rect 6891 67831 6977 67887
rect 7033 67831 7119 67887
rect 7175 67831 7261 67887
rect 7317 67831 7403 67887
rect 7459 67831 7545 67887
rect 7601 67831 7687 67887
rect 7743 67831 7829 67887
rect 7885 67831 7971 67887
rect 8027 67831 8113 67887
rect 8169 67831 8255 67887
rect 8311 67831 8397 67887
rect 8453 67831 8539 67887
rect 8595 67831 8681 67887
rect 8737 67831 8823 67887
rect 8879 67831 8965 67887
rect 9021 67831 9107 67887
rect 9163 67831 9249 67887
rect 9305 67831 9391 67887
rect 9447 67831 9533 67887
rect 9589 67831 9675 67887
rect 9731 67831 9817 67887
rect 9873 67831 9959 67887
rect 10015 67831 10101 67887
rect 10157 67831 10243 67887
rect 10299 67831 10385 67887
rect 10441 67831 10527 67887
rect 10583 67831 10669 67887
rect 10725 67831 10811 67887
rect 10867 67831 10953 67887
rect 11009 67831 11095 67887
rect 11151 67831 11237 67887
rect 11293 67831 11379 67887
rect 11435 67831 11521 67887
rect 11577 67831 11663 67887
rect 11719 67831 11805 67887
rect 11861 67831 11947 67887
rect 12003 67831 12089 67887
rect 12145 67831 12231 67887
rect 12287 67831 12373 67887
rect 12429 67831 12515 67887
rect 12571 67831 12657 67887
rect 12713 67831 12799 67887
rect 12855 67831 12941 67887
rect 12997 67831 13083 67887
rect 13139 67831 13225 67887
rect 13281 67831 13367 67887
rect 13423 67831 13509 67887
rect 13565 67831 13651 67887
rect 13707 67831 13793 67887
rect 13849 67831 13935 67887
rect 13991 67831 14077 67887
rect 14133 67831 14219 67887
rect 14275 67831 14361 67887
rect 14417 67831 14503 67887
rect 14559 67831 14645 67887
rect 14701 67831 14787 67887
rect 14843 67831 15000 67887
rect 0 67745 15000 67831
rect 0 67689 161 67745
rect 217 67689 303 67745
rect 359 67689 445 67745
rect 501 67689 587 67745
rect 643 67689 729 67745
rect 785 67689 871 67745
rect 927 67689 1013 67745
rect 1069 67689 1155 67745
rect 1211 67689 1297 67745
rect 1353 67689 1439 67745
rect 1495 67689 1581 67745
rect 1637 67689 1723 67745
rect 1779 67689 1865 67745
rect 1921 67689 2007 67745
rect 2063 67689 2149 67745
rect 2205 67689 2291 67745
rect 2347 67689 2433 67745
rect 2489 67689 2575 67745
rect 2631 67689 2717 67745
rect 2773 67689 2859 67745
rect 2915 67689 3001 67745
rect 3057 67689 3143 67745
rect 3199 67689 3285 67745
rect 3341 67689 3427 67745
rect 3483 67689 3569 67745
rect 3625 67689 3711 67745
rect 3767 67689 3853 67745
rect 3909 67689 3995 67745
rect 4051 67689 4137 67745
rect 4193 67689 4279 67745
rect 4335 67689 4421 67745
rect 4477 67689 4563 67745
rect 4619 67689 4705 67745
rect 4761 67689 4847 67745
rect 4903 67689 4989 67745
rect 5045 67689 5131 67745
rect 5187 67689 5273 67745
rect 5329 67689 5415 67745
rect 5471 67689 5557 67745
rect 5613 67689 5699 67745
rect 5755 67689 5841 67745
rect 5897 67689 5983 67745
rect 6039 67689 6125 67745
rect 6181 67689 6267 67745
rect 6323 67689 6409 67745
rect 6465 67689 6551 67745
rect 6607 67689 6693 67745
rect 6749 67689 6835 67745
rect 6891 67689 6977 67745
rect 7033 67689 7119 67745
rect 7175 67689 7261 67745
rect 7317 67689 7403 67745
rect 7459 67689 7545 67745
rect 7601 67689 7687 67745
rect 7743 67689 7829 67745
rect 7885 67689 7971 67745
rect 8027 67689 8113 67745
rect 8169 67689 8255 67745
rect 8311 67689 8397 67745
rect 8453 67689 8539 67745
rect 8595 67689 8681 67745
rect 8737 67689 8823 67745
rect 8879 67689 8965 67745
rect 9021 67689 9107 67745
rect 9163 67689 9249 67745
rect 9305 67689 9391 67745
rect 9447 67689 9533 67745
rect 9589 67689 9675 67745
rect 9731 67689 9817 67745
rect 9873 67689 9959 67745
rect 10015 67689 10101 67745
rect 10157 67689 10243 67745
rect 10299 67689 10385 67745
rect 10441 67689 10527 67745
rect 10583 67689 10669 67745
rect 10725 67689 10811 67745
rect 10867 67689 10953 67745
rect 11009 67689 11095 67745
rect 11151 67689 11237 67745
rect 11293 67689 11379 67745
rect 11435 67689 11521 67745
rect 11577 67689 11663 67745
rect 11719 67689 11805 67745
rect 11861 67689 11947 67745
rect 12003 67689 12089 67745
rect 12145 67689 12231 67745
rect 12287 67689 12373 67745
rect 12429 67689 12515 67745
rect 12571 67689 12657 67745
rect 12713 67689 12799 67745
rect 12855 67689 12941 67745
rect 12997 67689 13083 67745
rect 13139 67689 13225 67745
rect 13281 67689 13367 67745
rect 13423 67689 13509 67745
rect 13565 67689 13651 67745
rect 13707 67689 13793 67745
rect 13849 67689 13935 67745
rect 13991 67689 14077 67745
rect 14133 67689 14219 67745
rect 14275 67689 14361 67745
rect 14417 67689 14503 67745
rect 14559 67689 14645 67745
rect 14701 67689 14787 67745
rect 14843 67689 15000 67745
rect 0 67603 15000 67689
rect 0 67547 161 67603
rect 217 67547 303 67603
rect 359 67547 445 67603
rect 501 67547 587 67603
rect 643 67547 729 67603
rect 785 67547 871 67603
rect 927 67547 1013 67603
rect 1069 67547 1155 67603
rect 1211 67547 1297 67603
rect 1353 67547 1439 67603
rect 1495 67547 1581 67603
rect 1637 67547 1723 67603
rect 1779 67547 1865 67603
rect 1921 67547 2007 67603
rect 2063 67547 2149 67603
rect 2205 67547 2291 67603
rect 2347 67547 2433 67603
rect 2489 67547 2575 67603
rect 2631 67547 2717 67603
rect 2773 67547 2859 67603
rect 2915 67547 3001 67603
rect 3057 67547 3143 67603
rect 3199 67547 3285 67603
rect 3341 67547 3427 67603
rect 3483 67547 3569 67603
rect 3625 67547 3711 67603
rect 3767 67547 3853 67603
rect 3909 67547 3995 67603
rect 4051 67547 4137 67603
rect 4193 67547 4279 67603
rect 4335 67547 4421 67603
rect 4477 67547 4563 67603
rect 4619 67547 4705 67603
rect 4761 67547 4847 67603
rect 4903 67547 4989 67603
rect 5045 67547 5131 67603
rect 5187 67547 5273 67603
rect 5329 67547 5415 67603
rect 5471 67547 5557 67603
rect 5613 67547 5699 67603
rect 5755 67547 5841 67603
rect 5897 67547 5983 67603
rect 6039 67547 6125 67603
rect 6181 67547 6267 67603
rect 6323 67547 6409 67603
rect 6465 67547 6551 67603
rect 6607 67547 6693 67603
rect 6749 67547 6835 67603
rect 6891 67547 6977 67603
rect 7033 67547 7119 67603
rect 7175 67547 7261 67603
rect 7317 67547 7403 67603
rect 7459 67547 7545 67603
rect 7601 67547 7687 67603
rect 7743 67547 7829 67603
rect 7885 67547 7971 67603
rect 8027 67547 8113 67603
rect 8169 67547 8255 67603
rect 8311 67547 8397 67603
rect 8453 67547 8539 67603
rect 8595 67547 8681 67603
rect 8737 67547 8823 67603
rect 8879 67547 8965 67603
rect 9021 67547 9107 67603
rect 9163 67547 9249 67603
rect 9305 67547 9391 67603
rect 9447 67547 9533 67603
rect 9589 67547 9675 67603
rect 9731 67547 9817 67603
rect 9873 67547 9959 67603
rect 10015 67547 10101 67603
rect 10157 67547 10243 67603
rect 10299 67547 10385 67603
rect 10441 67547 10527 67603
rect 10583 67547 10669 67603
rect 10725 67547 10811 67603
rect 10867 67547 10953 67603
rect 11009 67547 11095 67603
rect 11151 67547 11237 67603
rect 11293 67547 11379 67603
rect 11435 67547 11521 67603
rect 11577 67547 11663 67603
rect 11719 67547 11805 67603
rect 11861 67547 11947 67603
rect 12003 67547 12089 67603
rect 12145 67547 12231 67603
rect 12287 67547 12373 67603
rect 12429 67547 12515 67603
rect 12571 67547 12657 67603
rect 12713 67547 12799 67603
rect 12855 67547 12941 67603
rect 12997 67547 13083 67603
rect 13139 67547 13225 67603
rect 13281 67547 13367 67603
rect 13423 67547 13509 67603
rect 13565 67547 13651 67603
rect 13707 67547 13793 67603
rect 13849 67547 13935 67603
rect 13991 67547 14077 67603
rect 14133 67547 14219 67603
rect 14275 67547 14361 67603
rect 14417 67547 14503 67603
rect 14559 67547 14645 67603
rect 14701 67547 14787 67603
rect 14843 67547 15000 67603
rect 0 67461 15000 67547
rect 0 67405 161 67461
rect 217 67405 303 67461
rect 359 67405 445 67461
rect 501 67405 587 67461
rect 643 67405 729 67461
rect 785 67405 871 67461
rect 927 67405 1013 67461
rect 1069 67405 1155 67461
rect 1211 67405 1297 67461
rect 1353 67405 1439 67461
rect 1495 67405 1581 67461
rect 1637 67405 1723 67461
rect 1779 67405 1865 67461
rect 1921 67405 2007 67461
rect 2063 67405 2149 67461
rect 2205 67405 2291 67461
rect 2347 67405 2433 67461
rect 2489 67405 2575 67461
rect 2631 67405 2717 67461
rect 2773 67405 2859 67461
rect 2915 67405 3001 67461
rect 3057 67405 3143 67461
rect 3199 67405 3285 67461
rect 3341 67405 3427 67461
rect 3483 67405 3569 67461
rect 3625 67405 3711 67461
rect 3767 67405 3853 67461
rect 3909 67405 3995 67461
rect 4051 67405 4137 67461
rect 4193 67405 4279 67461
rect 4335 67405 4421 67461
rect 4477 67405 4563 67461
rect 4619 67405 4705 67461
rect 4761 67405 4847 67461
rect 4903 67405 4989 67461
rect 5045 67405 5131 67461
rect 5187 67405 5273 67461
rect 5329 67405 5415 67461
rect 5471 67405 5557 67461
rect 5613 67405 5699 67461
rect 5755 67405 5841 67461
rect 5897 67405 5983 67461
rect 6039 67405 6125 67461
rect 6181 67405 6267 67461
rect 6323 67405 6409 67461
rect 6465 67405 6551 67461
rect 6607 67405 6693 67461
rect 6749 67405 6835 67461
rect 6891 67405 6977 67461
rect 7033 67405 7119 67461
rect 7175 67405 7261 67461
rect 7317 67405 7403 67461
rect 7459 67405 7545 67461
rect 7601 67405 7687 67461
rect 7743 67405 7829 67461
rect 7885 67405 7971 67461
rect 8027 67405 8113 67461
rect 8169 67405 8255 67461
rect 8311 67405 8397 67461
rect 8453 67405 8539 67461
rect 8595 67405 8681 67461
rect 8737 67405 8823 67461
rect 8879 67405 8965 67461
rect 9021 67405 9107 67461
rect 9163 67405 9249 67461
rect 9305 67405 9391 67461
rect 9447 67405 9533 67461
rect 9589 67405 9675 67461
rect 9731 67405 9817 67461
rect 9873 67405 9959 67461
rect 10015 67405 10101 67461
rect 10157 67405 10243 67461
rect 10299 67405 10385 67461
rect 10441 67405 10527 67461
rect 10583 67405 10669 67461
rect 10725 67405 10811 67461
rect 10867 67405 10953 67461
rect 11009 67405 11095 67461
rect 11151 67405 11237 67461
rect 11293 67405 11379 67461
rect 11435 67405 11521 67461
rect 11577 67405 11663 67461
rect 11719 67405 11805 67461
rect 11861 67405 11947 67461
rect 12003 67405 12089 67461
rect 12145 67405 12231 67461
rect 12287 67405 12373 67461
rect 12429 67405 12515 67461
rect 12571 67405 12657 67461
rect 12713 67405 12799 67461
rect 12855 67405 12941 67461
rect 12997 67405 13083 67461
rect 13139 67405 13225 67461
rect 13281 67405 13367 67461
rect 13423 67405 13509 67461
rect 13565 67405 13651 67461
rect 13707 67405 13793 67461
rect 13849 67405 13935 67461
rect 13991 67405 14077 67461
rect 14133 67405 14219 67461
rect 14275 67405 14361 67461
rect 14417 67405 14503 67461
rect 14559 67405 14645 67461
rect 14701 67405 14787 67461
rect 14843 67405 15000 67461
rect 0 67319 15000 67405
rect 0 67263 161 67319
rect 217 67263 303 67319
rect 359 67263 445 67319
rect 501 67263 587 67319
rect 643 67263 729 67319
rect 785 67263 871 67319
rect 927 67263 1013 67319
rect 1069 67263 1155 67319
rect 1211 67263 1297 67319
rect 1353 67263 1439 67319
rect 1495 67263 1581 67319
rect 1637 67263 1723 67319
rect 1779 67263 1865 67319
rect 1921 67263 2007 67319
rect 2063 67263 2149 67319
rect 2205 67263 2291 67319
rect 2347 67263 2433 67319
rect 2489 67263 2575 67319
rect 2631 67263 2717 67319
rect 2773 67263 2859 67319
rect 2915 67263 3001 67319
rect 3057 67263 3143 67319
rect 3199 67263 3285 67319
rect 3341 67263 3427 67319
rect 3483 67263 3569 67319
rect 3625 67263 3711 67319
rect 3767 67263 3853 67319
rect 3909 67263 3995 67319
rect 4051 67263 4137 67319
rect 4193 67263 4279 67319
rect 4335 67263 4421 67319
rect 4477 67263 4563 67319
rect 4619 67263 4705 67319
rect 4761 67263 4847 67319
rect 4903 67263 4989 67319
rect 5045 67263 5131 67319
rect 5187 67263 5273 67319
rect 5329 67263 5415 67319
rect 5471 67263 5557 67319
rect 5613 67263 5699 67319
rect 5755 67263 5841 67319
rect 5897 67263 5983 67319
rect 6039 67263 6125 67319
rect 6181 67263 6267 67319
rect 6323 67263 6409 67319
rect 6465 67263 6551 67319
rect 6607 67263 6693 67319
rect 6749 67263 6835 67319
rect 6891 67263 6977 67319
rect 7033 67263 7119 67319
rect 7175 67263 7261 67319
rect 7317 67263 7403 67319
rect 7459 67263 7545 67319
rect 7601 67263 7687 67319
rect 7743 67263 7829 67319
rect 7885 67263 7971 67319
rect 8027 67263 8113 67319
rect 8169 67263 8255 67319
rect 8311 67263 8397 67319
rect 8453 67263 8539 67319
rect 8595 67263 8681 67319
rect 8737 67263 8823 67319
rect 8879 67263 8965 67319
rect 9021 67263 9107 67319
rect 9163 67263 9249 67319
rect 9305 67263 9391 67319
rect 9447 67263 9533 67319
rect 9589 67263 9675 67319
rect 9731 67263 9817 67319
rect 9873 67263 9959 67319
rect 10015 67263 10101 67319
rect 10157 67263 10243 67319
rect 10299 67263 10385 67319
rect 10441 67263 10527 67319
rect 10583 67263 10669 67319
rect 10725 67263 10811 67319
rect 10867 67263 10953 67319
rect 11009 67263 11095 67319
rect 11151 67263 11237 67319
rect 11293 67263 11379 67319
rect 11435 67263 11521 67319
rect 11577 67263 11663 67319
rect 11719 67263 11805 67319
rect 11861 67263 11947 67319
rect 12003 67263 12089 67319
rect 12145 67263 12231 67319
rect 12287 67263 12373 67319
rect 12429 67263 12515 67319
rect 12571 67263 12657 67319
rect 12713 67263 12799 67319
rect 12855 67263 12941 67319
rect 12997 67263 13083 67319
rect 13139 67263 13225 67319
rect 13281 67263 13367 67319
rect 13423 67263 13509 67319
rect 13565 67263 13651 67319
rect 13707 67263 13793 67319
rect 13849 67263 13935 67319
rect 13991 67263 14077 67319
rect 14133 67263 14219 67319
rect 14275 67263 14361 67319
rect 14417 67263 14503 67319
rect 14559 67263 14645 67319
rect 14701 67263 14787 67319
rect 14843 67263 15000 67319
rect 0 67177 15000 67263
rect 0 67121 161 67177
rect 217 67121 303 67177
rect 359 67121 445 67177
rect 501 67121 587 67177
rect 643 67121 729 67177
rect 785 67121 871 67177
rect 927 67121 1013 67177
rect 1069 67121 1155 67177
rect 1211 67121 1297 67177
rect 1353 67121 1439 67177
rect 1495 67121 1581 67177
rect 1637 67121 1723 67177
rect 1779 67121 1865 67177
rect 1921 67121 2007 67177
rect 2063 67121 2149 67177
rect 2205 67121 2291 67177
rect 2347 67121 2433 67177
rect 2489 67121 2575 67177
rect 2631 67121 2717 67177
rect 2773 67121 2859 67177
rect 2915 67121 3001 67177
rect 3057 67121 3143 67177
rect 3199 67121 3285 67177
rect 3341 67121 3427 67177
rect 3483 67121 3569 67177
rect 3625 67121 3711 67177
rect 3767 67121 3853 67177
rect 3909 67121 3995 67177
rect 4051 67121 4137 67177
rect 4193 67121 4279 67177
rect 4335 67121 4421 67177
rect 4477 67121 4563 67177
rect 4619 67121 4705 67177
rect 4761 67121 4847 67177
rect 4903 67121 4989 67177
rect 5045 67121 5131 67177
rect 5187 67121 5273 67177
rect 5329 67121 5415 67177
rect 5471 67121 5557 67177
rect 5613 67121 5699 67177
rect 5755 67121 5841 67177
rect 5897 67121 5983 67177
rect 6039 67121 6125 67177
rect 6181 67121 6267 67177
rect 6323 67121 6409 67177
rect 6465 67121 6551 67177
rect 6607 67121 6693 67177
rect 6749 67121 6835 67177
rect 6891 67121 6977 67177
rect 7033 67121 7119 67177
rect 7175 67121 7261 67177
rect 7317 67121 7403 67177
rect 7459 67121 7545 67177
rect 7601 67121 7687 67177
rect 7743 67121 7829 67177
rect 7885 67121 7971 67177
rect 8027 67121 8113 67177
rect 8169 67121 8255 67177
rect 8311 67121 8397 67177
rect 8453 67121 8539 67177
rect 8595 67121 8681 67177
rect 8737 67121 8823 67177
rect 8879 67121 8965 67177
rect 9021 67121 9107 67177
rect 9163 67121 9249 67177
rect 9305 67121 9391 67177
rect 9447 67121 9533 67177
rect 9589 67121 9675 67177
rect 9731 67121 9817 67177
rect 9873 67121 9959 67177
rect 10015 67121 10101 67177
rect 10157 67121 10243 67177
rect 10299 67121 10385 67177
rect 10441 67121 10527 67177
rect 10583 67121 10669 67177
rect 10725 67121 10811 67177
rect 10867 67121 10953 67177
rect 11009 67121 11095 67177
rect 11151 67121 11237 67177
rect 11293 67121 11379 67177
rect 11435 67121 11521 67177
rect 11577 67121 11663 67177
rect 11719 67121 11805 67177
rect 11861 67121 11947 67177
rect 12003 67121 12089 67177
rect 12145 67121 12231 67177
rect 12287 67121 12373 67177
rect 12429 67121 12515 67177
rect 12571 67121 12657 67177
rect 12713 67121 12799 67177
rect 12855 67121 12941 67177
rect 12997 67121 13083 67177
rect 13139 67121 13225 67177
rect 13281 67121 13367 67177
rect 13423 67121 13509 67177
rect 13565 67121 13651 67177
rect 13707 67121 13793 67177
rect 13849 67121 13935 67177
rect 13991 67121 14077 67177
rect 14133 67121 14219 67177
rect 14275 67121 14361 67177
rect 14417 67121 14503 67177
rect 14559 67121 14645 67177
rect 14701 67121 14787 67177
rect 14843 67121 15000 67177
rect 0 67035 15000 67121
rect 0 66979 161 67035
rect 217 66979 303 67035
rect 359 66979 445 67035
rect 501 66979 587 67035
rect 643 66979 729 67035
rect 785 66979 871 67035
rect 927 66979 1013 67035
rect 1069 66979 1155 67035
rect 1211 66979 1297 67035
rect 1353 66979 1439 67035
rect 1495 66979 1581 67035
rect 1637 66979 1723 67035
rect 1779 66979 1865 67035
rect 1921 66979 2007 67035
rect 2063 66979 2149 67035
rect 2205 66979 2291 67035
rect 2347 66979 2433 67035
rect 2489 66979 2575 67035
rect 2631 66979 2717 67035
rect 2773 66979 2859 67035
rect 2915 66979 3001 67035
rect 3057 66979 3143 67035
rect 3199 66979 3285 67035
rect 3341 66979 3427 67035
rect 3483 66979 3569 67035
rect 3625 66979 3711 67035
rect 3767 66979 3853 67035
rect 3909 66979 3995 67035
rect 4051 66979 4137 67035
rect 4193 66979 4279 67035
rect 4335 66979 4421 67035
rect 4477 66979 4563 67035
rect 4619 66979 4705 67035
rect 4761 66979 4847 67035
rect 4903 66979 4989 67035
rect 5045 66979 5131 67035
rect 5187 66979 5273 67035
rect 5329 66979 5415 67035
rect 5471 66979 5557 67035
rect 5613 66979 5699 67035
rect 5755 66979 5841 67035
rect 5897 66979 5983 67035
rect 6039 66979 6125 67035
rect 6181 66979 6267 67035
rect 6323 66979 6409 67035
rect 6465 66979 6551 67035
rect 6607 66979 6693 67035
rect 6749 66979 6835 67035
rect 6891 66979 6977 67035
rect 7033 66979 7119 67035
rect 7175 66979 7261 67035
rect 7317 66979 7403 67035
rect 7459 66979 7545 67035
rect 7601 66979 7687 67035
rect 7743 66979 7829 67035
rect 7885 66979 7971 67035
rect 8027 66979 8113 67035
rect 8169 66979 8255 67035
rect 8311 66979 8397 67035
rect 8453 66979 8539 67035
rect 8595 66979 8681 67035
rect 8737 66979 8823 67035
rect 8879 66979 8965 67035
rect 9021 66979 9107 67035
rect 9163 66979 9249 67035
rect 9305 66979 9391 67035
rect 9447 66979 9533 67035
rect 9589 66979 9675 67035
rect 9731 66979 9817 67035
rect 9873 66979 9959 67035
rect 10015 66979 10101 67035
rect 10157 66979 10243 67035
rect 10299 66979 10385 67035
rect 10441 66979 10527 67035
rect 10583 66979 10669 67035
rect 10725 66979 10811 67035
rect 10867 66979 10953 67035
rect 11009 66979 11095 67035
rect 11151 66979 11237 67035
rect 11293 66979 11379 67035
rect 11435 66979 11521 67035
rect 11577 66979 11663 67035
rect 11719 66979 11805 67035
rect 11861 66979 11947 67035
rect 12003 66979 12089 67035
rect 12145 66979 12231 67035
rect 12287 66979 12373 67035
rect 12429 66979 12515 67035
rect 12571 66979 12657 67035
rect 12713 66979 12799 67035
rect 12855 66979 12941 67035
rect 12997 66979 13083 67035
rect 13139 66979 13225 67035
rect 13281 66979 13367 67035
rect 13423 66979 13509 67035
rect 13565 66979 13651 67035
rect 13707 66979 13793 67035
rect 13849 66979 13935 67035
rect 13991 66979 14077 67035
rect 14133 66979 14219 67035
rect 14275 66979 14361 67035
rect 14417 66979 14503 67035
rect 14559 66979 14645 67035
rect 14701 66979 14787 67035
rect 14843 66979 15000 67035
rect 0 66893 15000 66979
rect 0 66837 161 66893
rect 217 66837 303 66893
rect 359 66837 445 66893
rect 501 66837 587 66893
rect 643 66837 729 66893
rect 785 66837 871 66893
rect 927 66837 1013 66893
rect 1069 66837 1155 66893
rect 1211 66837 1297 66893
rect 1353 66837 1439 66893
rect 1495 66837 1581 66893
rect 1637 66837 1723 66893
rect 1779 66837 1865 66893
rect 1921 66837 2007 66893
rect 2063 66837 2149 66893
rect 2205 66837 2291 66893
rect 2347 66837 2433 66893
rect 2489 66837 2575 66893
rect 2631 66837 2717 66893
rect 2773 66837 2859 66893
rect 2915 66837 3001 66893
rect 3057 66837 3143 66893
rect 3199 66837 3285 66893
rect 3341 66837 3427 66893
rect 3483 66837 3569 66893
rect 3625 66837 3711 66893
rect 3767 66837 3853 66893
rect 3909 66837 3995 66893
rect 4051 66837 4137 66893
rect 4193 66837 4279 66893
rect 4335 66837 4421 66893
rect 4477 66837 4563 66893
rect 4619 66837 4705 66893
rect 4761 66837 4847 66893
rect 4903 66837 4989 66893
rect 5045 66837 5131 66893
rect 5187 66837 5273 66893
rect 5329 66837 5415 66893
rect 5471 66837 5557 66893
rect 5613 66837 5699 66893
rect 5755 66837 5841 66893
rect 5897 66837 5983 66893
rect 6039 66837 6125 66893
rect 6181 66837 6267 66893
rect 6323 66837 6409 66893
rect 6465 66837 6551 66893
rect 6607 66837 6693 66893
rect 6749 66837 6835 66893
rect 6891 66837 6977 66893
rect 7033 66837 7119 66893
rect 7175 66837 7261 66893
rect 7317 66837 7403 66893
rect 7459 66837 7545 66893
rect 7601 66837 7687 66893
rect 7743 66837 7829 66893
rect 7885 66837 7971 66893
rect 8027 66837 8113 66893
rect 8169 66837 8255 66893
rect 8311 66837 8397 66893
rect 8453 66837 8539 66893
rect 8595 66837 8681 66893
rect 8737 66837 8823 66893
rect 8879 66837 8965 66893
rect 9021 66837 9107 66893
rect 9163 66837 9249 66893
rect 9305 66837 9391 66893
rect 9447 66837 9533 66893
rect 9589 66837 9675 66893
rect 9731 66837 9817 66893
rect 9873 66837 9959 66893
rect 10015 66837 10101 66893
rect 10157 66837 10243 66893
rect 10299 66837 10385 66893
rect 10441 66837 10527 66893
rect 10583 66837 10669 66893
rect 10725 66837 10811 66893
rect 10867 66837 10953 66893
rect 11009 66837 11095 66893
rect 11151 66837 11237 66893
rect 11293 66837 11379 66893
rect 11435 66837 11521 66893
rect 11577 66837 11663 66893
rect 11719 66837 11805 66893
rect 11861 66837 11947 66893
rect 12003 66837 12089 66893
rect 12145 66837 12231 66893
rect 12287 66837 12373 66893
rect 12429 66837 12515 66893
rect 12571 66837 12657 66893
rect 12713 66837 12799 66893
rect 12855 66837 12941 66893
rect 12997 66837 13083 66893
rect 13139 66837 13225 66893
rect 13281 66837 13367 66893
rect 13423 66837 13509 66893
rect 13565 66837 13651 66893
rect 13707 66837 13793 66893
rect 13849 66837 13935 66893
rect 13991 66837 14077 66893
rect 14133 66837 14219 66893
rect 14275 66837 14361 66893
rect 14417 66837 14503 66893
rect 14559 66837 14645 66893
rect 14701 66837 14787 66893
rect 14843 66837 15000 66893
rect 0 66800 15000 66837
rect 0 66571 15000 66600
rect 0 66515 161 66571
rect 217 66515 303 66571
rect 359 66515 445 66571
rect 501 66515 587 66571
rect 643 66515 729 66571
rect 785 66515 871 66571
rect 927 66515 1013 66571
rect 1069 66515 1155 66571
rect 1211 66515 1297 66571
rect 1353 66515 1439 66571
rect 1495 66515 1581 66571
rect 1637 66515 1723 66571
rect 1779 66515 1865 66571
rect 1921 66515 2007 66571
rect 2063 66515 2149 66571
rect 2205 66515 2291 66571
rect 2347 66515 2433 66571
rect 2489 66515 2575 66571
rect 2631 66515 2717 66571
rect 2773 66515 2859 66571
rect 2915 66515 3001 66571
rect 3057 66515 3143 66571
rect 3199 66515 3285 66571
rect 3341 66515 3427 66571
rect 3483 66515 3569 66571
rect 3625 66515 3711 66571
rect 3767 66515 3853 66571
rect 3909 66515 3995 66571
rect 4051 66515 4137 66571
rect 4193 66515 4279 66571
rect 4335 66515 4421 66571
rect 4477 66515 4563 66571
rect 4619 66515 4705 66571
rect 4761 66515 4847 66571
rect 4903 66515 4989 66571
rect 5045 66515 5131 66571
rect 5187 66515 5273 66571
rect 5329 66515 5415 66571
rect 5471 66515 5557 66571
rect 5613 66515 5699 66571
rect 5755 66515 5841 66571
rect 5897 66515 5983 66571
rect 6039 66515 6125 66571
rect 6181 66515 6267 66571
rect 6323 66515 6409 66571
rect 6465 66515 6551 66571
rect 6607 66515 6693 66571
rect 6749 66515 6835 66571
rect 6891 66515 6977 66571
rect 7033 66515 7119 66571
rect 7175 66515 7261 66571
rect 7317 66515 7403 66571
rect 7459 66515 7545 66571
rect 7601 66515 7687 66571
rect 7743 66515 7829 66571
rect 7885 66515 7971 66571
rect 8027 66515 8113 66571
rect 8169 66515 8255 66571
rect 8311 66515 8397 66571
rect 8453 66515 8539 66571
rect 8595 66515 8681 66571
rect 8737 66515 8823 66571
rect 8879 66515 8965 66571
rect 9021 66515 9107 66571
rect 9163 66515 9249 66571
rect 9305 66515 9391 66571
rect 9447 66515 9533 66571
rect 9589 66515 9675 66571
rect 9731 66515 9817 66571
rect 9873 66515 9959 66571
rect 10015 66515 10101 66571
rect 10157 66515 10243 66571
rect 10299 66515 10385 66571
rect 10441 66515 10527 66571
rect 10583 66515 10669 66571
rect 10725 66515 10811 66571
rect 10867 66515 10953 66571
rect 11009 66515 11095 66571
rect 11151 66515 11237 66571
rect 11293 66515 11379 66571
rect 11435 66515 11521 66571
rect 11577 66515 11663 66571
rect 11719 66515 11805 66571
rect 11861 66515 11947 66571
rect 12003 66515 12089 66571
rect 12145 66515 12231 66571
rect 12287 66515 12373 66571
rect 12429 66515 12515 66571
rect 12571 66515 12657 66571
rect 12713 66515 12799 66571
rect 12855 66515 12941 66571
rect 12997 66515 13083 66571
rect 13139 66515 13225 66571
rect 13281 66515 13367 66571
rect 13423 66515 13509 66571
rect 13565 66515 13651 66571
rect 13707 66515 13793 66571
rect 13849 66515 13935 66571
rect 13991 66515 14077 66571
rect 14133 66515 14219 66571
rect 14275 66515 14361 66571
rect 14417 66515 14503 66571
rect 14559 66515 14645 66571
rect 14701 66515 14787 66571
rect 14843 66515 15000 66571
rect 0 66429 15000 66515
rect 0 66373 161 66429
rect 217 66373 303 66429
rect 359 66373 445 66429
rect 501 66373 587 66429
rect 643 66373 729 66429
rect 785 66373 871 66429
rect 927 66373 1013 66429
rect 1069 66373 1155 66429
rect 1211 66373 1297 66429
rect 1353 66373 1439 66429
rect 1495 66373 1581 66429
rect 1637 66373 1723 66429
rect 1779 66373 1865 66429
rect 1921 66373 2007 66429
rect 2063 66373 2149 66429
rect 2205 66373 2291 66429
rect 2347 66373 2433 66429
rect 2489 66373 2575 66429
rect 2631 66373 2717 66429
rect 2773 66373 2859 66429
rect 2915 66373 3001 66429
rect 3057 66373 3143 66429
rect 3199 66373 3285 66429
rect 3341 66373 3427 66429
rect 3483 66373 3569 66429
rect 3625 66373 3711 66429
rect 3767 66373 3853 66429
rect 3909 66373 3995 66429
rect 4051 66373 4137 66429
rect 4193 66373 4279 66429
rect 4335 66373 4421 66429
rect 4477 66373 4563 66429
rect 4619 66373 4705 66429
rect 4761 66373 4847 66429
rect 4903 66373 4989 66429
rect 5045 66373 5131 66429
rect 5187 66373 5273 66429
rect 5329 66373 5415 66429
rect 5471 66373 5557 66429
rect 5613 66373 5699 66429
rect 5755 66373 5841 66429
rect 5897 66373 5983 66429
rect 6039 66373 6125 66429
rect 6181 66373 6267 66429
rect 6323 66373 6409 66429
rect 6465 66373 6551 66429
rect 6607 66373 6693 66429
rect 6749 66373 6835 66429
rect 6891 66373 6977 66429
rect 7033 66373 7119 66429
rect 7175 66373 7261 66429
rect 7317 66373 7403 66429
rect 7459 66373 7545 66429
rect 7601 66373 7687 66429
rect 7743 66373 7829 66429
rect 7885 66373 7971 66429
rect 8027 66373 8113 66429
rect 8169 66373 8255 66429
rect 8311 66373 8397 66429
rect 8453 66373 8539 66429
rect 8595 66373 8681 66429
rect 8737 66373 8823 66429
rect 8879 66373 8965 66429
rect 9021 66373 9107 66429
rect 9163 66373 9249 66429
rect 9305 66373 9391 66429
rect 9447 66373 9533 66429
rect 9589 66373 9675 66429
rect 9731 66373 9817 66429
rect 9873 66373 9959 66429
rect 10015 66373 10101 66429
rect 10157 66373 10243 66429
rect 10299 66373 10385 66429
rect 10441 66373 10527 66429
rect 10583 66373 10669 66429
rect 10725 66373 10811 66429
rect 10867 66373 10953 66429
rect 11009 66373 11095 66429
rect 11151 66373 11237 66429
rect 11293 66373 11379 66429
rect 11435 66373 11521 66429
rect 11577 66373 11663 66429
rect 11719 66373 11805 66429
rect 11861 66373 11947 66429
rect 12003 66373 12089 66429
rect 12145 66373 12231 66429
rect 12287 66373 12373 66429
rect 12429 66373 12515 66429
rect 12571 66373 12657 66429
rect 12713 66373 12799 66429
rect 12855 66373 12941 66429
rect 12997 66373 13083 66429
rect 13139 66373 13225 66429
rect 13281 66373 13367 66429
rect 13423 66373 13509 66429
rect 13565 66373 13651 66429
rect 13707 66373 13793 66429
rect 13849 66373 13935 66429
rect 13991 66373 14077 66429
rect 14133 66373 14219 66429
rect 14275 66373 14361 66429
rect 14417 66373 14503 66429
rect 14559 66373 14645 66429
rect 14701 66373 14787 66429
rect 14843 66373 15000 66429
rect 0 66287 15000 66373
rect 0 66231 161 66287
rect 217 66231 303 66287
rect 359 66231 445 66287
rect 501 66231 587 66287
rect 643 66231 729 66287
rect 785 66231 871 66287
rect 927 66231 1013 66287
rect 1069 66231 1155 66287
rect 1211 66231 1297 66287
rect 1353 66231 1439 66287
rect 1495 66231 1581 66287
rect 1637 66231 1723 66287
rect 1779 66231 1865 66287
rect 1921 66231 2007 66287
rect 2063 66231 2149 66287
rect 2205 66231 2291 66287
rect 2347 66231 2433 66287
rect 2489 66231 2575 66287
rect 2631 66231 2717 66287
rect 2773 66231 2859 66287
rect 2915 66231 3001 66287
rect 3057 66231 3143 66287
rect 3199 66231 3285 66287
rect 3341 66231 3427 66287
rect 3483 66231 3569 66287
rect 3625 66231 3711 66287
rect 3767 66231 3853 66287
rect 3909 66231 3995 66287
rect 4051 66231 4137 66287
rect 4193 66231 4279 66287
rect 4335 66231 4421 66287
rect 4477 66231 4563 66287
rect 4619 66231 4705 66287
rect 4761 66231 4847 66287
rect 4903 66231 4989 66287
rect 5045 66231 5131 66287
rect 5187 66231 5273 66287
rect 5329 66231 5415 66287
rect 5471 66231 5557 66287
rect 5613 66231 5699 66287
rect 5755 66231 5841 66287
rect 5897 66231 5983 66287
rect 6039 66231 6125 66287
rect 6181 66231 6267 66287
rect 6323 66231 6409 66287
rect 6465 66231 6551 66287
rect 6607 66231 6693 66287
rect 6749 66231 6835 66287
rect 6891 66231 6977 66287
rect 7033 66231 7119 66287
rect 7175 66231 7261 66287
rect 7317 66231 7403 66287
rect 7459 66231 7545 66287
rect 7601 66231 7687 66287
rect 7743 66231 7829 66287
rect 7885 66231 7971 66287
rect 8027 66231 8113 66287
rect 8169 66231 8255 66287
rect 8311 66231 8397 66287
rect 8453 66231 8539 66287
rect 8595 66231 8681 66287
rect 8737 66231 8823 66287
rect 8879 66231 8965 66287
rect 9021 66231 9107 66287
rect 9163 66231 9249 66287
rect 9305 66231 9391 66287
rect 9447 66231 9533 66287
rect 9589 66231 9675 66287
rect 9731 66231 9817 66287
rect 9873 66231 9959 66287
rect 10015 66231 10101 66287
rect 10157 66231 10243 66287
rect 10299 66231 10385 66287
rect 10441 66231 10527 66287
rect 10583 66231 10669 66287
rect 10725 66231 10811 66287
rect 10867 66231 10953 66287
rect 11009 66231 11095 66287
rect 11151 66231 11237 66287
rect 11293 66231 11379 66287
rect 11435 66231 11521 66287
rect 11577 66231 11663 66287
rect 11719 66231 11805 66287
rect 11861 66231 11947 66287
rect 12003 66231 12089 66287
rect 12145 66231 12231 66287
rect 12287 66231 12373 66287
rect 12429 66231 12515 66287
rect 12571 66231 12657 66287
rect 12713 66231 12799 66287
rect 12855 66231 12941 66287
rect 12997 66231 13083 66287
rect 13139 66231 13225 66287
rect 13281 66231 13367 66287
rect 13423 66231 13509 66287
rect 13565 66231 13651 66287
rect 13707 66231 13793 66287
rect 13849 66231 13935 66287
rect 13991 66231 14077 66287
rect 14133 66231 14219 66287
rect 14275 66231 14361 66287
rect 14417 66231 14503 66287
rect 14559 66231 14645 66287
rect 14701 66231 14787 66287
rect 14843 66231 15000 66287
rect 0 66145 15000 66231
rect 0 66089 161 66145
rect 217 66089 303 66145
rect 359 66089 445 66145
rect 501 66089 587 66145
rect 643 66089 729 66145
rect 785 66089 871 66145
rect 927 66089 1013 66145
rect 1069 66089 1155 66145
rect 1211 66089 1297 66145
rect 1353 66089 1439 66145
rect 1495 66089 1581 66145
rect 1637 66089 1723 66145
rect 1779 66089 1865 66145
rect 1921 66089 2007 66145
rect 2063 66089 2149 66145
rect 2205 66089 2291 66145
rect 2347 66089 2433 66145
rect 2489 66089 2575 66145
rect 2631 66089 2717 66145
rect 2773 66089 2859 66145
rect 2915 66089 3001 66145
rect 3057 66089 3143 66145
rect 3199 66089 3285 66145
rect 3341 66089 3427 66145
rect 3483 66089 3569 66145
rect 3625 66089 3711 66145
rect 3767 66089 3853 66145
rect 3909 66089 3995 66145
rect 4051 66089 4137 66145
rect 4193 66089 4279 66145
rect 4335 66089 4421 66145
rect 4477 66089 4563 66145
rect 4619 66089 4705 66145
rect 4761 66089 4847 66145
rect 4903 66089 4989 66145
rect 5045 66089 5131 66145
rect 5187 66089 5273 66145
rect 5329 66089 5415 66145
rect 5471 66089 5557 66145
rect 5613 66089 5699 66145
rect 5755 66089 5841 66145
rect 5897 66089 5983 66145
rect 6039 66089 6125 66145
rect 6181 66089 6267 66145
rect 6323 66089 6409 66145
rect 6465 66089 6551 66145
rect 6607 66089 6693 66145
rect 6749 66089 6835 66145
rect 6891 66089 6977 66145
rect 7033 66089 7119 66145
rect 7175 66089 7261 66145
rect 7317 66089 7403 66145
rect 7459 66089 7545 66145
rect 7601 66089 7687 66145
rect 7743 66089 7829 66145
rect 7885 66089 7971 66145
rect 8027 66089 8113 66145
rect 8169 66089 8255 66145
rect 8311 66089 8397 66145
rect 8453 66089 8539 66145
rect 8595 66089 8681 66145
rect 8737 66089 8823 66145
rect 8879 66089 8965 66145
rect 9021 66089 9107 66145
rect 9163 66089 9249 66145
rect 9305 66089 9391 66145
rect 9447 66089 9533 66145
rect 9589 66089 9675 66145
rect 9731 66089 9817 66145
rect 9873 66089 9959 66145
rect 10015 66089 10101 66145
rect 10157 66089 10243 66145
rect 10299 66089 10385 66145
rect 10441 66089 10527 66145
rect 10583 66089 10669 66145
rect 10725 66089 10811 66145
rect 10867 66089 10953 66145
rect 11009 66089 11095 66145
rect 11151 66089 11237 66145
rect 11293 66089 11379 66145
rect 11435 66089 11521 66145
rect 11577 66089 11663 66145
rect 11719 66089 11805 66145
rect 11861 66089 11947 66145
rect 12003 66089 12089 66145
rect 12145 66089 12231 66145
rect 12287 66089 12373 66145
rect 12429 66089 12515 66145
rect 12571 66089 12657 66145
rect 12713 66089 12799 66145
rect 12855 66089 12941 66145
rect 12997 66089 13083 66145
rect 13139 66089 13225 66145
rect 13281 66089 13367 66145
rect 13423 66089 13509 66145
rect 13565 66089 13651 66145
rect 13707 66089 13793 66145
rect 13849 66089 13935 66145
rect 13991 66089 14077 66145
rect 14133 66089 14219 66145
rect 14275 66089 14361 66145
rect 14417 66089 14503 66145
rect 14559 66089 14645 66145
rect 14701 66089 14787 66145
rect 14843 66089 15000 66145
rect 0 66003 15000 66089
rect 0 65947 161 66003
rect 217 65947 303 66003
rect 359 65947 445 66003
rect 501 65947 587 66003
rect 643 65947 729 66003
rect 785 65947 871 66003
rect 927 65947 1013 66003
rect 1069 65947 1155 66003
rect 1211 65947 1297 66003
rect 1353 65947 1439 66003
rect 1495 65947 1581 66003
rect 1637 65947 1723 66003
rect 1779 65947 1865 66003
rect 1921 65947 2007 66003
rect 2063 65947 2149 66003
rect 2205 65947 2291 66003
rect 2347 65947 2433 66003
rect 2489 65947 2575 66003
rect 2631 65947 2717 66003
rect 2773 65947 2859 66003
rect 2915 65947 3001 66003
rect 3057 65947 3143 66003
rect 3199 65947 3285 66003
rect 3341 65947 3427 66003
rect 3483 65947 3569 66003
rect 3625 65947 3711 66003
rect 3767 65947 3853 66003
rect 3909 65947 3995 66003
rect 4051 65947 4137 66003
rect 4193 65947 4279 66003
rect 4335 65947 4421 66003
rect 4477 65947 4563 66003
rect 4619 65947 4705 66003
rect 4761 65947 4847 66003
rect 4903 65947 4989 66003
rect 5045 65947 5131 66003
rect 5187 65947 5273 66003
rect 5329 65947 5415 66003
rect 5471 65947 5557 66003
rect 5613 65947 5699 66003
rect 5755 65947 5841 66003
rect 5897 65947 5983 66003
rect 6039 65947 6125 66003
rect 6181 65947 6267 66003
rect 6323 65947 6409 66003
rect 6465 65947 6551 66003
rect 6607 65947 6693 66003
rect 6749 65947 6835 66003
rect 6891 65947 6977 66003
rect 7033 65947 7119 66003
rect 7175 65947 7261 66003
rect 7317 65947 7403 66003
rect 7459 65947 7545 66003
rect 7601 65947 7687 66003
rect 7743 65947 7829 66003
rect 7885 65947 7971 66003
rect 8027 65947 8113 66003
rect 8169 65947 8255 66003
rect 8311 65947 8397 66003
rect 8453 65947 8539 66003
rect 8595 65947 8681 66003
rect 8737 65947 8823 66003
rect 8879 65947 8965 66003
rect 9021 65947 9107 66003
rect 9163 65947 9249 66003
rect 9305 65947 9391 66003
rect 9447 65947 9533 66003
rect 9589 65947 9675 66003
rect 9731 65947 9817 66003
rect 9873 65947 9959 66003
rect 10015 65947 10101 66003
rect 10157 65947 10243 66003
rect 10299 65947 10385 66003
rect 10441 65947 10527 66003
rect 10583 65947 10669 66003
rect 10725 65947 10811 66003
rect 10867 65947 10953 66003
rect 11009 65947 11095 66003
rect 11151 65947 11237 66003
rect 11293 65947 11379 66003
rect 11435 65947 11521 66003
rect 11577 65947 11663 66003
rect 11719 65947 11805 66003
rect 11861 65947 11947 66003
rect 12003 65947 12089 66003
rect 12145 65947 12231 66003
rect 12287 65947 12373 66003
rect 12429 65947 12515 66003
rect 12571 65947 12657 66003
rect 12713 65947 12799 66003
rect 12855 65947 12941 66003
rect 12997 65947 13083 66003
rect 13139 65947 13225 66003
rect 13281 65947 13367 66003
rect 13423 65947 13509 66003
rect 13565 65947 13651 66003
rect 13707 65947 13793 66003
rect 13849 65947 13935 66003
rect 13991 65947 14077 66003
rect 14133 65947 14219 66003
rect 14275 65947 14361 66003
rect 14417 65947 14503 66003
rect 14559 65947 14645 66003
rect 14701 65947 14787 66003
rect 14843 65947 15000 66003
rect 0 65861 15000 65947
rect 0 65805 161 65861
rect 217 65805 303 65861
rect 359 65805 445 65861
rect 501 65805 587 65861
rect 643 65805 729 65861
rect 785 65805 871 65861
rect 927 65805 1013 65861
rect 1069 65805 1155 65861
rect 1211 65805 1297 65861
rect 1353 65805 1439 65861
rect 1495 65805 1581 65861
rect 1637 65805 1723 65861
rect 1779 65805 1865 65861
rect 1921 65805 2007 65861
rect 2063 65805 2149 65861
rect 2205 65805 2291 65861
rect 2347 65805 2433 65861
rect 2489 65805 2575 65861
rect 2631 65805 2717 65861
rect 2773 65805 2859 65861
rect 2915 65805 3001 65861
rect 3057 65805 3143 65861
rect 3199 65805 3285 65861
rect 3341 65805 3427 65861
rect 3483 65805 3569 65861
rect 3625 65805 3711 65861
rect 3767 65805 3853 65861
rect 3909 65805 3995 65861
rect 4051 65805 4137 65861
rect 4193 65805 4279 65861
rect 4335 65805 4421 65861
rect 4477 65805 4563 65861
rect 4619 65805 4705 65861
rect 4761 65805 4847 65861
rect 4903 65805 4989 65861
rect 5045 65805 5131 65861
rect 5187 65805 5273 65861
rect 5329 65805 5415 65861
rect 5471 65805 5557 65861
rect 5613 65805 5699 65861
rect 5755 65805 5841 65861
rect 5897 65805 5983 65861
rect 6039 65805 6125 65861
rect 6181 65805 6267 65861
rect 6323 65805 6409 65861
rect 6465 65805 6551 65861
rect 6607 65805 6693 65861
rect 6749 65805 6835 65861
rect 6891 65805 6977 65861
rect 7033 65805 7119 65861
rect 7175 65805 7261 65861
rect 7317 65805 7403 65861
rect 7459 65805 7545 65861
rect 7601 65805 7687 65861
rect 7743 65805 7829 65861
rect 7885 65805 7971 65861
rect 8027 65805 8113 65861
rect 8169 65805 8255 65861
rect 8311 65805 8397 65861
rect 8453 65805 8539 65861
rect 8595 65805 8681 65861
rect 8737 65805 8823 65861
rect 8879 65805 8965 65861
rect 9021 65805 9107 65861
rect 9163 65805 9249 65861
rect 9305 65805 9391 65861
rect 9447 65805 9533 65861
rect 9589 65805 9675 65861
rect 9731 65805 9817 65861
rect 9873 65805 9959 65861
rect 10015 65805 10101 65861
rect 10157 65805 10243 65861
rect 10299 65805 10385 65861
rect 10441 65805 10527 65861
rect 10583 65805 10669 65861
rect 10725 65805 10811 65861
rect 10867 65805 10953 65861
rect 11009 65805 11095 65861
rect 11151 65805 11237 65861
rect 11293 65805 11379 65861
rect 11435 65805 11521 65861
rect 11577 65805 11663 65861
rect 11719 65805 11805 65861
rect 11861 65805 11947 65861
rect 12003 65805 12089 65861
rect 12145 65805 12231 65861
rect 12287 65805 12373 65861
rect 12429 65805 12515 65861
rect 12571 65805 12657 65861
rect 12713 65805 12799 65861
rect 12855 65805 12941 65861
rect 12997 65805 13083 65861
rect 13139 65805 13225 65861
rect 13281 65805 13367 65861
rect 13423 65805 13509 65861
rect 13565 65805 13651 65861
rect 13707 65805 13793 65861
rect 13849 65805 13935 65861
rect 13991 65805 14077 65861
rect 14133 65805 14219 65861
rect 14275 65805 14361 65861
rect 14417 65805 14503 65861
rect 14559 65805 14645 65861
rect 14701 65805 14787 65861
rect 14843 65805 15000 65861
rect 0 65719 15000 65805
rect 0 65663 161 65719
rect 217 65663 303 65719
rect 359 65663 445 65719
rect 501 65663 587 65719
rect 643 65663 729 65719
rect 785 65663 871 65719
rect 927 65663 1013 65719
rect 1069 65663 1155 65719
rect 1211 65663 1297 65719
rect 1353 65663 1439 65719
rect 1495 65663 1581 65719
rect 1637 65663 1723 65719
rect 1779 65663 1865 65719
rect 1921 65663 2007 65719
rect 2063 65663 2149 65719
rect 2205 65663 2291 65719
rect 2347 65663 2433 65719
rect 2489 65663 2575 65719
rect 2631 65663 2717 65719
rect 2773 65663 2859 65719
rect 2915 65663 3001 65719
rect 3057 65663 3143 65719
rect 3199 65663 3285 65719
rect 3341 65663 3427 65719
rect 3483 65663 3569 65719
rect 3625 65663 3711 65719
rect 3767 65663 3853 65719
rect 3909 65663 3995 65719
rect 4051 65663 4137 65719
rect 4193 65663 4279 65719
rect 4335 65663 4421 65719
rect 4477 65663 4563 65719
rect 4619 65663 4705 65719
rect 4761 65663 4847 65719
rect 4903 65663 4989 65719
rect 5045 65663 5131 65719
rect 5187 65663 5273 65719
rect 5329 65663 5415 65719
rect 5471 65663 5557 65719
rect 5613 65663 5699 65719
rect 5755 65663 5841 65719
rect 5897 65663 5983 65719
rect 6039 65663 6125 65719
rect 6181 65663 6267 65719
rect 6323 65663 6409 65719
rect 6465 65663 6551 65719
rect 6607 65663 6693 65719
rect 6749 65663 6835 65719
rect 6891 65663 6977 65719
rect 7033 65663 7119 65719
rect 7175 65663 7261 65719
rect 7317 65663 7403 65719
rect 7459 65663 7545 65719
rect 7601 65663 7687 65719
rect 7743 65663 7829 65719
rect 7885 65663 7971 65719
rect 8027 65663 8113 65719
rect 8169 65663 8255 65719
rect 8311 65663 8397 65719
rect 8453 65663 8539 65719
rect 8595 65663 8681 65719
rect 8737 65663 8823 65719
rect 8879 65663 8965 65719
rect 9021 65663 9107 65719
rect 9163 65663 9249 65719
rect 9305 65663 9391 65719
rect 9447 65663 9533 65719
rect 9589 65663 9675 65719
rect 9731 65663 9817 65719
rect 9873 65663 9959 65719
rect 10015 65663 10101 65719
rect 10157 65663 10243 65719
rect 10299 65663 10385 65719
rect 10441 65663 10527 65719
rect 10583 65663 10669 65719
rect 10725 65663 10811 65719
rect 10867 65663 10953 65719
rect 11009 65663 11095 65719
rect 11151 65663 11237 65719
rect 11293 65663 11379 65719
rect 11435 65663 11521 65719
rect 11577 65663 11663 65719
rect 11719 65663 11805 65719
rect 11861 65663 11947 65719
rect 12003 65663 12089 65719
rect 12145 65663 12231 65719
rect 12287 65663 12373 65719
rect 12429 65663 12515 65719
rect 12571 65663 12657 65719
rect 12713 65663 12799 65719
rect 12855 65663 12941 65719
rect 12997 65663 13083 65719
rect 13139 65663 13225 65719
rect 13281 65663 13367 65719
rect 13423 65663 13509 65719
rect 13565 65663 13651 65719
rect 13707 65663 13793 65719
rect 13849 65663 13935 65719
rect 13991 65663 14077 65719
rect 14133 65663 14219 65719
rect 14275 65663 14361 65719
rect 14417 65663 14503 65719
rect 14559 65663 14645 65719
rect 14701 65663 14787 65719
rect 14843 65663 15000 65719
rect 0 65577 15000 65663
rect 0 65521 161 65577
rect 217 65521 303 65577
rect 359 65521 445 65577
rect 501 65521 587 65577
rect 643 65521 729 65577
rect 785 65521 871 65577
rect 927 65521 1013 65577
rect 1069 65521 1155 65577
rect 1211 65521 1297 65577
rect 1353 65521 1439 65577
rect 1495 65521 1581 65577
rect 1637 65521 1723 65577
rect 1779 65521 1865 65577
rect 1921 65521 2007 65577
rect 2063 65521 2149 65577
rect 2205 65521 2291 65577
rect 2347 65521 2433 65577
rect 2489 65521 2575 65577
rect 2631 65521 2717 65577
rect 2773 65521 2859 65577
rect 2915 65521 3001 65577
rect 3057 65521 3143 65577
rect 3199 65521 3285 65577
rect 3341 65521 3427 65577
rect 3483 65521 3569 65577
rect 3625 65521 3711 65577
rect 3767 65521 3853 65577
rect 3909 65521 3995 65577
rect 4051 65521 4137 65577
rect 4193 65521 4279 65577
rect 4335 65521 4421 65577
rect 4477 65521 4563 65577
rect 4619 65521 4705 65577
rect 4761 65521 4847 65577
rect 4903 65521 4989 65577
rect 5045 65521 5131 65577
rect 5187 65521 5273 65577
rect 5329 65521 5415 65577
rect 5471 65521 5557 65577
rect 5613 65521 5699 65577
rect 5755 65521 5841 65577
rect 5897 65521 5983 65577
rect 6039 65521 6125 65577
rect 6181 65521 6267 65577
rect 6323 65521 6409 65577
rect 6465 65521 6551 65577
rect 6607 65521 6693 65577
rect 6749 65521 6835 65577
rect 6891 65521 6977 65577
rect 7033 65521 7119 65577
rect 7175 65521 7261 65577
rect 7317 65521 7403 65577
rect 7459 65521 7545 65577
rect 7601 65521 7687 65577
rect 7743 65521 7829 65577
rect 7885 65521 7971 65577
rect 8027 65521 8113 65577
rect 8169 65521 8255 65577
rect 8311 65521 8397 65577
rect 8453 65521 8539 65577
rect 8595 65521 8681 65577
rect 8737 65521 8823 65577
rect 8879 65521 8965 65577
rect 9021 65521 9107 65577
rect 9163 65521 9249 65577
rect 9305 65521 9391 65577
rect 9447 65521 9533 65577
rect 9589 65521 9675 65577
rect 9731 65521 9817 65577
rect 9873 65521 9959 65577
rect 10015 65521 10101 65577
rect 10157 65521 10243 65577
rect 10299 65521 10385 65577
rect 10441 65521 10527 65577
rect 10583 65521 10669 65577
rect 10725 65521 10811 65577
rect 10867 65521 10953 65577
rect 11009 65521 11095 65577
rect 11151 65521 11237 65577
rect 11293 65521 11379 65577
rect 11435 65521 11521 65577
rect 11577 65521 11663 65577
rect 11719 65521 11805 65577
rect 11861 65521 11947 65577
rect 12003 65521 12089 65577
rect 12145 65521 12231 65577
rect 12287 65521 12373 65577
rect 12429 65521 12515 65577
rect 12571 65521 12657 65577
rect 12713 65521 12799 65577
rect 12855 65521 12941 65577
rect 12997 65521 13083 65577
rect 13139 65521 13225 65577
rect 13281 65521 13367 65577
rect 13423 65521 13509 65577
rect 13565 65521 13651 65577
rect 13707 65521 13793 65577
rect 13849 65521 13935 65577
rect 13991 65521 14077 65577
rect 14133 65521 14219 65577
rect 14275 65521 14361 65577
rect 14417 65521 14503 65577
rect 14559 65521 14645 65577
rect 14701 65521 14787 65577
rect 14843 65521 15000 65577
rect 0 65435 15000 65521
rect 0 65379 161 65435
rect 217 65379 303 65435
rect 359 65379 445 65435
rect 501 65379 587 65435
rect 643 65379 729 65435
rect 785 65379 871 65435
rect 927 65379 1013 65435
rect 1069 65379 1155 65435
rect 1211 65379 1297 65435
rect 1353 65379 1439 65435
rect 1495 65379 1581 65435
rect 1637 65379 1723 65435
rect 1779 65379 1865 65435
rect 1921 65379 2007 65435
rect 2063 65379 2149 65435
rect 2205 65379 2291 65435
rect 2347 65379 2433 65435
rect 2489 65379 2575 65435
rect 2631 65379 2717 65435
rect 2773 65379 2859 65435
rect 2915 65379 3001 65435
rect 3057 65379 3143 65435
rect 3199 65379 3285 65435
rect 3341 65379 3427 65435
rect 3483 65379 3569 65435
rect 3625 65379 3711 65435
rect 3767 65379 3853 65435
rect 3909 65379 3995 65435
rect 4051 65379 4137 65435
rect 4193 65379 4279 65435
rect 4335 65379 4421 65435
rect 4477 65379 4563 65435
rect 4619 65379 4705 65435
rect 4761 65379 4847 65435
rect 4903 65379 4989 65435
rect 5045 65379 5131 65435
rect 5187 65379 5273 65435
rect 5329 65379 5415 65435
rect 5471 65379 5557 65435
rect 5613 65379 5699 65435
rect 5755 65379 5841 65435
rect 5897 65379 5983 65435
rect 6039 65379 6125 65435
rect 6181 65379 6267 65435
rect 6323 65379 6409 65435
rect 6465 65379 6551 65435
rect 6607 65379 6693 65435
rect 6749 65379 6835 65435
rect 6891 65379 6977 65435
rect 7033 65379 7119 65435
rect 7175 65379 7261 65435
rect 7317 65379 7403 65435
rect 7459 65379 7545 65435
rect 7601 65379 7687 65435
rect 7743 65379 7829 65435
rect 7885 65379 7971 65435
rect 8027 65379 8113 65435
rect 8169 65379 8255 65435
rect 8311 65379 8397 65435
rect 8453 65379 8539 65435
rect 8595 65379 8681 65435
rect 8737 65379 8823 65435
rect 8879 65379 8965 65435
rect 9021 65379 9107 65435
rect 9163 65379 9249 65435
rect 9305 65379 9391 65435
rect 9447 65379 9533 65435
rect 9589 65379 9675 65435
rect 9731 65379 9817 65435
rect 9873 65379 9959 65435
rect 10015 65379 10101 65435
rect 10157 65379 10243 65435
rect 10299 65379 10385 65435
rect 10441 65379 10527 65435
rect 10583 65379 10669 65435
rect 10725 65379 10811 65435
rect 10867 65379 10953 65435
rect 11009 65379 11095 65435
rect 11151 65379 11237 65435
rect 11293 65379 11379 65435
rect 11435 65379 11521 65435
rect 11577 65379 11663 65435
rect 11719 65379 11805 65435
rect 11861 65379 11947 65435
rect 12003 65379 12089 65435
rect 12145 65379 12231 65435
rect 12287 65379 12373 65435
rect 12429 65379 12515 65435
rect 12571 65379 12657 65435
rect 12713 65379 12799 65435
rect 12855 65379 12941 65435
rect 12997 65379 13083 65435
rect 13139 65379 13225 65435
rect 13281 65379 13367 65435
rect 13423 65379 13509 65435
rect 13565 65379 13651 65435
rect 13707 65379 13793 65435
rect 13849 65379 13935 65435
rect 13991 65379 14077 65435
rect 14133 65379 14219 65435
rect 14275 65379 14361 65435
rect 14417 65379 14503 65435
rect 14559 65379 14645 65435
rect 14701 65379 14787 65435
rect 14843 65379 15000 65435
rect 0 65293 15000 65379
rect 0 65237 161 65293
rect 217 65237 303 65293
rect 359 65237 445 65293
rect 501 65237 587 65293
rect 643 65237 729 65293
rect 785 65237 871 65293
rect 927 65237 1013 65293
rect 1069 65237 1155 65293
rect 1211 65237 1297 65293
rect 1353 65237 1439 65293
rect 1495 65237 1581 65293
rect 1637 65237 1723 65293
rect 1779 65237 1865 65293
rect 1921 65237 2007 65293
rect 2063 65237 2149 65293
rect 2205 65237 2291 65293
rect 2347 65237 2433 65293
rect 2489 65237 2575 65293
rect 2631 65237 2717 65293
rect 2773 65237 2859 65293
rect 2915 65237 3001 65293
rect 3057 65237 3143 65293
rect 3199 65237 3285 65293
rect 3341 65237 3427 65293
rect 3483 65237 3569 65293
rect 3625 65237 3711 65293
rect 3767 65237 3853 65293
rect 3909 65237 3995 65293
rect 4051 65237 4137 65293
rect 4193 65237 4279 65293
rect 4335 65237 4421 65293
rect 4477 65237 4563 65293
rect 4619 65237 4705 65293
rect 4761 65237 4847 65293
rect 4903 65237 4989 65293
rect 5045 65237 5131 65293
rect 5187 65237 5273 65293
rect 5329 65237 5415 65293
rect 5471 65237 5557 65293
rect 5613 65237 5699 65293
rect 5755 65237 5841 65293
rect 5897 65237 5983 65293
rect 6039 65237 6125 65293
rect 6181 65237 6267 65293
rect 6323 65237 6409 65293
rect 6465 65237 6551 65293
rect 6607 65237 6693 65293
rect 6749 65237 6835 65293
rect 6891 65237 6977 65293
rect 7033 65237 7119 65293
rect 7175 65237 7261 65293
rect 7317 65237 7403 65293
rect 7459 65237 7545 65293
rect 7601 65237 7687 65293
rect 7743 65237 7829 65293
rect 7885 65237 7971 65293
rect 8027 65237 8113 65293
rect 8169 65237 8255 65293
rect 8311 65237 8397 65293
rect 8453 65237 8539 65293
rect 8595 65237 8681 65293
rect 8737 65237 8823 65293
rect 8879 65237 8965 65293
rect 9021 65237 9107 65293
rect 9163 65237 9249 65293
rect 9305 65237 9391 65293
rect 9447 65237 9533 65293
rect 9589 65237 9675 65293
rect 9731 65237 9817 65293
rect 9873 65237 9959 65293
rect 10015 65237 10101 65293
rect 10157 65237 10243 65293
rect 10299 65237 10385 65293
rect 10441 65237 10527 65293
rect 10583 65237 10669 65293
rect 10725 65237 10811 65293
rect 10867 65237 10953 65293
rect 11009 65237 11095 65293
rect 11151 65237 11237 65293
rect 11293 65237 11379 65293
rect 11435 65237 11521 65293
rect 11577 65237 11663 65293
rect 11719 65237 11805 65293
rect 11861 65237 11947 65293
rect 12003 65237 12089 65293
rect 12145 65237 12231 65293
rect 12287 65237 12373 65293
rect 12429 65237 12515 65293
rect 12571 65237 12657 65293
rect 12713 65237 12799 65293
rect 12855 65237 12941 65293
rect 12997 65237 13083 65293
rect 13139 65237 13225 65293
rect 13281 65237 13367 65293
rect 13423 65237 13509 65293
rect 13565 65237 13651 65293
rect 13707 65237 13793 65293
rect 13849 65237 13935 65293
rect 13991 65237 14077 65293
rect 14133 65237 14219 65293
rect 14275 65237 14361 65293
rect 14417 65237 14503 65293
rect 14559 65237 14645 65293
rect 14701 65237 14787 65293
rect 14843 65237 15000 65293
rect 0 65200 15000 65237
rect 0 64963 15000 65000
rect 0 64907 161 64963
rect 217 64907 303 64963
rect 359 64907 445 64963
rect 501 64907 587 64963
rect 643 64907 729 64963
rect 785 64907 871 64963
rect 927 64907 1013 64963
rect 1069 64907 1155 64963
rect 1211 64907 1297 64963
rect 1353 64907 1439 64963
rect 1495 64907 1581 64963
rect 1637 64907 1723 64963
rect 1779 64907 1865 64963
rect 1921 64907 2007 64963
rect 2063 64907 2149 64963
rect 2205 64907 2291 64963
rect 2347 64907 2433 64963
rect 2489 64907 2575 64963
rect 2631 64907 2717 64963
rect 2773 64907 2859 64963
rect 2915 64907 3001 64963
rect 3057 64907 3143 64963
rect 3199 64907 3285 64963
rect 3341 64907 3427 64963
rect 3483 64907 3569 64963
rect 3625 64907 3711 64963
rect 3767 64907 3853 64963
rect 3909 64907 3995 64963
rect 4051 64907 4137 64963
rect 4193 64907 4279 64963
rect 4335 64907 4421 64963
rect 4477 64907 4563 64963
rect 4619 64907 4705 64963
rect 4761 64907 4847 64963
rect 4903 64907 4989 64963
rect 5045 64907 5131 64963
rect 5187 64907 5273 64963
rect 5329 64907 5415 64963
rect 5471 64907 5557 64963
rect 5613 64907 5699 64963
rect 5755 64907 5841 64963
rect 5897 64907 5983 64963
rect 6039 64907 6125 64963
rect 6181 64907 6267 64963
rect 6323 64907 6409 64963
rect 6465 64907 6551 64963
rect 6607 64907 6693 64963
rect 6749 64907 6835 64963
rect 6891 64907 6977 64963
rect 7033 64907 7119 64963
rect 7175 64907 7261 64963
rect 7317 64907 7403 64963
rect 7459 64907 7545 64963
rect 7601 64907 7687 64963
rect 7743 64907 7829 64963
rect 7885 64907 7971 64963
rect 8027 64907 8113 64963
rect 8169 64907 8255 64963
rect 8311 64907 8397 64963
rect 8453 64907 8539 64963
rect 8595 64907 8681 64963
rect 8737 64907 8823 64963
rect 8879 64907 8965 64963
rect 9021 64907 9107 64963
rect 9163 64907 9249 64963
rect 9305 64907 9391 64963
rect 9447 64907 9533 64963
rect 9589 64907 9675 64963
rect 9731 64907 9817 64963
rect 9873 64907 9959 64963
rect 10015 64907 10101 64963
rect 10157 64907 10243 64963
rect 10299 64907 10385 64963
rect 10441 64907 10527 64963
rect 10583 64907 10669 64963
rect 10725 64907 10811 64963
rect 10867 64907 10953 64963
rect 11009 64907 11095 64963
rect 11151 64907 11237 64963
rect 11293 64907 11379 64963
rect 11435 64907 11521 64963
rect 11577 64907 11663 64963
rect 11719 64907 11805 64963
rect 11861 64907 11947 64963
rect 12003 64907 12089 64963
rect 12145 64907 12231 64963
rect 12287 64907 12373 64963
rect 12429 64907 12515 64963
rect 12571 64907 12657 64963
rect 12713 64907 12799 64963
rect 12855 64907 12941 64963
rect 12997 64907 13083 64963
rect 13139 64907 13225 64963
rect 13281 64907 13367 64963
rect 13423 64907 13509 64963
rect 13565 64907 13651 64963
rect 13707 64907 13793 64963
rect 13849 64907 13935 64963
rect 13991 64907 14077 64963
rect 14133 64907 14219 64963
rect 14275 64907 14361 64963
rect 14417 64907 14503 64963
rect 14559 64907 14645 64963
rect 14701 64907 14787 64963
rect 14843 64907 15000 64963
rect 0 64821 15000 64907
rect 0 64765 161 64821
rect 217 64765 303 64821
rect 359 64765 445 64821
rect 501 64765 587 64821
rect 643 64765 729 64821
rect 785 64765 871 64821
rect 927 64765 1013 64821
rect 1069 64765 1155 64821
rect 1211 64765 1297 64821
rect 1353 64765 1439 64821
rect 1495 64765 1581 64821
rect 1637 64765 1723 64821
rect 1779 64765 1865 64821
rect 1921 64765 2007 64821
rect 2063 64765 2149 64821
rect 2205 64765 2291 64821
rect 2347 64765 2433 64821
rect 2489 64765 2575 64821
rect 2631 64765 2717 64821
rect 2773 64765 2859 64821
rect 2915 64765 3001 64821
rect 3057 64765 3143 64821
rect 3199 64765 3285 64821
rect 3341 64765 3427 64821
rect 3483 64765 3569 64821
rect 3625 64765 3711 64821
rect 3767 64765 3853 64821
rect 3909 64765 3995 64821
rect 4051 64765 4137 64821
rect 4193 64765 4279 64821
rect 4335 64765 4421 64821
rect 4477 64765 4563 64821
rect 4619 64765 4705 64821
rect 4761 64765 4847 64821
rect 4903 64765 4989 64821
rect 5045 64765 5131 64821
rect 5187 64765 5273 64821
rect 5329 64765 5415 64821
rect 5471 64765 5557 64821
rect 5613 64765 5699 64821
rect 5755 64765 5841 64821
rect 5897 64765 5983 64821
rect 6039 64765 6125 64821
rect 6181 64765 6267 64821
rect 6323 64765 6409 64821
rect 6465 64765 6551 64821
rect 6607 64765 6693 64821
rect 6749 64765 6835 64821
rect 6891 64765 6977 64821
rect 7033 64765 7119 64821
rect 7175 64765 7261 64821
rect 7317 64765 7403 64821
rect 7459 64765 7545 64821
rect 7601 64765 7687 64821
rect 7743 64765 7829 64821
rect 7885 64765 7971 64821
rect 8027 64765 8113 64821
rect 8169 64765 8255 64821
rect 8311 64765 8397 64821
rect 8453 64765 8539 64821
rect 8595 64765 8681 64821
rect 8737 64765 8823 64821
rect 8879 64765 8965 64821
rect 9021 64765 9107 64821
rect 9163 64765 9249 64821
rect 9305 64765 9391 64821
rect 9447 64765 9533 64821
rect 9589 64765 9675 64821
rect 9731 64765 9817 64821
rect 9873 64765 9959 64821
rect 10015 64765 10101 64821
rect 10157 64765 10243 64821
rect 10299 64765 10385 64821
rect 10441 64765 10527 64821
rect 10583 64765 10669 64821
rect 10725 64765 10811 64821
rect 10867 64765 10953 64821
rect 11009 64765 11095 64821
rect 11151 64765 11237 64821
rect 11293 64765 11379 64821
rect 11435 64765 11521 64821
rect 11577 64765 11663 64821
rect 11719 64765 11805 64821
rect 11861 64765 11947 64821
rect 12003 64765 12089 64821
rect 12145 64765 12231 64821
rect 12287 64765 12373 64821
rect 12429 64765 12515 64821
rect 12571 64765 12657 64821
rect 12713 64765 12799 64821
rect 12855 64765 12941 64821
rect 12997 64765 13083 64821
rect 13139 64765 13225 64821
rect 13281 64765 13367 64821
rect 13423 64765 13509 64821
rect 13565 64765 13651 64821
rect 13707 64765 13793 64821
rect 13849 64765 13935 64821
rect 13991 64765 14077 64821
rect 14133 64765 14219 64821
rect 14275 64765 14361 64821
rect 14417 64765 14503 64821
rect 14559 64765 14645 64821
rect 14701 64765 14787 64821
rect 14843 64765 15000 64821
rect 0 64679 15000 64765
rect 0 64623 161 64679
rect 217 64623 303 64679
rect 359 64623 445 64679
rect 501 64623 587 64679
rect 643 64623 729 64679
rect 785 64623 871 64679
rect 927 64623 1013 64679
rect 1069 64623 1155 64679
rect 1211 64623 1297 64679
rect 1353 64623 1439 64679
rect 1495 64623 1581 64679
rect 1637 64623 1723 64679
rect 1779 64623 1865 64679
rect 1921 64623 2007 64679
rect 2063 64623 2149 64679
rect 2205 64623 2291 64679
rect 2347 64623 2433 64679
rect 2489 64623 2575 64679
rect 2631 64623 2717 64679
rect 2773 64623 2859 64679
rect 2915 64623 3001 64679
rect 3057 64623 3143 64679
rect 3199 64623 3285 64679
rect 3341 64623 3427 64679
rect 3483 64623 3569 64679
rect 3625 64623 3711 64679
rect 3767 64623 3853 64679
rect 3909 64623 3995 64679
rect 4051 64623 4137 64679
rect 4193 64623 4279 64679
rect 4335 64623 4421 64679
rect 4477 64623 4563 64679
rect 4619 64623 4705 64679
rect 4761 64623 4847 64679
rect 4903 64623 4989 64679
rect 5045 64623 5131 64679
rect 5187 64623 5273 64679
rect 5329 64623 5415 64679
rect 5471 64623 5557 64679
rect 5613 64623 5699 64679
rect 5755 64623 5841 64679
rect 5897 64623 5983 64679
rect 6039 64623 6125 64679
rect 6181 64623 6267 64679
rect 6323 64623 6409 64679
rect 6465 64623 6551 64679
rect 6607 64623 6693 64679
rect 6749 64623 6835 64679
rect 6891 64623 6977 64679
rect 7033 64623 7119 64679
rect 7175 64623 7261 64679
rect 7317 64623 7403 64679
rect 7459 64623 7545 64679
rect 7601 64623 7687 64679
rect 7743 64623 7829 64679
rect 7885 64623 7971 64679
rect 8027 64623 8113 64679
rect 8169 64623 8255 64679
rect 8311 64623 8397 64679
rect 8453 64623 8539 64679
rect 8595 64623 8681 64679
rect 8737 64623 8823 64679
rect 8879 64623 8965 64679
rect 9021 64623 9107 64679
rect 9163 64623 9249 64679
rect 9305 64623 9391 64679
rect 9447 64623 9533 64679
rect 9589 64623 9675 64679
rect 9731 64623 9817 64679
rect 9873 64623 9959 64679
rect 10015 64623 10101 64679
rect 10157 64623 10243 64679
rect 10299 64623 10385 64679
rect 10441 64623 10527 64679
rect 10583 64623 10669 64679
rect 10725 64623 10811 64679
rect 10867 64623 10953 64679
rect 11009 64623 11095 64679
rect 11151 64623 11237 64679
rect 11293 64623 11379 64679
rect 11435 64623 11521 64679
rect 11577 64623 11663 64679
rect 11719 64623 11805 64679
rect 11861 64623 11947 64679
rect 12003 64623 12089 64679
rect 12145 64623 12231 64679
rect 12287 64623 12373 64679
rect 12429 64623 12515 64679
rect 12571 64623 12657 64679
rect 12713 64623 12799 64679
rect 12855 64623 12941 64679
rect 12997 64623 13083 64679
rect 13139 64623 13225 64679
rect 13281 64623 13367 64679
rect 13423 64623 13509 64679
rect 13565 64623 13651 64679
rect 13707 64623 13793 64679
rect 13849 64623 13935 64679
rect 13991 64623 14077 64679
rect 14133 64623 14219 64679
rect 14275 64623 14361 64679
rect 14417 64623 14503 64679
rect 14559 64623 14645 64679
rect 14701 64623 14787 64679
rect 14843 64623 15000 64679
rect 0 64537 15000 64623
rect 0 64481 161 64537
rect 217 64481 303 64537
rect 359 64481 445 64537
rect 501 64481 587 64537
rect 643 64481 729 64537
rect 785 64481 871 64537
rect 927 64481 1013 64537
rect 1069 64481 1155 64537
rect 1211 64481 1297 64537
rect 1353 64481 1439 64537
rect 1495 64481 1581 64537
rect 1637 64481 1723 64537
rect 1779 64481 1865 64537
rect 1921 64481 2007 64537
rect 2063 64481 2149 64537
rect 2205 64481 2291 64537
rect 2347 64481 2433 64537
rect 2489 64481 2575 64537
rect 2631 64481 2717 64537
rect 2773 64481 2859 64537
rect 2915 64481 3001 64537
rect 3057 64481 3143 64537
rect 3199 64481 3285 64537
rect 3341 64481 3427 64537
rect 3483 64481 3569 64537
rect 3625 64481 3711 64537
rect 3767 64481 3853 64537
rect 3909 64481 3995 64537
rect 4051 64481 4137 64537
rect 4193 64481 4279 64537
rect 4335 64481 4421 64537
rect 4477 64481 4563 64537
rect 4619 64481 4705 64537
rect 4761 64481 4847 64537
rect 4903 64481 4989 64537
rect 5045 64481 5131 64537
rect 5187 64481 5273 64537
rect 5329 64481 5415 64537
rect 5471 64481 5557 64537
rect 5613 64481 5699 64537
rect 5755 64481 5841 64537
rect 5897 64481 5983 64537
rect 6039 64481 6125 64537
rect 6181 64481 6267 64537
rect 6323 64481 6409 64537
rect 6465 64481 6551 64537
rect 6607 64481 6693 64537
rect 6749 64481 6835 64537
rect 6891 64481 6977 64537
rect 7033 64481 7119 64537
rect 7175 64481 7261 64537
rect 7317 64481 7403 64537
rect 7459 64481 7545 64537
rect 7601 64481 7687 64537
rect 7743 64481 7829 64537
rect 7885 64481 7971 64537
rect 8027 64481 8113 64537
rect 8169 64481 8255 64537
rect 8311 64481 8397 64537
rect 8453 64481 8539 64537
rect 8595 64481 8681 64537
rect 8737 64481 8823 64537
rect 8879 64481 8965 64537
rect 9021 64481 9107 64537
rect 9163 64481 9249 64537
rect 9305 64481 9391 64537
rect 9447 64481 9533 64537
rect 9589 64481 9675 64537
rect 9731 64481 9817 64537
rect 9873 64481 9959 64537
rect 10015 64481 10101 64537
rect 10157 64481 10243 64537
rect 10299 64481 10385 64537
rect 10441 64481 10527 64537
rect 10583 64481 10669 64537
rect 10725 64481 10811 64537
rect 10867 64481 10953 64537
rect 11009 64481 11095 64537
rect 11151 64481 11237 64537
rect 11293 64481 11379 64537
rect 11435 64481 11521 64537
rect 11577 64481 11663 64537
rect 11719 64481 11805 64537
rect 11861 64481 11947 64537
rect 12003 64481 12089 64537
rect 12145 64481 12231 64537
rect 12287 64481 12373 64537
rect 12429 64481 12515 64537
rect 12571 64481 12657 64537
rect 12713 64481 12799 64537
rect 12855 64481 12941 64537
rect 12997 64481 13083 64537
rect 13139 64481 13225 64537
rect 13281 64481 13367 64537
rect 13423 64481 13509 64537
rect 13565 64481 13651 64537
rect 13707 64481 13793 64537
rect 13849 64481 13935 64537
rect 13991 64481 14077 64537
rect 14133 64481 14219 64537
rect 14275 64481 14361 64537
rect 14417 64481 14503 64537
rect 14559 64481 14645 64537
rect 14701 64481 14787 64537
rect 14843 64481 15000 64537
rect 0 64395 15000 64481
rect 0 64339 161 64395
rect 217 64339 303 64395
rect 359 64339 445 64395
rect 501 64339 587 64395
rect 643 64339 729 64395
rect 785 64339 871 64395
rect 927 64339 1013 64395
rect 1069 64339 1155 64395
rect 1211 64339 1297 64395
rect 1353 64339 1439 64395
rect 1495 64339 1581 64395
rect 1637 64339 1723 64395
rect 1779 64339 1865 64395
rect 1921 64339 2007 64395
rect 2063 64339 2149 64395
rect 2205 64339 2291 64395
rect 2347 64339 2433 64395
rect 2489 64339 2575 64395
rect 2631 64339 2717 64395
rect 2773 64339 2859 64395
rect 2915 64339 3001 64395
rect 3057 64339 3143 64395
rect 3199 64339 3285 64395
rect 3341 64339 3427 64395
rect 3483 64339 3569 64395
rect 3625 64339 3711 64395
rect 3767 64339 3853 64395
rect 3909 64339 3995 64395
rect 4051 64339 4137 64395
rect 4193 64339 4279 64395
rect 4335 64339 4421 64395
rect 4477 64339 4563 64395
rect 4619 64339 4705 64395
rect 4761 64339 4847 64395
rect 4903 64339 4989 64395
rect 5045 64339 5131 64395
rect 5187 64339 5273 64395
rect 5329 64339 5415 64395
rect 5471 64339 5557 64395
rect 5613 64339 5699 64395
rect 5755 64339 5841 64395
rect 5897 64339 5983 64395
rect 6039 64339 6125 64395
rect 6181 64339 6267 64395
rect 6323 64339 6409 64395
rect 6465 64339 6551 64395
rect 6607 64339 6693 64395
rect 6749 64339 6835 64395
rect 6891 64339 6977 64395
rect 7033 64339 7119 64395
rect 7175 64339 7261 64395
rect 7317 64339 7403 64395
rect 7459 64339 7545 64395
rect 7601 64339 7687 64395
rect 7743 64339 7829 64395
rect 7885 64339 7971 64395
rect 8027 64339 8113 64395
rect 8169 64339 8255 64395
rect 8311 64339 8397 64395
rect 8453 64339 8539 64395
rect 8595 64339 8681 64395
rect 8737 64339 8823 64395
rect 8879 64339 8965 64395
rect 9021 64339 9107 64395
rect 9163 64339 9249 64395
rect 9305 64339 9391 64395
rect 9447 64339 9533 64395
rect 9589 64339 9675 64395
rect 9731 64339 9817 64395
rect 9873 64339 9959 64395
rect 10015 64339 10101 64395
rect 10157 64339 10243 64395
rect 10299 64339 10385 64395
rect 10441 64339 10527 64395
rect 10583 64339 10669 64395
rect 10725 64339 10811 64395
rect 10867 64339 10953 64395
rect 11009 64339 11095 64395
rect 11151 64339 11237 64395
rect 11293 64339 11379 64395
rect 11435 64339 11521 64395
rect 11577 64339 11663 64395
rect 11719 64339 11805 64395
rect 11861 64339 11947 64395
rect 12003 64339 12089 64395
rect 12145 64339 12231 64395
rect 12287 64339 12373 64395
rect 12429 64339 12515 64395
rect 12571 64339 12657 64395
rect 12713 64339 12799 64395
rect 12855 64339 12941 64395
rect 12997 64339 13083 64395
rect 13139 64339 13225 64395
rect 13281 64339 13367 64395
rect 13423 64339 13509 64395
rect 13565 64339 13651 64395
rect 13707 64339 13793 64395
rect 13849 64339 13935 64395
rect 13991 64339 14077 64395
rect 14133 64339 14219 64395
rect 14275 64339 14361 64395
rect 14417 64339 14503 64395
rect 14559 64339 14645 64395
rect 14701 64339 14787 64395
rect 14843 64339 15000 64395
rect 0 64253 15000 64339
rect 0 64197 161 64253
rect 217 64197 303 64253
rect 359 64197 445 64253
rect 501 64197 587 64253
rect 643 64197 729 64253
rect 785 64197 871 64253
rect 927 64197 1013 64253
rect 1069 64197 1155 64253
rect 1211 64197 1297 64253
rect 1353 64197 1439 64253
rect 1495 64197 1581 64253
rect 1637 64197 1723 64253
rect 1779 64197 1865 64253
rect 1921 64197 2007 64253
rect 2063 64197 2149 64253
rect 2205 64197 2291 64253
rect 2347 64197 2433 64253
rect 2489 64197 2575 64253
rect 2631 64197 2717 64253
rect 2773 64197 2859 64253
rect 2915 64197 3001 64253
rect 3057 64197 3143 64253
rect 3199 64197 3285 64253
rect 3341 64197 3427 64253
rect 3483 64197 3569 64253
rect 3625 64197 3711 64253
rect 3767 64197 3853 64253
rect 3909 64197 3995 64253
rect 4051 64197 4137 64253
rect 4193 64197 4279 64253
rect 4335 64197 4421 64253
rect 4477 64197 4563 64253
rect 4619 64197 4705 64253
rect 4761 64197 4847 64253
rect 4903 64197 4989 64253
rect 5045 64197 5131 64253
rect 5187 64197 5273 64253
rect 5329 64197 5415 64253
rect 5471 64197 5557 64253
rect 5613 64197 5699 64253
rect 5755 64197 5841 64253
rect 5897 64197 5983 64253
rect 6039 64197 6125 64253
rect 6181 64197 6267 64253
rect 6323 64197 6409 64253
rect 6465 64197 6551 64253
rect 6607 64197 6693 64253
rect 6749 64197 6835 64253
rect 6891 64197 6977 64253
rect 7033 64197 7119 64253
rect 7175 64197 7261 64253
rect 7317 64197 7403 64253
rect 7459 64197 7545 64253
rect 7601 64197 7687 64253
rect 7743 64197 7829 64253
rect 7885 64197 7971 64253
rect 8027 64197 8113 64253
rect 8169 64197 8255 64253
rect 8311 64197 8397 64253
rect 8453 64197 8539 64253
rect 8595 64197 8681 64253
rect 8737 64197 8823 64253
rect 8879 64197 8965 64253
rect 9021 64197 9107 64253
rect 9163 64197 9249 64253
rect 9305 64197 9391 64253
rect 9447 64197 9533 64253
rect 9589 64197 9675 64253
rect 9731 64197 9817 64253
rect 9873 64197 9959 64253
rect 10015 64197 10101 64253
rect 10157 64197 10243 64253
rect 10299 64197 10385 64253
rect 10441 64197 10527 64253
rect 10583 64197 10669 64253
rect 10725 64197 10811 64253
rect 10867 64197 10953 64253
rect 11009 64197 11095 64253
rect 11151 64197 11237 64253
rect 11293 64197 11379 64253
rect 11435 64197 11521 64253
rect 11577 64197 11663 64253
rect 11719 64197 11805 64253
rect 11861 64197 11947 64253
rect 12003 64197 12089 64253
rect 12145 64197 12231 64253
rect 12287 64197 12373 64253
rect 12429 64197 12515 64253
rect 12571 64197 12657 64253
rect 12713 64197 12799 64253
rect 12855 64197 12941 64253
rect 12997 64197 13083 64253
rect 13139 64197 13225 64253
rect 13281 64197 13367 64253
rect 13423 64197 13509 64253
rect 13565 64197 13651 64253
rect 13707 64197 13793 64253
rect 13849 64197 13935 64253
rect 13991 64197 14077 64253
rect 14133 64197 14219 64253
rect 14275 64197 14361 64253
rect 14417 64197 14503 64253
rect 14559 64197 14645 64253
rect 14701 64197 14787 64253
rect 14843 64197 15000 64253
rect 0 64111 15000 64197
rect 0 64055 161 64111
rect 217 64055 303 64111
rect 359 64055 445 64111
rect 501 64055 587 64111
rect 643 64055 729 64111
rect 785 64055 871 64111
rect 927 64055 1013 64111
rect 1069 64055 1155 64111
rect 1211 64055 1297 64111
rect 1353 64055 1439 64111
rect 1495 64055 1581 64111
rect 1637 64055 1723 64111
rect 1779 64055 1865 64111
rect 1921 64055 2007 64111
rect 2063 64055 2149 64111
rect 2205 64055 2291 64111
rect 2347 64055 2433 64111
rect 2489 64055 2575 64111
rect 2631 64055 2717 64111
rect 2773 64055 2859 64111
rect 2915 64055 3001 64111
rect 3057 64055 3143 64111
rect 3199 64055 3285 64111
rect 3341 64055 3427 64111
rect 3483 64055 3569 64111
rect 3625 64055 3711 64111
rect 3767 64055 3853 64111
rect 3909 64055 3995 64111
rect 4051 64055 4137 64111
rect 4193 64055 4279 64111
rect 4335 64055 4421 64111
rect 4477 64055 4563 64111
rect 4619 64055 4705 64111
rect 4761 64055 4847 64111
rect 4903 64055 4989 64111
rect 5045 64055 5131 64111
rect 5187 64055 5273 64111
rect 5329 64055 5415 64111
rect 5471 64055 5557 64111
rect 5613 64055 5699 64111
rect 5755 64055 5841 64111
rect 5897 64055 5983 64111
rect 6039 64055 6125 64111
rect 6181 64055 6267 64111
rect 6323 64055 6409 64111
rect 6465 64055 6551 64111
rect 6607 64055 6693 64111
rect 6749 64055 6835 64111
rect 6891 64055 6977 64111
rect 7033 64055 7119 64111
rect 7175 64055 7261 64111
rect 7317 64055 7403 64111
rect 7459 64055 7545 64111
rect 7601 64055 7687 64111
rect 7743 64055 7829 64111
rect 7885 64055 7971 64111
rect 8027 64055 8113 64111
rect 8169 64055 8255 64111
rect 8311 64055 8397 64111
rect 8453 64055 8539 64111
rect 8595 64055 8681 64111
rect 8737 64055 8823 64111
rect 8879 64055 8965 64111
rect 9021 64055 9107 64111
rect 9163 64055 9249 64111
rect 9305 64055 9391 64111
rect 9447 64055 9533 64111
rect 9589 64055 9675 64111
rect 9731 64055 9817 64111
rect 9873 64055 9959 64111
rect 10015 64055 10101 64111
rect 10157 64055 10243 64111
rect 10299 64055 10385 64111
rect 10441 64055 10527 64111
rect 10583 64055 10669 64111
rect 10725 64055 10811 64111
rect 10867 64055 10953 64111
rect 11009 64055 11095 64111
rect 11151 64055 11237 64111
rect 11293 64055 11379 64111
rect 11435 64055 11521 64111
rect 11577 64055 11663 64111
rect 11719 64055 11805 64111
rect 11861 64055 11947 64111
rect 12003 64055 12089 64111
rect 12145 64055 12231 64111
rect 12287 64055 12373 64111
rect 12429 64055 12515 64111
rect 12571 64055 12657 64111
rect 12713 64055 12799 64111
rect 12855 64055 12941 64111
rect 12997 64055 13083 64111
rect 13139 64055 13225 64111
rect 13281 64055 13367 64111
rect 13423 64055 13509 64111
rect 13565 64055 13651 64111
rect 13707 64055 13793 64111
rect 13849 64055 13935 64111
rect 13991 64055 14077 64111
rect 14133 64055 14219 64111
rect 14275 64055 14361 64111
rect 14417 64055 14503 64111
rect 14559 64055 14645 64111
rect 14701 64055 14787 64111
rect 14843 64055 15000 64111
rect 0 63969 15000 64055
rect 0 63913 161 63969
rect 217 63913 303 63969
rect 359 63913 445 63969
rect 501 63913 587 63969
rect 643 63913 729 63969
rect 785 63913 871 63969
rect 927 63913 1013 63969
rect 1069 63913 1155 63969
rect 1211 63913 1297 63969
rect 1353 63913 1439 63969
rect 1495 63913 1581 63969
rect 1637 63913 1723 63969
rect 1779 63913 1865 63969
rect 1921 63913 2007 63969
rect 2063 63913 2149 63969
rect 2205 63913 2291 63969
rect 2347 63913 2433 63969
rect 2489 63913 2575 63969
rect 2631 63913 2717 63969
rect 2773 63913 2859 63969
rect 2915 63913 3001 63969
rect 3057 63913 3143 63969
rect 3199 63913 3285 63969
rect 3341 63913 3427 63969
rect 3483 63913 3569 63969
rect 3625 63913 3711 63969
rect 3767 63913 3853 63969
rect 3909 63913 3995 63969
rect 4051 63913 4137 63969
rect 4193 63913 4279 63969
rect 4335 63913 4421 63969
rect 4477 63913 4563 63969
rect 4619 63913 4705 63969
rect 4761 63913 4847 63969
rect 4903 63913 4989 63969
rect 5045 63913 5131 63969
rect 5187 63913 5273 63969
rect 5329 63913 5415 63969
rect 5471 63913 5557 63969
rect 5613 63913 5699 63969
rect 5755 63913 5841 63969
rect 5897 63913 5983 63969
rect 6039 63913 6125 63969
rect 6181 63913 6267 63969
rect 6323 63913 6409 63969
rect 6465 63913 6551 63969
rect 6607 63913 6693 63969
rect 6749 63913 6835 63969
rect 6891 63913 6977 63969
rect 7033 63913 7119 63969
rect 7175 63913 7261 63969
rect 7317 63913 7403 63969
rect 7459 63913 7545 63969
rect 7601 63913 7687 63969
rect 7743 63913 7829 63969
rect 7885 63913 7971 63969
rect 8027 63913 8113 63969
rect 8169 63913 8255 63969
rect 8311 63913 8397 63969
rect 8453 63913 8539 63969
rect 8595 63913 8681 63969
rect 8737 63913 8823 63969
rect 8879 63913 8965 63969
rect 9021 63913 9107 63969
rect 9163 63913 9249 63969
rect 9305 63913 9391 63969
rect 9447 63913 9533 63969
rect 9589 63913 9675 63969
rect 9731 63913 9817 63969
rect 9873 63913 9959 63969
rect 10015 63913 10101 63969
rect 10157 63913 10243 63969
rect 10299 63913 10385 63969
rect 10441 63913 10527 63969
rect 10583 63913 10669 63969
rect 10725 63913 10811 63969
rect 10867 63913 10953 63969
rect 11009 63913 11095 63969
rect 11151 63913 11237 63969
rect 11293 63913 11379 63969
rect 11435 63913 11521 63969
rect 11577 63913 11663 63969
rect 11719 63913 11805 63969
rect 11861 63913 11947 63969
rect 12003 63913 12089 63969
rect 12145 63913 12231 63969
rect 12287 63913 12373 63969
rect 12429 63913 12515 63969
rect 12571 63913 12657 63969
rect 12713 63913 12799 63969
rect 12855 63913 12941 63969
rect 12997 63913 13083 63969
rect 13139 63913 13225 63969
rect 13281 63913 13367 63969
rect 13423 63913 13509 63969
rect 13565 63913 13651 63969
rect 13707 63913 13793 63969
rect 13849 63913 13935 63969
rect 13991 63913 14077 63969
rect 14133 63913 14219 63969
rect 14275 63913 14361 63969
rect 14417 63913 14503 63969
rect 14559 63913 14645 63969
rect 14701 63913 14787 63969
rect 14843 63913 15000 63969
rect 0 63827 15000 63913
rect 0 63771 161 63827
rect 217 63771 303 63827
rect 359 63771 445 63827
rect 501 63771 587 63827
rect 643 63771 729 63827
rect 785 63771 871 63827
rect 927 63771 1013 63827
rect 1069 63771 1155 63827
rect 1211 63771 1297 63827
rect 1353 63771 1439 63827
rect 1495 63771 1581 63827
rect 1637 63771 1723 63827
rect 1779 63771 1865 63827
rect 1921 63771 2007 63827
rect 2063 63771 2149 63827
rect 2205 63771 2291 63827
rect 2347 63771 2433 63827
rect 2489 63771 2575 63827
rect 2631 63771 2717 63827
rect 2773 63771 2859 63827
rect 2915 63771 3001 63827
rect 3057 63771 3143 63827
rect 3199 63771 3285 63827
rect 3341 63771 3427 63827
rect 3483 63771 3569 63827
rect 3625 63771 3711 63827
rect 3767 63771 3853 63827
rect 3909 63771 3995 63827
rect 4051 63771 4137 63827
rect 4193 63771 4279 63827
rect 4335 63771 4421 63827
rect 4477 63771 4563 63827
rect 4619 63771 4705 63827
rect 4761 63771 4847 63827
rect 4903 63771 4989 63827
rect 5045 63771 5131 63827
rect 5187 63771 5273 63827
rect 5329 63771 5415 63827
rect 5471 63771 5557 63827
rect 5613 63771 5699 63827
rect 5755 63771 5841 63827
rect 5897 63771 5983 63827
rect 6039 63771 6125 63827
rect 6181 63771 6267 63827
rect 6323 63771 6409 63827
rect 6465 63771 6551 63827
rect 6607 63771 6693 63827
rect 6749 63771 6835 63827
rect 6891 63771 6977 63827
rect 7033 63771 7119 63827
rect 7175 63771 7261 63827
rect 7317 63771 7403 63827
rect 7459 63771 7545 63827
rect 7601 63771 7687 63827
rect 7743 63771 7829 63827
rect 7885 63771 7971 63827
rect 8027 63771 8113 63827
rect 8169 63771 8255 63827
rect 8311 63771 8397 63827
rect 8453 63771 8539 63827
rect 8595 63771 8681 63827
rect 8737 63771 8823 63827
rect 8879 63771 8965 63827
rect 9021 63771 9107 63827
rect 9163 63771 9249 63827
rect 9305 63771 9391 63827
rect 9447 63771 9533 63827
rect 9589 63771 9675 63827
rect 9731 63771 9817 63827
rect 9873 63771 9959 63827
rect 10015 63771 10101 63827
rect 10157 63771 10243 63827
rect 10299 63771 10385 63827
rect 10441 63771 10527 63827
rect 10583 63771 10669 63827
rect 10725 63771 10811 63827
rect 10867 63771 10953 63827
rect 11009 63771 11095 63827
rect 11151 63771 11237 63827
rect 11293 63771 11379 63827
rect 11435 63771 11521 63827
rect 11577 63771 11663 63827
rect 11719 63771 11805 63827
rect 11861 63771 11947 63827
rect 12003 63771 12089 63827
rect 12145 63771 12231 63827
rect 12287 63771 12373 63827
rect 12429 63771 12515 63827
rect 12571 63771 12657 63827
rect 12713 63771 12799 63827
rect 12855 63771 12941 63827
rect 12997 63771 13083 63827
rect 13139 63771 13225 63827
rect 13281 63771 13367 63827
rect 13423 63771 13509 63827
rect 13565 63771 13651 63827
rect 13707 63771 13793 63827
rect 13849 63771 13935 63827
rect 13991 63771 14077 63827
rect 14133 63771 14219 63827
rect 14275 63771 14361 63827
rect 14417 63771 14503 63827
rect 14559 63771 14645 63827
rect 14701 63771 14787 63827
rect 14843 63771 15000 63827
rect 0 63685 15000 63771
rect 0 63629 161 63685
rect 217 63629 303 63685
rect 359 63629 445 63685
rect 501 63629 587 63685
rect 643 63629 729 63685
rect 785 63629 871 63685
rect 927 63629 1013 63685
rect 1069 63629 1155 63685
rect 1211 63629 1297 63685
rect 1353 63629 1439 63685
rect 1495 63629 1581 63685
rect 1637 63629 1723 63685
rect 1779 63629 1865 63685
rect 1921 63629 2007 63685
rect 2063 63629 2149 63685
rect 2205 63629 2291 63685
rect 2347 63629 2433 63685
rect 2489 63629 2575 63685
rect 2631 63629 2717 63685
rect 2773 63629 2859 63685
rect 2915 63629 3001 63685
rect 3057 63629 3143 63685
rect 3199 63629 3285 63685
rect 3341 63629 3427 63685
rect 3483 63629 3569 63685
rect 3625 63629 3711 63685
rect 3767 63629 3853 63685
rect 3909 63629 3995 63685
rect 4051 63629 4137 63685
rect 4193 63629 4279 63685
rect 4335 63629 4421 63685
rect 4477 63629 4563 63685
rect 4619 63629 4705 63685
rect 4761 63629 4847 63685
rect 4903 63629 4989 63685
rect 5045 63629 5131 63685
rect 5187 63629 5273 63685
rect 5329 63629 5415 63685
rect 5471 63629 5557 63685
rect 5613 63629 5699 63685
rect 5755 63629 5841 63685
rect 5897 63629 5983 63685
rect 6039 63629 6125 63685
rect 6181 63629 6267 63685
rect 6323 63629 6409 63685
rect 6465 63629 6551 63685
rect 6607 63629 6693 63685
rect 6749 63629 6835 63685
rect 6891 63629 6977 63685
rect 7033 63629 7119 63685
rect 7175 63629 7261 63685
rect 7317 63629 7403 63685
rect 7459 63629 7545 63685
rect 7601 63629 7687 63685
rect 7743 63629 7829 63685
rect 7885 63629 7971 63685
rect 8027 63629 8113 63685
rect 8169 63629 8255 63685
rect 8311 63629 8397 63685
rect 8453 63629 8539 63685
rect 8595 63629 8681 63685
rect 8737 63629 8823 63685
rect 8879 63629 8965 63685
rect 9021 63629 9107 63685
rect 9163 63629 9249 63685
rect 9305 63629 9391 63685
rect 9447 63629 9533 63685
rect 9589 63629 9675 63685
rect 9731 63629 9817 63685
rect 9873 63629 9959 63685
rect 10015 63629 10101 63685
rect 10157 63629 10243 63685
rect 10299 63629 10385 63685
rect 10441 63629 10527 63685
rect 10583 63629 10669 63685
rect 10725 63629 10811 63685
rect 10867 63629 10953 63685
rect 11009 63629 11095 63685
rect 11151 63629 11237 63685
rect 11293 63629 11379 63685
rect 11435 63629 11521 63685
rect 11577 63629 11663 63685
rect 11719 63629 11805 63685
rect 11861 63629 11947 63685
rect 12003 63629 12089 63685
rect 12145 63629 12231 63685
rect 12287 63629 12373 63685
rect 12429 63629 12515 63685
rect 12571 63629 12657 63685
rect 12713 63629 12799 63685
rect 12855 63629 12941 63685
rect 12997 63629 13083 63685
rect 13139 63629 13225 63685
rect 13281 63629 13367 63685
rect 13423 63629 13509 63685
rect 13565 63629 13651 63685
rect 13707 63629 13793 63685
rect 13849 63629 13935 63685
rect 13991 63629 14077 63685
rect 14133 63629 14219 63685
rect 14275 63629 14361 63685
rect 14417 63629 14503 63685
rect 14559 63629 14645 63685
rect 14701 63629 14787 63685
rect 14843 63629 15000 63685
rect 0 63600 15000 63629
rect 0 63371 15000 63400
rect 0 63315 161 63371
rect 217 63315 303 63371
rect 359 63315 445 63371
rect 501 63315 587 63371
rect 643 63315 729 63371
rect 785 63315 871 63371
rect 927 63315 1013 63371
rect 1069 63315 1155 63371
rect 1211 63315 1297 63371
rect 1353 63315 1439 63371
rect 1495 63315 1581 63371
rect 1637 63315 1723 63371
rect 1779 63315 1865 63371
rect 1921 63315 2007 63371
rect 2063 63315 2149 63371
rect 2205 63315 2291 63371
rect 2347 63315 2433 63371
rect 2489 63315 2575 63371
rect 2631 63315 2717 63371
rect 2773 63315 2859 63371
rect 2915 63315 3001 63371
rect 3057 63315 3143 63371
rect 3199 63315 3285 63371
rect 3341 63315 3427 63371
rect 3483 63315 3569 63371
rect 3625 63315 3711 63371
rect 3767 63315 3853 63371
rect 3909 63315 3995 63371
rect 4051 63315 4137 63371
rect 4193 63315 4279 63371
rect 4335 63315 4421 63371
rect 4477 63315 4563 63371
rect 4619 63315 4705 63371
rect 4761 63315 4847 63371
rect 4903 63315 4989 63371
rect 5045 63315 5131 63371
rect 5187 63315 5273 63371
rect 5329 63315 5415 63371
rect 5471 63315 5557 63371
rect 5613 63315 5699 63371
rect 5755 63315 5841 63371
rect 5897 63315 5983 63371
rect 6039 63315 6125 63371
rect 6181 63315 6267 63371
rect 6323 63315 6409 63371
rect 6465 63315 6551 63371
rect 6607 63315 6693 63371
rect 6749 63315 6835 63371
rect 6891 63315 6977 63371
rect 7033 63315 7119 63371
rect 7175 63315 7261 63371
rect 7317 63315 7403 63371
rect 7459 63315 7545 63371
rect 7601 63315 7687 63371
rect 7743 63315 7829 63371
rect 7885 63315 7971 63371
rect 8027 63315 8113 63371
rect 8169 63315 8255 63371
rect 8311 63315 8397 63371
rect 8453 63315 8539 63371
rect 8595 63315 8681 63371
rect 8737 63315 8823 63371
rect 8879 63315 8965 63371
rect 9021 63315 9107 63371
rect 9163 63315 9249 63371
rect 9305 63315 9391 63371
rect 9447 63315 9533 63371
rect 9589 63315 9675 63371
rect 9731 63315 9817 63371
rect 9873 63315 9959 63371
rect 10015 63315 10101 63371
rect 10157 63315 10243 63371
rect 10299 63315 10385 63371
rect 10441 63315 10527 63371
rect 10583 63315 10669 63371
rect 10725 63315 10811 63371
rect 10867 63315 10953 63371
rect 11009 63315 11095 63371
rect 11151 63315 11237 63371
rect 11293 63315 11379 63371
rect 11435 63315 11521 63371
rect 11577 63315 11663 63371
rect 11719 63315 11805 63371
rect 11861 63315 11947 63371
rect 12003 63315 12089 63371
rect 12145 63315 12231 63371
rect 12287 63315 12373 63371
rect 12429 63315 12515 63371
rect 12571 63315 12657 63371
rect 12713 63315 12799 63371
rect 12855 63315 12941 63371
rect 12997 63315 13083 63371
rect 13139 63315 13225 63371
rect 13281 63315 13367 63371
rect 13423 63315 13509 63371
rect 13565 63315 13651 63371
rect 13707 63315 13793 63371
rect 13849 63315 13935 63371
rect 13991 63315 14077 63371
rect 14133 63315 14219 63371
rect 14275 63315 14361 63371
rect 14417 63315 14503 63371
rect 14559 63315 14645 63371
rect 14701 63315 14787 63371
rect 14843 63315 15000 63371
rect 0 63229 15000 63315
rect 0 63173 161 63229
rect 217 63173 303 63229
rect 359 63173 445 63229
rect 501 63173 587 63229
rect 643 63173 729 63229
rect 785 63173 871 63229
rect 927 63173 1013 63229
rect 1069 63173 1155 63229
rect 1211 63173 1297 63229
rect 1353 63173 1439 63229
rect 1495 63173 1581 63229
rect 1637 63173 1723 63229
rect 1779 63173 1865 63229
rect 1921 63173 2007 63229
rect 2063 63173 2149 63229
rect 2205 63173 2291 63229
rect 2347 63173 2433 63229
rect 2489 63173 2575 63229
rect 2631 63173 2717 63229
rect 2773 63173 2859 63229
rect 2915 63173 3001 63229
rect 3057 63173 3143 63229
rect 3199 63173 3285 63229
rect 3341 63173 3427 63229
rect 3483 63173 3569 63229
rect 3625 63173 3711 63229
rect 3767 63173 3853 63229
rect 3909 63173 3995 63229
rect 4051 63173 4137 63229
rect 4193 63173 4279 63229
rect 4335 63173 4421 63229
rect 4477 63173 4563 63229
rect 4619 63173 4705 63229
rect 4761 63173 4847 63229
rect 4903 63173 4989 63229
rect 5045 63173 5131 63229
rect 5187 63173 5273 63229
rect 5329 63173 5415 63229
rect 5471 63173 5557 63229
rect 5613 63173 5699 63229
rect 5755 63173 5841 63229
rect 5897 63173 5983 63229
rect 6039 63173 6125 63229
rect 6181 63173 6267 63229
rect 6323 63173 6409 63229
rect 6465 63173 6551 63229
rect 6607 63173 6693 63229
rect 6749 63173 6835 63229
rect 6891 63173 6977 63229
rect 7033 63173 7119 63229
rect 7175 63173 7261 63229
rect 7317 63173 7403 63229
rect 7459 63173 7545 63229
rect 7601 63173 7687 63229
rect 7743 63173 7829 63229
rect 7885 63173 7971 63229
rect 8027 63173 8113 63229
rect 8169 63173 8255 63229
rect 8311 63173 8397 63229
rect 8453 63173 8539 63229
rect 8595 63173 8681 63229
rect 8737 63173 8823 63229
rect 8879 63173 8965 63229
rect 9021 63173 9107 63229
rect 9163 63173 9249 63229
rect 9305 63173 9391 63229
rect 9447 63173 9533 63229
rect 9589 63173 9675 63229
rect 9731 63173 9817 63229
rect 9873 63173 9959 63229
rect 10015 63173 10101 63229
rect 10157 63173 10243 63229
rect 10299 63173 10385 63229
rect 10441 63173 10527 63229
rect 10583 63173 10669 63229
rect 10725 63173 10811 63229
rect 10867 63173 10953 63229
rect 11009 63173 11095 63229
rect 11151 63173 11237 63229
rect 11293 63173 11379 63229
rect 11435 63173 11521 63229
rect 11577 63173 11663 63229
rect 11719 63173 11805 63229
rect 11861 63173 11947 63229
rect 12003 63173 12089 63229
rect 12145 63173 12231 63229
rect 12287 63173 12373 63229
rect 12429 63173 12515 63229
rect 12571 63173 12657 63229
rect 12713 63173 12799 63229
rect 12855 63173 12941 63229
rect 12997 63173 13083 63229
rect 13139 63173 13225 63229
rect 13281 63173 13367 63229
rect 13423 63173 13509 63229
rect 13565 63173 13651 63229
rect 13707 63173 13793 63229
rect 13849 63173 13935 63229
rect 13991 63173 14077 63229
rect 14133 63173 14219 63229
rect 14275 63173 14361 63229
rect 14417 63173 14503 63229
rect 14559 63173 14645 63229
rect 14701 63173 14787 63229
rect 14843 63173 15000 63229
rect 0 63087 15000 63173
rect 0 63031 161 63087
rect 217 63031 303 63087
rect 359 63031 445 63087
rect 501 63031 587 63087
rect 643 63031 729 63087
rect 785 63031 871 63087
rect 927 63031 1013 63087
rect 1069 63031 1155 63087
rect 1211 63031 1297 63087
rect 1353 63031 1439 63087
rect 1495 63031 1581 63087
rect 1637 63031 1723 63087
rect 1779 63031 1865 63087
rect 1921 63031 2007 63087
rect 2063 63031 2149 63087
rect 2205 63031 2291 63087
rect 2347 63031 2433 63087
rect 2489 63031 2575 63087
rect 2631 63031 2717 63087
rect 2773 63031 2859 63087
rect 2915 63031 3001 63087
rect 3057 63031 3143 63087
rect 3199 63031 3285 63087
rect 3341 63031 3427 63087
rect 3483 63031 3569 63087
rect 3625 63031 3711 63087
rect 3767 63031 3853 63087
rect 3909 63031 3995 63087
rect 4051 63031 4137 63087
rect 4193 63031 4279 63087
rect 4335 63031 4421 63087
rect 4477 63031 4563 63087
rect 4619 63031 4705 63087
rect 4761 63031 4847 63087
rect 4903 63031 4989 63087
rect 5045 63031 5131 63087
rect 5187 63031 5273 63087
rect 5329 63031 5415 63087
rect 5471 63031 5557 63087
rect 5613 63031 5699 63087
rect 5755 63031 5841 63087
rect 5897 63031 5983 63087
rect 6039 63031 6125 63087
rect 6181 63031 6267 63087
rect 6323 63031 6409 63087
rect 6465 63031 6551 63087
rect 6607 63031 6693 63087
rect 6749 63031 6835 63087
rect 6891 63031 6977 63087
rect 7033 63031 7119 63087
rect 7175 63031 7261 63087
rect 7317 63031 7403 63087
rect 7459 63031 7545 63087
rect 7601 63031 7687 63087
rect 7743 63031 7829 63087
rect 7885 63031 7971 63087
rect 8027 63031 8113 63087
rect 8169 63031 8255 63087
rect 8311 63031 8397 63087
rect 8453 63031 8539 63087
rect 8595 63031 8681 63087
rect 8737 63031 8823 63087
rect 8879 63031 8965 63087
rect 9021 63031 9107 63087
rect 9163 63031 9249 63087
rect 9305 63031 9391 63087
rect 9447 63031 9533 63087
rect 9589 63031 9675 63087
rect 9731 63031 9817 63087
rect 9873 63031 9959 63087
rect 10015 63031 10101 63087
rect 10157 63031 10243 63087
rect 10299 63031 10385 63087
rect 10441 63031 10527 63087
rect 10583 63031 10669 63087
rect 10725 63031 10811 63087
rect 10867 63031 10953 63087
rect 11009 63031 11095 63087
rect 11151 63031 11237 63087
rect 11293 63031 11379 63087
rect 11435 63031 11521 63087
rect 11577 63031 11663 63087
rect 11719 63031 11805 63087
rect 11861 63031 11947 63087
rect 12003 63031 12089 63087
rect 12145 63031 12231 63087
rect 12287 63031 12373 63087
rect 12429 63031 12515 63087
rect 12571 63031 12657 63087
rect 12713 63031 12799 63087
rect 12855 63031 12941 63087
rect 12997 63031 13083 63087
rect 13139 63031 13225 63087
rect 13281 63031 13367 63087
rect 13423 63031 13509 63087
rect 13565 63031 13651 63087
rect 13707 63031 13793 63087
rect 13849 63031 13935 63087
rect 13991 63031 14077 63087
rect 14133 63031 14219 63087
rect 14275 63031 14361 63087
rect 14417 63031 14503 63087
rect 14559 63031 14645 63087
rect 14701 63031 14787 63087
rect 14843 63031 15000 63087
rect 0 62945 15000 63031
rect 0 62889 161 62945
rect 217 62889 303 62945
rect 359 62889 445 62945
rect 501 62889 587 62945
rect 643 62889 729 62945
rect 785 62889 871 62945
rect 927 62889 1013 62945
rect 1069 62889 1155 62945
rect 1211 62889 1297 62945
rect 1353 62889 1439 62945
rect 1495 62889 1581 62945
rect 1637 62889 1723 62945
rect 1779 62889 1865 62945
rect 1921 62889 2007 62945
rect 2063 62889 2149 62945
rect 2205 62889 2291 62945
rect 2347 62889 2433 62945
rect 2489 62889 2575 62945
rect 2631 62889 2717 62945
rect 2773 62889 2859 62945
rect 2915 62889 3001 62945
rect 3057 62889 3143 62945
rect 3199 62889 3285 62945
rect 3341 62889 3427 62945
rect 3483 62889 3569 62945
rect 3625 62889 3711 62945
rect 3767 62889 3853 62945
rect 3909 62889 3995 62945
rect 4051 62889 4137 62945
rect 4193 62889 4279 62945
rect 4335 62889 4421 62945
rect 4477 62889 4563 62945
rect 4619 62889 4705 62945
rect 4761 62889 4847 62945
rect 4903 62889 4989 62945
rect 5045 62889 5131 62945
rect 5187 62889 5273 62945
rect 5329 62889 5415 62945
rect 5471 62889 5557 62945
rect 5613 62889 5699 62945
rect 5755 62889 5841 62945
rect 5897 62889 5983 62945
rect 6039 62889 6125 62945
rect 6181 62889 6267 62945
rect 6323 62889 6409 62945
rect 6465 62889 6551 62945
rect 6607 62889 6693 62945
rect 6749 62889 6835 62945
rect 6891 62889 6977 62945
rect 7033 62889 7119 62945
rect 7175 62889 7261 62945
rect 7317 62889 7403 62945
rect 7459 62889 7545 62945
rect 7601 62889 7687 62945
rect 7743 62889 7829 62945
rect 7885 62889 7971 62945
rect 8027 62889 8113 62945
rect 8169 62889 8255 62945
rect 8311 62889 8397 62945
rect 8453 62889 8539 62945
rect 8595 62889 8681 62945
rect 8737 62889 8823 62945
rect 8879 62889 8965 62945
rect 9021 62889 9107 62945
rect 9163 62889 9249 62945
rect 9305 62889 9391 62945
rect 9447 62889 9533 62945
rect 9589 62889 9675 62945
rect 9731 62889 9817 62945
rect 9873 62889 9959 62945
rect 10015 62889 10101 62945
rect 10157 62889 10243 62945
rect 10299 62889 10385 62945
rect 10441 62889 10527 62945
rect 10583 62889 10669 62945
rect 10725 62889 10811 62945
rect 10867 62889 10953 62945
rect 11009 62889 11095 62945
rect 11151 62889 11237 62945
rect 11293 62889 11379 62945
rect 11435 62889 11521 62945
rect 11577 62889 11663 62945
rect 11719 62889 11805 62945
rect 11861 62889 11947 62945
rect 12003 62889 12089 62945
rect 12145 62889 12231 62945
rect 12287 62889 12373 62945
rect 12429 62889 12515 62945
rect 12571 62889 12657 62945
rect 12713 62889 12799 62945
rect 12855 62889 12941 62945
rect 12997 62889 13083 62945
rect 13139 62889 13225 62945
rect 13281 62889 13367 62945
rect 13423 62889 13509 62945
rect 13565 62889 13651 62945
rect 13707 62889 13793 62945
rect 13849 62889 13935 62945
rect 13991 62889 14077 62945
rect 14133 62889 14219 62945
rect 14275 62889 14361 62945
rect 14417 62889 14503 62945
rect 14559 62889 14645 62945
rect 14701 62889 14787 62945
rect 14843 62889 15000 62945
rect 0 62803 15000 62889
rect 0 62747 161 62803
rect 217 62747 303 62803
rect 359 62747 445 62803
rect 501 62747 587 62803
rect 643 62747 729 62803
rect 785 62747 871 62803
rect 927 62747 1013 62803
rect 1069 62747 1155 62803
rect 1211 62747 1297 62803
rect 1353 62747 1439 62803
rect 1495 62747 1581 62803
rect 1637 62747 1723 62803
rect 1779 62747 1865 62803
rect 1921 62747 2007 62803
rect 2063 62747 2149 62803
rect 2205 62747 2291 62803
rect 2347 62747 2433 62803
rect 2489 62747 2575 62803
rect 2631 62747 2717 62803
rect 2773 62747 2859 62803
rect 2915 62747 3001 62803
rect 3057 62747 3143 62803
rect 3199 62747 3285 62803
rect 3341 62747 3427 62803
rect 3483 62747 3569 62803
rect 3625 62747 3711 62803
rect 3767 62747 3853 62803
rect 3909 62747 3995 62803
rect 4051 62747 4137 62803
rect 4193 62747 4279 62803
rect 4335 62747 4421 62803
rect 4477 62747 4563 62803
rect 4619 62747 4705 62803
rect 4761 62747 4847 62803
rect 4903 62747 4989 62803
rect 5045 62747 5131 62803
rect 5187 62747 5273 62803
rect 5329 62747 5415 62803
rect 5471 62747 5557 62803
rect 5613 62747 5699 62803
rect 5755 62747 5841 62803
rect 5897 62747 5983 62803
rect 6039 62747 6125 62803
rect 6181 62747 6267 62803
rect 6323 62747 6409 62803
rect 6465 62747 6551 62803
rect 6607 62747 6693 62803
rect 6749 62747 6835 62803
rect 6891 62747 6977 62803
rect 7033 62747 7119 62803
rect 7175 62747 7261 62803
rect 7317 62747 7403 62803
rect 7459 62747 7545 62803
rect 7601 62747 7687 62803
rect 7743 62747 7829 62803
rect 7885 62747 7971 62803
rect 8027 62747 8113 62803
rect 8169 62747 8255 62803
rect 8311 62747 8397 62803
rect 8453 62747 8539 62803
rect 8595 62747 8681 62803
rect 8737 62747 8823 62803
rect 8879 62747 8965 62803
rect 9021 62747 9107 62803
rect 9163 62747 9249 62803
rect 9305 62747 9391 62803
rect 9447 62747 9533 62803
rect 9589 62747 9675 62803
rect 9731 62747 9817 62803
rect 9873 62747 9959 62803
rect 10015 62747 10101 62803
rect 10157 62747 10243 62803
rect 10299 62747 10385 62803
rect 10441 62747 10527 62803
rect 10583 62747 10669 62803
rect 10725 62747 10811 62803
rect 10867 62747 10953 62803
rect 11009 62747 11095 62803
rect 11151 62747 11237 62803
rect 11293 62747 11379 62803
rect 11435 62747 11521 62803
rect 11577 62747 11663 62803
rect 11719 62747 11805 62803
rect 11861 62747 11947 62803
rect 12003 62747 12089 62803
rect 12145 62747 12231 62803
rect 12287 62747 12373 62803
rect 12429 62747 12515 62803
rect 12571 62747 12657 62803
rect 12713 62747 12799 62803
rect 12855 62747 12941 62803
rect 12997 62747 13083 62803
rect 13139 62747 13225 62803
rect 13281 62747 13367 62803
rect 13423 62747 13509 62803
rect 13565 62747 13651 62803
rect 13707 62747 13793 62803
rect 13849 62747 13935 62803
rect 13991 62747 14077 62803
rect 14133 62747 14219 62803
rect 14275 62747 14361 62803
rect 14417 62747 14503 62803
rect 14559 62747 14645 62803
rect 14701 62747 14787 62803
rect 14843 62747 15000 62803
rect 0 62661 15000 62747
rect 0 62605 161 62661
rect 217 62605 303 62661
rect 359 62605 445 62661
rect 501 62605 587 62661
rect 643 62605 729 62661
rect 785 62605 871 62661
rect 927 62605 1013 62661
rect 1069 62605 1155 62661
rect 1211 62605 1297 62661
rect 1353 62605 1439 62661
rect 1495 62605 1581 62661
rect 1637 62605 1723 62661
rect 1779 62605 1865 62661
rect 1921 62605 2007 62661
rect 2063 62605 2149 62661
rect 2205 62605 2291 62661
rect 2347 62605 2433 62661
rect 2489 62605 2575 62661
rect 2631 62605 2717 62661
rect 2773 62605 2859 62661
rect 2915 62605 3001 62661
rect 3057 62605 3143 62661
rect 3199 62605 3285 62661
rect 3341 62605 3427 62661
rect 3483 62605 3569 62661
rect 3625 62605 3711 62661
rect 3767 62605 3853 62661
rect 3909 62605 3995 62661
rect 4051 62605 4137 62661
rect 4193 62605 4279 62661
rect 4335 62605 4421 62661
rect 4477 62605 4563 62661
rect 4619 62605 4705 62661
rect 4761 62605 4847 62661
rect 4903 62605 4989 62661
rect 5045 62605 5131 62661
rect 5187 62605 5273 62661
rect 5329 62605 5415 62661
rect 5471 62605 5557 62661
rect 5613 62605 5699 62661
rect 5755 62605 5841 62661
rect 5897 62605 5983 62661
rect 6039 62605 6125 62661
rect 6181 62605 6267 62661
rect 6323 62605 6409 62661
rect 6465 62605 6551 62661
rect 6607 62605 6693 62661
rect 6749 62605 6835 62661
rect 6891 62605 6977 62661
rect 7033 62605 7119 62661
rect 7175 62605 7261 62661
rect 7317 62605 7403 62661
rect 7459 62605 7545 62661
rect 7601 62605 7687 62661
rect 7743 62605 7829 62661
rect 7885 62605 7971 62661
rect 8027 62605 8113 62661
rect 8169 62605 8255 62661
rect 8311 62605 8397 62661
rect 8453 62605 8539 62661
rect 8595 62605 8681 62661
rect 8737 62605 8823 62661
rect 8879 62605 8965 62661
rect 9021 62605 9107 62661
rect 9163 62605 9249 62661
rect 9305 62605 9391 62661
rect 9447 62605 9533 62661
rect 9589 62605 9675 62661
rect 9731 62605 9817 62661
rect 9873 62605 9959 62661
rect 10015 62605 10101 62661
rect 10157 62605 10243 62661
rect 10299 62605 10385 62661
rect 10441 62605 10527 62661
rect 10583 62605 10669 62661
rect 10725 62605 10811 62661
rect 10867 62605 10953 62661
rect 11009 62605 11095 62661
rect 11151 62605 11237 62661
rect 11293 62605 11379 62661
rect 11435 62605 11521 62661
rect 11577 62605 11663 62661
rect 11719 62605 11805 62661
rect 11861 62605 11947 62661
rect 12003 62605 12089 62661
rect 12145 62605 12231 62661
rect 12287 62605 12373 62661
rect 12429 62605 12515 62661
rect 12571 62605 12657 62661
rect 12713 62605 12799 62661
rect 12855 62605 12941 62661
rect 12997 62605 13083 62661
rect 13139 62605 13225 62661
rect 13281 62605 13367 62661
rect 13423 62605 13509 62661
rect 13565 62605 13651 62661
rect 13707 62605 13793 62661
rect 13849 62605 13935 62661
rect 13991 62605 14077 62661
rect 14133 62605 14219 62661
rect 14275 62605 14361 62661
rect 14417 62605 14503 62661
rect 14559 62605 14645 62661
rect 14701 62605 14787 62661
rect 14843 62605 15000 62661
rect 0 62519 15000 62605
rect 0 62463 161 62519
rect 217 62463 303 62519
rect 359 62463 445 62519
rect 501 62463 587 62519
rect 643 62463 729 62519
rect 785 62463 871 62519
rect 927 62463 1013 62519
rect 1069 62463 1155 62519
rect 1211 62463 1297 62519
rect 1353 62463 1439 62519
rect 1495 62463 1581 62519
rect 1637 62463 1723 62519
rect 1779 62463 1865 62519
rect 1921 62463 2007 62519
rect 2063 62463 2149 62519
rect 2205 62463 2291 62519
rect 2347 62463 2433 62519
rect 2489 62463 2575 62519
rect 2631 62463 2717 62519
rect 2773 62463 2859 62519
rect 2915 62463 3001 62519
rect 3057 62463 3143 62519
rect 3199 62463 3285 62519
rect 3341 62463 3427 62519
rect 3483 62463 3569 62519
rect 3625 62463 3711 62519
rect 3767 62463 3853 62519
rect 3909 62463 3995 62519
rect 4051 62463 4137 62519
rect 4193 62463 4279 62519
rect 4335 62463 4421 62519
rect 4477 62463 4563 62519
rect 4619 62463 4705 62519
rect 4761 62463 4847 62519
rect 4903 62463 4989 62519
rect 5045 62463 5131 62519
rect 5187 62463 5273 62519
rect 5329 62463 5415 62519
rect 5471 62463 5557 62519
rect 5613 62463 5699 62519
rect 5755 62463 5841 62519
rect 5897 62463 5983 62519
rect 6039 62463 6125 62519
rect 6181 62463 6267 62519
rect 6323 62463 6409 62519
rect 6465 62463 6551 62519
rect 6607 62463 6693 62519
rect 6749 62463 6835 62519
rect 6891 62463 6977 62519
rect 7033 62463 7119 62519
rect 7175 62463 7261 62519
rect 7317 62463 7403 62519
rect 7459 62463 7545 62519
rect 7601 62463 7687 62519
rect 7743 62463 7829 62519
rect 7885 62463 7971 62519
rect 8027 62463 8113 62519
rect 8169 62463 8255 62519
rect 8311 62463 8397 62519
rect 8453 62463 8539 62519
rect 8595 62463 8681 62519
rect 8737 62463 8823 62519
rect 8879 62463 8965 62519
rect 9021 62463 9107 62519
rect 9163 62463 9249 62519
rect 9305 62463 9391 62519
rect 9447 62463 9533 62519
rect 9589 62463 9675 62519
rect 9731 62463 9817 62519
rect 9873 62463 9959 62519
rect 10015 62463 10101 62519
rect 10157 62463 10243 62519
rect 10299 62463 10385 62519
rect 10441 62463 10527 62519
rect 10583 62463 10669 62519
rect 10725 62463 10811 62519
rect 10867 62463 10953 62519
rect 11009 62463 11095 62519
rect 11151 62463 11237 62519
rect 11293 62463 11379 62519
rect 11435 62463 11521 62519
rect 11577 62463 11663 62519
rect 11719 62463 11805 62519
rect 11861 62463 11947 62519
rect 12003 62463 12089 62519
rect 12145 62463 12231 62519
rect 12287 62463 12373 62519
rect 12429 62463 12515 62519
rect 12571 62463 12657 62519
rect 12713 62463 12799 62519
rect 12855 62463 12941 62519
rect 12997 62463 13083 62519
rect 13139 62463 13225 62519
rect 13281 62463 13367 62519
rect 13423 62463 13509 62519
rect 13565 62463 13651 62519
rect 13707 62463 13793 62519
rect 13849 62463 13935 62519
rect 13991 62463 14077 62519
rect 14133 62463 14219 62519
rect 14275 62463 14361 62519
rect 14417 62463 14503 62519
rect 14559 62463 14645 62519
rect 14701 62463 14787 62519
rect 14843 62463 15000 62519
rect 0 62377 15000 62463
rect 0 62321 161 62377
rect 217 62321 303 62377
rect 359 62321 445 62377
rect 501 62321 587 62377
rect 643 62321 729 62377
rect 785 62321 871 62377
rect 927 62321 1013 62377
rect 1069 62321 1155 62377
rect 1211 62321 1297 62377
rect 1353 62321 1439 62377
rect 1495 62321 1581 62377
rect 1637 62321 1723 62377
rect 1779 62321 1865 62377
rect 1921 62321 2007 62377
rect 2063 62321 2149 62377
rect 2205 62321 2291 62377
rect 2347 62321 2433 62377
rect 2489 62321 2575 62377
rect 2631 62321 2717 62377
rect 2773 62321 2859 62377
rect 2915 62321 3001 62377
rect 3057 62321 3143 62377
rect 3199 62321 3285 62377
rect 3341 62321 3427 62377
rect 3483 62321 3569 62377
rect 3625 62321 3711 62377
rect 3767 62321 3853 62377
rect 3909 62321 3995 62377
rect 4051 62321 4137 62377
rect 4193 62321 4279 62377
rect 4335 62321 4421 62377
rect 4477 62321 4563 62377
rect 4619 62321 4705 62377
rect 4761 62321 4847 62377
rect 4903 62321 4989 62377
rect 5045 62321 5131 62377
rect 5187 62321 5273 62377
rect 5329 62321 5415 62377
rect 5471 62321 5557 62377
rect 5613 62321 5699 62377
rect 5755 62321 5841 62377
rect 5897 62321 5983 62377
rect 6039 62321 6125 62377
rect 6181 62321 6267 62377
rect 6323 62321 6409 62377
rect 6465 62321 6551 62377
rect 6607 62321 6693 62377
rect 6749 62321 6835 62377
rect 6891 62321 6977 62377
rect 7033 62321 7119 62377
rect 7175 62321 7261 62377
rect 7317 62321 7403 62377
rect 7459 62321 7545 62377
rect 7601 62321 7687 62377
rect 7743 62321 7829 62377
rect 7885 62321 7971 62377
rect 8027 62321 8113 62377
rect 8169 62321 8255 62377
rect 8311 62321 8397 62377
rect 8453 62321 8539 62377
rect 8595 62321 8681 62377
rect 8737 62321 8823 62377
rect 8879 62321 8965 62377
rect 9021 62321 9107 62377
rect 9163 62321 9249 62377
rect 9305 62321 9391 62377
rect 9447 62321 9533 62377
rect 9589 62321 9675 62377
rect 9731 62321 9817 62377
rect 9873 62321 9959 62377
rect 10015 62321 10101 62377
rect 10157 62321 10243 62377
rect 10299 62321 10385 62377
rect 10441 62321 10527 62377
rect 10583 62321 10669 62377
rect 10725 62321 10811 62377
rect 10867 62321 10953 62377
rect 11009 62321 11095 62377
rect 11151 62321 11237 62377
rect 11293 62321 11379 62377
rect 11435 62321 11521 62377
rect 11577 62321 11663 62377
rect 11719 62321 11805 62377
rect 11861 62321 11947 62377
rect 12003 62321 12089 62377
rect 12145 62321 12231 62377
rect 12287 62321 12373 62377
rect 12429 62321 12515 62377
rect 12571 62321 12657 62377
rect 12713 62321 12799 62377
rect 12855 62321 12941 62377
rect 12997 62321 13083 62377
rect 13139 62321 13225 62377
rect 13281 62321 13367 62377
rect 13423 62321 13509 62377
rect 13565 62321 13651 62377
rect 13707 62321 13793 62377
rect 13849 62321 13935 62377
rect 13991 62321 14077 62377
rect 14133 62321 14219 62377
rect 14275 62321 14361 62377
rect 14417 62321 14503 62377
rect 14559 62321 14645 62377
rect 14701 62321 14787 62377
rect 14843 62321 15000 62377
rect 0 62235 15000 62321
rect 0 62179 161 62235
rect 217 62179 303 62235
rect 359 62179 445 62235
rect 501 62179 587 62235
rect 643 62179 729 62235
rect 785 62179 871 62235
rect 927 62179 1013 62235
rect 1069 62179 1155 62235
rect 1211 62179 1297 62235
rect 1353 62179 1439 62235
rect 1495 62179 1581 62235
rect 1637 62179 1723 62235
rect 1779 62179 1865 62235
rect 1921 62179 2007 62235
rect 2063 62179 2149 62235
rect 2205 62179 2291 62235
rect 2347 62179 2433 62235
rect 2489 62179 2575 62235
rect 2631 62179 2717 62235
rect 2773 62179 2859 62235
rect 2915 62179 3001 62235
rect 3057 62179 3143 62235
rect 3199 62179 3285 62235
rect 3341 62179 3427 62235
rect 3483 62179 3569 62235
rect 3625 62179 3711 62235
rect 3767 62179 3853 62235
rect 3909 62179 3995 62235
rect 4051 62179 4137 62235
rect 4193 62179 4279 62235
rect 4335 62179 4421 62235
rect 4477 62179 4563 62235
rect 4619 62179 4705 62235
rect 4761 62179 4847 62235
rect 4903 62179 4989 62235
rect 5045 62179 5131 62235
rect 5187 62179 5273 62235
rect 5329 62179 5415 62235
rect 5471 62179 5557 62235
rect 5613 62179 5699 62235
rect 5755 62179 5841 62235
rect 5897 62179 5983 62235
rect 6039 62179 6125 62235
rect 6181 62179 6267 62235
rect 6323 62179 6409 62235
rect 6465 62179 6551 62235
rect 6607 62179 6693 62235
rect 6749 62179 6835 62235
rect 6891 62179 6977 62235
rect 7033 62179 7119 62235
rect 7175 62179 7261 62235
rect 7317 62179 7403 62235
rect 7459 62179 7545 62235
rect 7601 62179 7687 62235
rect 7743 62179 7829 62235
rect 7885 62179 7971 62235
rect 8027 62179 8113 62235
rect 8169 62179 8255 62235
rect 8311 62179 8397 62235
rect 8453 62179 8539 62235
rect 8595 62179 8681 62235
rect 8737 62179 8823 62235
rect 8879 62179 8965 62235
rect 9021 62179 9107 62235
rect 9163 62179 9249 62235
rect 9305 62179 9391 62235
rect 9447 62179 9533 62235
rect 9589 62179 9675 62235
rect 9731 62179 9817 62235
rect 9873 62179 9959 62235
rect 10015 62179 10101 62235
rect 10157 62179 10243 62235
rect 10299 62179 10385 62235
rect 10441 62179 10527 62235
rect 10583 62179 10669 62235
rect 10725 62179 10811 62235
rect 10867 62179 10953 62235
rect 11009 62179 11095 62235
rect 11151 62179 11237 62235
rect 11293 62179 11379 62235
rect 11435 62179 11521 62235
rect 11577 62179 11663 62235
rect 11719 62179 11805 62235
rect 11861 62179 11947 62235
rect 12003 62179 12089 62235
rect 12145 62179 12231 62235
rect 12287 62179 12373 62235
rect 12429 62179 12515 62235
rect 12571 62179 12657 62235
rect 12713 62179 12799 62235
rect 12855 62179 12941 62235
rect 12997 62179 13083 62235
rect 13139 62179 13225 62235
rect 13281 62179 13367 62235
rect 13423 62179 13509 62235
rect 13565 62179 13651 62235
rect 13707 62179 13793 62235
rect 13849 62179 13935 62235
rect 13991 62179 14077 62235
rect 14133 62179 14219 62235
rect 14275 62179 14361 62235
rect 14417 62179 14503 62235
rect 14559 62179 14645 62235
rect 14701 62179 14787 62235
rect 14843 62179 15000 62235
rect 0 62093 15000 62179
rect 0 62037 161 62093
rect 217 62037 303 62093
rect 359 62037 445 62093
rect 501 62037 587 62093
rect 643 62037 729 62093
rect 785 62037 871 62093
rect 927 62037 1013 62093
rect 1069 62037 1155 62093
rect 1211 62037 1297 62093
rect 1353 62037 1439 62093
rect 1495 62037 1581 62093
rect 1637 62037 1723 62093
rect 1779 62037 1865 62093
rect 1921 62037 2007 62093
rect 2063 62037 2149 62093
rect 2205 62037 2291 62093
rect 2347 62037 2433 62093
rect 2489 62037 2575 62093
rect 2631 62037 2717 62093
rect 2773 62037 2859 62093
rect 2915 62037 3001 62093
rect 3057 62037 3143 62093
rect 3199 62037 3285 62093
rect 3341 62037 3427 62093
rect 3483 62037 3569 62093
rect 3625 62037 3711 62093
rect 3767 62037 3853 62093
rect 3909 62037 3995 62093
rect 4051 62037 4137 62093
rect 4193 62037 4279 62093
rect 4335 62037 4421 62093
rect 4477 62037 4563 62093
rect 4619 62037 4705 62093
rect 4761 62037 4847 62093
rect 4903 62037 4989 62093
rect 5045 62037 5131 62093
rect 5187 62037 5273 62093
rect 5329 62037 5415 62093
rect 5471 62037 5557 62093
rect 5613 62037 5699 62093
rect 5755 62037 5841 62093
rect 5897 62037 5983 62093
rect 6039 62037 6125 62093
rect 6181 62037 6267 62093
rect 6323 62037 6409 62093
rect 6465 62037 6551 62093
rect 6607 62037 6693 62093
rect 6749 62037 6835 62093
rect 6891 62037 6977 62093
rect 7033 62037 7119 62093
rect 7175 62037 7261 62093
rect 7317 62037 7403 62093
rect 7459 62037 7545 62093
rect 7601 62037 7687 62093
rect 7743 62037 7829 62093
rect 7885 62037 7971 62093
rect 8027 62037 8113 62093
rect 8169 62037 8255 62093
rect 8311 62037 8397 62093
rect 8453 62037 8539 62093
rect 8595 62037 8681 62093
rect 8737 62037 8823 62093
rect 8879 62037 8965 62093
rect 9021 62037 9107 62093
rect 9163 62037 9249 62093
rect 9305 62037 9391 62093
rect 9447 62037 9533 62093
rect 9589 62037 9675 62093
rect 9731 62037 9817 62093
rect 9873 62037 9959 62093
rect 10015 62037 10101 62093
rect 10157 62037 10243 62093
rect 10299 62037 10385 62093
rect 10441 62037 10527 62093
rect 10583 62037 10669 62093
rect 10725 62037 10811 62093
rect 10867 62037 10953 62093
rect 11009 62037 11095 62093
rect 11151 62037 11237 62093
rect 11293 62037 11379 62093
rect 11435 62037 11521 62093
rect 11577 62037 11663 62093
rect 11719 62037 11805 62093
rect 11861 62037 11947 62093
rect 12003 62037 12089 62093
rect 12145 62037 12231 62093
rect 12287 62037 12373 62093
rect 12429 62037 12515 62093
rect 12571 62037 12657 62093
rect 12713 62037 12799 62093
rect 12855 62037 12941 62093
rect 12997 62037 13083 62093
rect 13139 62037 13225 62093
rect 13281 62037 13367 62093
rect 13423 62037 13509 62093
rect 13565 62037 13651 62093
rect 13707 62037 13793 62093
rect 13849 62037 13935 62093
rect 13991 62037 14077 62093
rect 14133 62037 14219 62093
rect 14275 62037 14361 62093
rect 14417 62037 14503 62093
rect 14559 62037 14645 62093
rect 14701 62037 14787 62093
rect 14843 62037 15000 62093
rect 0 62000 15000 62037
rect 0 61763 15000 61800
rect 0 61707 161 61763
rect 217 61707 303 61763
rect 359 61707 445 61763
rect 501 61707 587 61763
rect 643 61707 729 61763
rect 785 61707 871 61763
rect 927 61707 1013 61763
rect 1069 61707 1155 61763
rect 1211 61707 1297 61763
rect 1353 61707 1439 61763
rect 1495 61707 1581 61763
rect 1637 61707 1723 61763
rect 1779 61707 1865 61763
rect 1921 61707 2007 61763
rect 2063 61707 2149 61763
rect 2205 61707 2291 61763
rect 2347 61707 2433 61763
rect 2489 61707 2575 61763
rect 2631 61707 2717 61763
rect 2773 61707 2859 61763
rect 2915 61707 3001 61763
rect 3057 61707 3143 61763
rect 3199 61707 3285 61763
rect 3341 61707 3427 61763
rect 3483 61707 3569 61763
rect 3625 61707 3711 61763
rect 3767 61707 3853 61763
rect 3909 61707 3995 61763
rect 4051 61707 4137 61763
rect 4193 61707 4279 61763
rect 4335 61707 4421 61763
rect 4477 61707 4563 61763
rect 4619 61707 4705 61763
rect 4761 61707 4847 61763
rect 4903 61707 4989 61763
rect 5045 61707 5131 61763
rect 5187 61707 5273 61763
rect 5329 61707 5415 61763
rect 5471 61707 5557 61763
rect 5613 61707 5699 61763
rect 5755 61707 5841 61763
rect 5897 61707 5983 61763
rect 6039 61707 6125 61763
rect 6181 61707 6267 61763
rect 6323 61707 6409 61763
rect 6465 61707 6551 61763
rect 6607 61707 6693 61763
rect 6749 61707 6835 61763
rect 6891 61707 6977 61763
rect 7033 61707 7119 61763
rect 7175 61707 7261 61763
rect 7317 61707 7403 61763
rect 7459 61707 7545 61763
rect 7601 61707 7687 61763
rect 7743 61707 7829 61763
rect 7885 61707 7971 61763
rect 8027 61707 8113 61763
rect 8169 61707 8255 61763
rect 8311 61707 8397 61763
rect 8453 61707 8539 61763
rect 8595 61707 8681 61763
rect 8737 61707 8823 61763
rect 8879 61707 8965 61763
rect 9021 61707 9107 61763
rect 9163 61707 9249 61763
rect 9305 61707 9391 61763
rect 9447 61707 9533 61763
rect 9589 61707 9675 61763
rect 9731 61707 9817 61763
rect 9873 61707 9959 61763
rect 10015 61707 10101 61763
rect 10157 61707 10243 61763
rect 10299 61707 10385 61763
rect 10441 61707 10527 61763
rect 10583 61707 10669 61763
rect 10725 61707 10811 61763
rect 10867 61707 10953 61763
rect 11009 61707 11095 61763
rect 11151 61707 11237 61763
rect 11293 61707 11379 61763
rect 11435 61707 11521 61763
rect 11577 61707 11663 61763
rect 11719 61707 11805 61763
rect 11861 61707 11947 61763
rect 12003 61707 12089 61763
rect 12145 61707 12231 61763
rect 12287 61707 12373 61763
rect 12429 61707 12515 61763
rect 12571 61707 12657 61763
rect 12713 61707 12799 61763
rect 12855 61707 12941 61763
rect 12997 61707 13083 61763
rect 13139 61707 13225 61763
rect 13281 61707 13367 61763
rect 13423 61707 13509 61763
rect 13565 61707 13651 61763
rect 13707 61707 13793 61763
rect 13849 61707 13935 61763
rect 13991 61707 14077 61763
rect 14133 61707 14219 61763
rect 14275 61707 14361 61763
rect 14417 61707 14503 61763
rect 14559 61707 14645 61763
rect 14701 61707 14787 61763
rect 14843 61707 15000 61763
rect 0 61621 15000 61707
rect 0 61565 161 61621
rect 217 61565 303 61621
rect 359 61565 445 61621
rect 501 61565 587 61621
rect 643 61565 729 61621
rect 785 61565 871 61621
rect 927 61565 1013 61621
rect 1069 61565 1155 61621
rect 1211 61565 1297 61621
rect 1353 61565 1439 61621
rect 1495 61565 1581 61621
rect 1637 61565 1723 61621
rect 1779 61565 1865 61621
rect 1921 61565 2007 61621
rect 2063 61565 2149 61621
rect 2205 61565 2291 61621
rect 2347 61565 2433 61621
rect 2489 61565 2575 61621
rect 2631 61565 2717 61621
rect 2773 61565 2859 61621
rect 2915 61565 3001 61621
rect 3057 61565 3143 61621
rect 3199 61565 3285 61621
rect 3341 61565 3427 61621
rect 3483 61565 3569 61621
rect 3625 61565 3711 61621
rect 3767 61565 3853 61621
rect 3909 61565 3995 61621
rect 4051 61565 4137 61621
rect 4193 61565 4279 61621
rect 4335 61565 4421 61621
rect 4477 61565 4563 61621
rect 4619 61565 4705 61621
rect 4761 61565 4847 61621
rect 4903 61565 4989 61621
rect 5045 61565 5131 61621
rect 5187 61565 5273 61621
rect 5329 61565 5415 61621
rect 5471 61565 5557 61621
rect 5613 61565 5699 61621
rect 5755 61565 5841 61621
rect 5897 61565 5983 61621
rect 6039 61565 6125 61621
rect 6181 61565 6267 61621
rect 6323 61565 6409 61621
rect 6465 61565 6551 61621
rect 6607 61565 6693 61621
rect 6749 61565 6835 61621
rect 6891 61565 6977 61621
rect 7033 61565 7119 61621
rect 7175 61565 7261 61621
rect 7317 61565 7403 61621
rect 7459 61565 7545 61621
rect 7601 61565 7687 61621
rect 7743 61565 7829 61621
rect 7885 61565 7971 61621
rect 8027 61565 8113 61621
rect 8169 61565 8255 61621
rect 8311 61565 8397 61621
rect 8453 61565 8539 61621
rect 8595 61565 8681 61621
rect 8737 61565 8823 61621
rect 8879 61565 8965 61621
rect 9021 61565 9107 61621
rect 9163 61565 9249 61621
rect 9305 61565 9391 61621
rect 9447 61565 9533 61621
rect 9589 61565 9675 61621
rect 9731 61565 9817 61621
rect 9873 61565 9959 61621
rect 10015 61565 10101 61621
rect 10157 61565 10243 61621
rect 10299 61565 10385 61621
rect 10441 61565 10527 61621
rect 10583 61565 10669 61621
rect 10725 61565 10811 61621
rect 10867 61565 10953 61621
rect 11009 61565 11095 61621
rect 11151 61565 11237 61621
rect 11293 61565 11379 61621
rect 11435 61565 11521 61621
rect 11577 61565 11663 61621
rect 11719 61565 11805 61621
rect 11861 61565 11947 61621
rect 12003 61565 12089 61621
rect 12145 61565 12231 61621
rect 12287 61565 12373 61621
rect 12429 61565 12515 61621
rect 12571 61565 12657 61621
rect 12713 61565 12799 61621
rect 12855 61565 12941 61621
rect 12997 61565 13083 61621
rect 13139 61565 13225 61621
rect 13281 61565 13367 61621
rect 13423 61565 13509 61621
rect 13565 61565 13651 61621
rect 13707 61565 13793 61621
rect 13849 61565 13935 61621
rect 13991 61565 14077 61621
rect 14133 61565 14219 61621
rect 14275 61565 14361 61621
rect 14417 61565 14503 61621
rect 14559 61565 14645 61621
rect 14701 61565 14787 61621
rect 14843 61565 15000 61621
rect 0 61479 15000 61565
rect 0 61423 161 61479
rect 217 61423 303 61479
rect 359 61423 445 61479
rect 501 61423 587 61479
rect 643 61423 729 61479
rect 785 61423 871 61479
rect 927 61423 1013 61479
rect 1069 61423 1155 61479
rect 1211 61423 1297 61479
rect 1353 61423 1439 61479
rect 1495 61423 1581 61479
rect 1637 61423 1723 61479
rect 1779 61423 1865 61479
rect 1921 61423 2007 61479
rect 2063 61423 2149 61479
rect 2205 61423 2291 61479
rect 2347 61423 2433 61479
rect 2489 61423 2575 61479
rect 2631 61423 2717 61479
rect 2773 61423 2859 61479
rect 2915 61423 3001 61479
rect 3057 61423 3143 61479
rect 3199 61423 3285 61479
rect 3341 61423 3427 61479
rect 3483 61423 3569 61479
rect 3625 61423 3711 61479
rect 3767 61423 3853 61479
rect 3909 61423 3995 61479
rect 4051 61423 4137 61479
rect 4193 61423 4279 61479
rect 4335 61423 4421 61479
rect 4477 61423 4563 61479
rect 4619 61423 4705 61479
rect 4761 61423 4847 61479
rect 4903 61423 4989 61479
rect 5045 61423 5131 61479
rect 5187 61423 5273 61479
rect 5329 61423 5415 61479
rect 5471 61423 5557 61479
rect 5613 61423 5699 61479
rect 5755 61423 5841 61479
rect 5897 61423 5983 61479
rect 6039 61423 6125 61479
rect 6181 61423 6267 61479
rect 6323 61423 6409 61479
rect 6465 61423 6551 61479
rect 6607 61423 6693 61479
rect 6749 61423 6835 61479
rect 6891 61423 6977 61479
rect 7033 61423 7119 61479
rect 7175 61423 7261 61479
rect 7317 61423 7403 61479
rect 7459 61423 7545 61479
rect 7601 61423 7687 61479
rect 7743 61423 7829 61479
rect 7885 61423 7971 61479
rect 8027 61423 8113 61479
rect 8169 61423 8255 61479
rect 8311 61423 8397 61479
rect 8453 61423 8539 61479
rect 8595 61423 8681 61479
rect 8737 61423 8823 61479
rect 8879 61423 8965 61479
rect 9021 61423 9107 61479
rect 9163 61423 9249 61479
rect 9305 61423 9391 61479
rect 9447 61423 9533 61479
rect 9589 61423 9675 61479
rect 9731 61423 9817 61479
rect 9873 61423 9959 61479
rect 10015 61423 10101 61479
rect 10157 61423 10243 61479
rect 10299 61423 10385 61479
rect 10441 61423 10527 61479
rect 10583 61423 10669 61479
rect 10725 61423 10811 61479
rect 10867 61423 10953 61479
rect 11009 61423 11095 61479
rect 11151 61423 11237 61479
rect 11293 61423 11379 61479
rect 11435 61423 11521 61479
rect 11577 61423 11663 61479
rect 11719 61423 11805 61479
rect 11861 61423 11947 61479
rect 12003 61423 12089 61479
rect 12145 61423 12231 61479
rect 12287 61423 12373 61479
rect 12429 61423 12515 61479
rect 12571 61423 12657 61479
rect 12713 61423 12799 61479
rect 12855 61423 12941 61479
rect 12997 61423 13083 61479
rect 13139 61423 13225 61479
rect 13281 61423 13367 61479
rect 13423 61423 13509 61479
rect 13565 61423 13651 61479
rect 13707 61423 13793 61479
rect 13849 61423 13935 61479
rect 13991 61423 14077 61479
rect 14133 61423 14219 61479
rect 14275 61423 14361 61479
rect 14417 61423 14503 61479
rect 14559 61423 14645 61479
rect 14701 61423 14787 61479
rect 14843 61423 15000 61479
rect 0 61337 15000 61423
rect 0 61281 161 61337
rect 217 61281 303 61337
rect 359 61281 445 61337
rect 501 61281 587 61337
rect 643 61281 729 61337
rect 785 61281 871 61337
rect 927 61281 1013 61337
rect 1069 61281 1155 61337
rect 1211 61281 1297 61337
rect 1353 61281 1439 61337
rect 1495 61281 1581 61337
rect 1637 61281 1723 61337
rect 1779 61281 1865 61337
rect 1921 61281 2007 61337
rect 2063 61281 2149 61337
rect 2205 61281 2291 61337
rect 2347 61281 2433 61337
rect 2489 61281 2575 61337
rect 2631 61281 2717 61337
rect 2773 61281 2859 61337
rect 2915 61281 3001 61337
rect 3057 61281 3143 61337
rect 3199 61281 3285 61337
rect 3341 61281 3427 61337
rect 3483 61281 3569 61337
rect 3625 61281 3711 61337
rect 3767 61281 3853 61337
rect 3909 61281 3995 61337
rect 4051 61281 4137 61337
rect 4193 61281 4279 61337
rect 4335 61281 4421 61337
rect 4477 61281 4563 61337
rect 4619 61281 4705 61337
rect 4761 61281 4847 61337
rect 4903 61281 4989 61337
rect 5045 61281 5131 61337
rect 5187 61281 5273 61337
rect 5329 61281 5415 61337
rect 5471 61281 5557 61337
rect 5613 61281 5699 61337
rect 5755 61281 5841 61337
rect 5897 61281 5983 61337
rect 6039 61281 6125 61337
rect 6181 61281 6267 61337
rect 6323 61281 6409 61337
rect 6465 61281 6551 61337
rect 6607 61281 6693 61337
rect 6749 61281 6835 61337
rect 6891 61281 6977 61337
rect 7033 61281 7119 61337
rect 7175 61281 7261 61337
rect 7317 61281 7403 61337
rect 7459 61281 7545 61337
rect 7601 61281 7687 61337
rect 7743 61281 7829 61337
rect 7885 61281 7971 61337
rect 8027 61281 8113 61337
rect 8169 61281 8255 61337
rect 8311 61281 8397 61337
rect 8453 61281 8539 61337
rect 8595 61281 8681 61337
rect 8737 61281 8823 61337
rect 8879 61281 8965 61337
rect 9021 61281 9107 61337
rect 9163 61281 9249 61337
rect 9305 61281 9391 61337
rect 9447 61281 9533 61337
rect 9589 61281 9675 61337
rect 9731 61281 9817 61337
rect 9873 61281 9959 61337
rect 10015 61281 10101 61337
rect 10157 61281 10243 61337
rect 10299 61281 10385 61337
rect 10441 61281 10527 61337
rect 10583 61281 10669 61337
rect 10725 61281 10811 61337
rect 10867 61281 10953 61337
rect 11009 61281 11095 61337
rect 11151 61281 11237 61337
rect 11293 61281 11379 61337
rect 11435 61281 11521 61337
rect 11577 61281 11663 61337
rect 11719 61281 11805 61337
rect 11861 61281 11947 61337
rect 12003 61281 12089 61337
rect 12145 61281 12231 61337
rect 12287 61281 12373 61337
rect 12429 61281 12515 61337
rect 12571 61281 12657 61337
rect 12713 61281 12799 61337
rect 12855 61281 12941 61337
rect 12997 61281 13083 61337
rect 13139 61281 13225 61337
rect 13281 61281 13367 61337
rect 13423 61281 13509 61337
rect 13565 61281 13651 61337
rect 13707 61281 13793 61337
rect 13849 61281 13935 61337
rect 13991 61281 14077 61337
rect 14133 61281 14219 61337
rect 14275 61281 14361 61337
rect 14417 61281 14503 61337
rect 14559 61281 14645 61337
rect 14701 61281 14787 61337
rect 14843 61281 15000 61337
rect 0 61195 15000 61281
rect 0 61139 161 61195
rect 217 61139 303 61195
rect 359 61139 445 61195
rect 501 61139 587 61195
rect 643 61139 729 61195
rect 785 61139 871 61195
rect 927 61139 1013 61195
rect 1069 61139 1155 61195
rect 1211 61139 1297 61195
rect 1353 61139 1439 61195
rect 1495 61139 1581 61195
rect 1637 61139 1723 61195
rect 1779 61139 1865 61195
rect 1921 61139 2007 61195
rect 2063 61139 2149 61195
rect 2205 61139 2291 61195
rect 2347 61139 2433 61195
rect 2489 61139 2575 61195
rect 2631 61139 2717 61195
rect 2773 61139 2859 61195
rect 2915 61139 3001 61195
rect 3057 61139 3143 61195
rect 3199 61139 3285 61195
rect 3341 61139 3427 61195
rect 3483 61139 3569 61195
rect 3625 61139 3711 61195
rect 3767 61139 3853 61195
rect 3909 61139 3995 61195
rect 4051 61139 4137 61195
rect 4193 61139 4279 61195
rect 4335 61139 4421 61195
rect 4477 61139 4563 61195
rect 4619 61139 4705 61195
rect 4761 61139 4847 61195
rect 4903 61139 4989 61195
rect 5045 61139 5131 61195
rect 5187 61139 5273 61195
rect 5329 61139 5415 61195
rect 5471 61139 5557 61195
rect 5613 61139 5699 61195
rect 5755 61139 5841 61195
rect 5897 61139 5983 61195
rect 6039 61139 6125 61195
rect 6181 61139 6267 61195
rect 6323 61139 6409 61195
rect 6465 61139 6551 61195
rect 6607 61139 6693 61195
rect 6749 61139 6835 61195
rect 6891 61139 6977 61195
rect 7033 61139 7119 61195
rect 7175 61139 7261 61195
rect 7317 61139 7403 61195
rect 7459 61139 7545 61195
rect 7601 61139 7687 61195
rect 7743 61139 7829 61195
rect 7885 61139 7971 61195
rect 8027 61139 8113 61195
rect 8169 61139 8255 61195
rect 8311 61139 8397 61195
rect 8453 61139 8539 61195
rect 8595 61139 8681 61195
rect 8737 61139 8823 61195
rect 8879 61139 8965 61195
rect 9021 61139 9107 61195
rect 9163 61139 9249 61195
rect 9305 61139 9391 61195
rect 9447 61139 9533 61195
rect 9589 61139 9675 61195
rect 9731 61139 9817 61195
rect 9873 61139 9959 61195
rect 10015 61139 10101 61195
rect 10157 61139 10243 61195
rect 10299 61139 10385 61195
rect 10441 61139 10527 61195
rect 10583 61139 10669 61195
rect 10725 61139 10811 61195
rect 10867 61139 10953 61195
rect 11009 61139 11095 61195
rect 11151 61139 11237 61195
rect 11293 61139 11379 61195
rect 11435 61139 11521 61195
rect 11577 61139 11663 61195
rect 11719 61139 11805 61195
rect 11861 61139 11947 61195
rect 12003 61139 12089 61195
rect 12145 61139 12231 61195
rect 12287 61139 12373 61195
rect 12429 61139 12515 61195
rect 12571 61139 12657 61195
rect 12713 61139 12799 61195
rect 12855 61139 12941 61195
rect 12997 61139 13083 61195
rect 13139 61139 13225 61195
rect 13281 61139 13367 61195
rect 13423 61139 13509 61195
rect 13565 61139 13651 61195
rect 13707 61139 13793 61195
rect 13849 61139 13935 61195
rect 13991 61139 14077 61195
rect 14133 61139 14219 61195
rect 14275 61139 14361 61195
rect 14417 61139 14503 61195
rect 14559 61139 14645 61195
rect 14701 61139 14787 61195
rect 14843 61139 15000 61195
rect 0 61053 15000 61139
rect 0 60997 161 61053
rect 217 60997 303 61053
rect 359 60997 445 61053
rect 501 60997 587 61053
rect 643 60997 729 61053
rect 785 60997 871 61053
rect 927 60997 1013 61053
rect 1069 60997 1155 61053
rect 1211 60997 1297 61053
rect 1353 60997 1439 61053
rect 1495 60997 1581 61053
rect 1637 60997 1723 61053
rect 1779 60997 1865 61053
rect 1921 60997 2007 61053
rect 2063 60997 2149 61053
rect 2205 60997 2291 61053
rect 2347 60997 2433 61053
rect 2489 60997 2575 61053
rect 2631 60997 2717 61053
rect 2773 60997 2859 61053
rect 2915 60997 3001 61053
rect 3057 60997 3143 61053
rect 3199 60997 3285 61053
rect 3341 60997 3427 61053
rect 3483 60997 3569 61053
rect 3625 60997 3711 61053
rect 3767 60997 3853 61053
rect 3909 60997 3995 61053
rect 4051 60997 4137 61053
rect 4193 60997 4279 61053
rect 4335 60997 4421 61053
rect 4477 60997 4563 61053
rect 4619 60997 4705 61053
rect 4761 60997 4847 61053
rect 4903 60997 4989 61053
rect 5045 60997 5131 61053
rect 5187 60997 5273 61053
rect 5329 60997 5415 61053
rect 5471 60997 5557 61053
rect 5613 60997 5699 61053
rect 5755 60997 5841 61053
rect 5897 60997 5983 61053
rect 6039 60997 6125 61053
rect 6181 60997 6267 61053
rect 6323 60997 6409 61053
rect 6465 60997 6551 61053
rect 6607 60997 6693 61053
rect 6749 60997 6835 61053
rect 6891 60997 6977 61053
rect 7033 60997 7119 61053
rect 7175 60997 7261 61053
rect 7317 60997 7403 61053
rect 7459 60997 7545 61053
rect 7601 60997 7687 61053
rect 7743 60997 7829 61053
rect 7885 60997 7971 61053
rect 8027 60997 8113 61053
rect 8169 60997 8255 61053
rect 8311 60997 8397 61053
rect 8453 60997 8539 61053
rect 8595 60997 8681 61053
rect 8737 60997 8823 61053
rect 8879 60997 8965 61053
rect 9021 60997 9107 61053
rect 9163 60997 9249 61053
rect 9305 60997 9391 61053
rect 9447 60997 9533 61053
rect 9589 60997 9675 61053
rect 9731 60997 9817 61053
rect 9873 60997 9959 61053
rect 10015 60997 10101 61053
rect 10157 60997 10243 61053
rect 10299 60997 10385 61053
rect 10441 60997 10527 61053
rect 10583 60997 10669 61053
rect 10725 60997 10811 61053
rect 10867 60997 10953 61053
rect 11009 60997 11095 61053
rect 11151 60997 11237 61053
rect 11293 60997 11379 61053
rect 11435 60997 11521 61053
rect 11577 60997 11663 61053
rect 11719 60997 11805 61053
rect 11861 60997 11947 61053
rect 12003 60997 12089 61053
rect 12145 60997 12231 61053
rect 12287 60997 12373 61053
rect 12429 60997 12515 61053
rect 12571 60997 12657 61053
rect 12713 60997 12799 61053
rect 12855 60997 12941 61053
rect 12997 60997 13083 61053
rect 13139 60997 13225 61053
rect 13281 60997 13367 61053
rect 13423 60997 13509 61053
rect 13565 60997 13651 61053
rect 13707 60997 13793 61053
rect 13849 60997 13935 61053
rect 13991 60997 14077 61053
rect 14133 60997 14219 61053
rect 14275 60997 14361 61053
rect 14417 60997 14503 61053
rect 14559 60997 14645 61053
rect 14701 60997 14787 61053
rect 14843 60997 15000 61053
rect 0 60911 15000 60997
rect 0 60855 161 60911
rect 217 60855 303 60911
rect 359 60855 445 60911
rect 501 60855 587 60911
rect 643 60855 729 60911
rect 785 60855 871 60911
rect 927 60855 1013 60911
rect 1069 60855 1155 60911
rect 1211 60855 1297 60911
rect 1353 60855 1439 60911
rect 1495 60855 1581 60911
rect 1637 60855 1723 60911
rect 1779 60855 1865 60911
rect 1921 60855 2007 60911
rect 2063 60855 2149 60911
rect 2205 60855 2291 60911
rect 2347 60855 2433 60911
rect 2489 60855 2575 60911
rect 2631 60855 2717 60911
rect 2773 60855 2859 60911
rect 2915 60855 3001 60911
rect 3057 60855 3143 60911
rect 3199 60855 3285 60911
rect 3341 60855 3427 60911
rect 3483 60855 3569 60911
rect 3625 60855 3711 60911
rect 3767 60855 3853 60911
rect 3909 60855 3995 60911
rect 4051 60855 4137 60911
rect 4193 60855 4279 60911
rect 4335 60855 4421 60911
rect 4477 60855 4563 60911
rect 4619 60855 4705 60911
rect 4761 60855 4847 60911
rect 4903 60855 4989 60911
rect 5045 60855 5131 60911
rect 5187 60855 5273 60911
rect 5329 60855 5415 60911
rect 5471 60855 5557 60911
rect 5613 60855 5699 60911
rect 5755 60855 5841 60911
rect 5897 60855 5983 60911
rect 6039 60855 6125 60911
rect 6181 60855 6267 60911
rect 6323 60855 6409 60911
rect 6465 60855 6551 60911
rect 6607 60855 6693 60911
rect 6749 60855 6835 60911
rect 6891 60855 6977 60911
rect 7033 60855 7119 60911
rect 7175 60855 7261 60911
rect 7317 60855 7403 60911
rect 7459 60855 7545 60911
rect 7601 60855 7687 60911
rect 7743 60855 7829 60911
rect 7885 60855 7971 60911
rect 8027 60855 8113 60911
rect 8169 60855 8255 60911
rect 8311 60855 8397 60911
rect 8453 60855 8539 60911
rect 8595 60855 8681 60911
rect 8737 60855 8823 60911
rect 8879 60855 8965 60911
rect 9021 60855 9107 60911
rect 9163 60855 9249 60911
rect 9305 60855 9391 60911
rect 9447 60855 9533 60911
rect 9589 60855 9675 60911
rect 9731 60855 9817 60911
rect 9873 60855 9959 60911
rect 10015 60855 10101 60911
rect 10157 60855 10243 60911
rect 10299 60855 10385 60911
rect 10441 60855 10527 60911
rect 10583 60855 10669 60911
rect 10725 60855 10811 60911
rect 10867 60855 10953 60911
rect 11009 60855 11095 60911
rect 11151 60855 11237 60911
rect 11293 60855 11379 60911
rect 11435 60855 11521 60911
rect 11577 60855 11663 60911
rect 11719 60855 11805 60911
rect 11861 60855 11947 60911
rect 12003 60855 12089 60911
rect 12145 60855 12231 60911
rect 12287 60855 12373 60911
rect 12429 60855 12515 60911
rect 12571 60855 12657 60911
rect 12713 60855 12799 60911
rect 12855 60855 12941 60911
rect 12997 60855 13083 60911
rect 13139 60855 13225 60911
rect 13281 60855 13367 60911
rect 13423 60855 13509 60911
rect 13565 60855 13651 60911
rect 13707 60855 13793 60911
rect 13849 60855 13935 60911
rect 13991 60855 14077 60911
rect 14133 60855 14219 60911
rect 14275 60855 14361 60911
rect 14417 60855 14503 60911
rect 14559 60855 14645 60911
rect 14701 60855 14787 60911
rect 14843 60855 15000 60911
rect 0 60769 15000 60855
rect 0 60713 161 60769
rect 217 60713 303 60769
rect 359 60713 445 60769
rect 501 60713 587 60769
rect 643 60713 729 60769
rect 785 60713 871 60769
rect 927 60713 1013 60769
rect 1069 60713 1155 60769
rect 1211 60713 1297 60769
rect 1353 60713 1439 60769
rect 1495 60713 1581 60769
rect 1637 60713 1723 60769
rect 1779 60713 1865 60769
rect 1921 60713 2007 60769
rect 2063 60713 2149 60769
rect 2205 60713 2291 60769
rect 2347 60713 2433 60769
rect 2489 60713 2575 60769
rect 2631 60713 2717 60769
rect 2773 60713 2859 60769
rect 2915 60713 3001 60769
rect 3057 60713 3143 60769
rect 3199 60713 3285 60769
rect 3341 60713 3427 60769
rect 3483 60713 3569 60769
rect 3625 60713 3711 60769
rect 3767 60713 3853 60769
rect 3909 60713 3995 60769
rect 4051 60713 4137 60769
rect 4193 60713 4279 60769
rect 4335 60713 4421 60769
rect 4477 60713 4563 60769
rect 4619 60713 4705 60769
rect 4761 60713 4847 60769
rect 4903 60713 4989 60769
rect 5045 60713 5131 60769
rect 5187 60713 5273 60769
rect 5329 60713 5415 60769
rect 5471 60713 5557 60769
rect 5613 60713 5699 60769
rect 5755 60713 5841 60769
rect 5897 60713 5983 60769
rect 6039 60713 6125 60769
rect 6181 60713 6267 60769
rect 6323 60713 6409 60769
rect 6465 60713 6551 60769
rect 6607 60713 6693 60769
rect 6749 60713 6835 60769
rect 6891 60713 6977 60769
rect 7033 60713 7119 60769
rect 7175 60713 7261 60769
rect 7317 60713 7403 60769
rect 7459 60713 7545 60769
rect 7601 60713 7687 60769
rect 7743 60713 7829 60769
rect 7885 60713 7971 60769
rect 8027 60713 8113 60769
rect 8169 60713 8255 60769
rect 8311 60713 8397 60769
rect 8453 60713 8539 60769
rect 8595 60713 8681 60769
rect 8737 60713 8823 60769
rect 8879 60713 8965 60769
rect 9021 60713 9107 60769
rect 9163 60713 9249 60769
rect 9305 60713 9391 60769
rect 9447 60713 9533 60769
rect 9589 60713 9675 60769
rect 9731 60713 9817 60769
rect 9873 60713 9959 60769
rect 10015 60713 10101 60769
rect 10157 60713 10243 60769
rect 10299 60713 10385 60769
rect 10441 60713 10527 60769
rect 10583 60713 10669 60769
rect 10725 60713 10811 60769
rect 10867 60713 10953 60769
rect 11009 60713 11095 60769
rect 11151 60713 11237 60769
rect 11293 60713 11379 60769
rect 11435 60713 11521 60769
rect 11577 60713 11663 60769
rect 11719 60713 11805 60769
rect 11861 60713 11947 60769
rect 12003 60713 12089 60769
rect 12145 60713 12231 60769
rect 12287 60713 12373 60769
rect 12429 60713 12515 60769
rect 12571 60713 12657 60769
rect 12713 60713 12799 60769
rect 12855 60713 12941 60769
rect 12997 60713 13083 60769
rect 13139 60713 13225 60769
rect 13281 60713 13367 60769
rect 13423 60713 13509 60769
rect 13565 60713 13651 60769
rect 13707 60713 13793 60769
rect 13849 60713 13935 60769
rect 13991 60713 14077 60769
rect 14133 60713 14219 60769
rect 14275 60713 14361 60769
rect 14417 60713 14503 60769
rect 14559 60713 14645 60769
rect 14701 60713 14787 60769
rect 14843 60713 15000 60769
rect 0 60627 15000 60713
rect 0 60571 161 60627
rect 217 60571 303 60627
rect 359 60571 445 60627
rect 501 60571 587 60627
rect 643 60571 729 60627
rect 785 60571 871 60627
rect 927 60571 1013 60627
rect 1069 60571 1155 60627
rect 1211 60571 1297 60627
rect 1353 60571 1439 60627
rect 1495 60571 1581 60627
rect 1637 60571 1723 60627
rect 1779 60571 1865 60627
rect 1921 60571 2007 60627
rect 2063 60571 2149 60627
rect 2205 60571 2291 60627
rect 2347 60571 2433 60627
rect 2489 60571 2575 60627
rect 2631 60571 2717 60627
rect 2773 60571 2859 60627
rect 2915 60571 3001 60627
rect 3057 60571 3143 60627
rect 3199 60571 3285 60627
rect 3341 60571 3427 60627
rect 3483 60571 3569 60627
rect 3625 60571 3711 60627
rect 3767 60571 3853 60627
rect 3909 60571 3995 60627
rect 4051 60571 4137 60627
rect 4193 60571 4279 60627
rect 4335 60571 4421 60627
rect 4477 60571 4563 60627
rect 4619 60571 4705 60627
rect 4761 60571 4847 60627
rect 4903 60571 4989 60627
rect 5045 60571 5131 60627
rect 5187 60571 5273 60627
rect 5329 60571 5415 60627
rect 5471 60571 5557 60627
rect 5613 60571 5699 60627
rect 5755 60571 5841 60627
rect 5897 60571 5983 60627
rect 6039 60571 6125 60627
rect 6181 60571 6267 60627
rect 6323 60571 6409 60627
rect 6465 60571 6551 60627
rect 6607 60571 6693 60627
rect 6749 60571 6835 60627
rect 6891 60571 6977 60627
rect 7033 60571 7119 60627
rect 7175 60571 7261 60627
rect 7317 60571 7403 60627
rect 7459 60571 7545 60627
rect 7601 60571 7687 60627
rect 7743 60571 7829 60627
rect 7885 60571 7971 60627
rect 8027 60571 8113 60627
rect 8169 60571 8255 60627
rect 8311 60571 8397 60627
rect 8453 60571 8539 60627
rect 8595 60571 8681 60627
rect 8737 60571 8823 60627
rect 8879 60571 8965 60627
rect 9021 60571 9107 60627
rect 9163 60571 9249 60627
rect 9305 60571 9391 60627
rect 9447 60571 9533 60627
rect 9589 60571 9675 60627
rect 9731 60571 9817 60627
rect 9873 60571 9959 60627
rect 10015 60571 10101 60627
rect 10157 60571 10243 60627
rect 10299 60571 10385 60627
rect 10441 60571 10527 60627
rect 10583 60571 10669 60627
rect 10725 60571 10811 60627
rect 10867 60571 10953 60627
rect 11009 60571 11095 60627
rect 11151 60571 11237 60627
rect 11293 60571 11379 60627
rect 11435 60571 11521 60627
rect 11577 60571 11663 60627
rect 11719 60571 11805 60627
rect 11861 60571 11947 60627
rect 12003 60571 12089 60627
rect 12145 60571 12231 60627
rect 12287 60571 12373 60627
rect 12429 60571 12515 60627
rect 12571 60571 12657 60627
rect 12713 60571 12799 60627
rect 12855 60571 12941 60627
rect 12997 60571 13083 60627
rect 13139 60571 13225 60627
rect 13281 60571 13367 60627
rect 13423 60571 13509 60627
rect 13565 60571 13651 60627
rect 13707 60571 13793 60627
rect 13849 60571 13935 60627
rect 13991 60571 14077 60627
rect 14133 60571 14219 60627
rect 14275 60571 14361 60627
rect 14417 60571 14503 60627
rect 14559 60571 14645 60627
rect 14701 60571 14787 60627
rect 14843 60571 15000 60627
rect 0 60485 15000 60571
rect 0 60429 161 60485
rect 217 60429 303 60485
rect 359 60429 445 60485
rect 501 60429 587 60485
rect 643 60429 729 60485
rect 785 60429 871 60485
rect 927 60429 1013 60485
rect 1069 60429 1155 60485
rect 1211 60429 1297 60485
rect 1353 60429 1439 60485
rect 1495 60429 1581 60485
rect 1637 60429 1723 60485
rect 1779 60429 1865 60485
rect 1921 60429 2007 60485
rect 2063 60429 2149 60485
rect 2205 60429 2291 60485
rect 2347 60429 2433 60485
rect 2489 60429 2575 60485
rect 2631 60429 2717 60485
rect 2773 60429 2859 60485
rect 2915 60429 3001 60485
rect 3057 60429 3143 60485
rect 3199 60429 3285 60485
rect 3341 60429 3427 60485
rect 3483 60429 3569 60485
rect 3625 60429 3711 60485
rect 3767 60429 3853 60485
rect 3909 60429 3995 60485
rect 4051 60429 4137 60485
rect 4193 60429 4279 60485
rect 4335 60429 4421 60485
rect 4477 60429 4563 60485
rect 4619 60429 4705 60485
rect 4761 60429 4847 60485
rect 4903 60429 4989 60485
rect 5045 60429 5131 60485
rect 5187 60429 5273 60485
rect 5329 60429 5415 60485
rect 5471 60429 5557 60485
rect 5613 60429 5699 60485
rect 5755 60429 5841 60485
rect 5897 60429 5983 60485
rect 6039 60429 6125 60485
rect 6181 60429 6267 60485
rect 6323 60429 6409 60485
rect 6465 60429 6551 60485
rect 6607 60429 6693 60485
rect 6749 60429 6835 60485
rect 6891 60429 6977 60485
rect 7033 60429 7119 60485
rect 7175 60429 7261 60485
rect 7317 60429 7403 60485
rect 7459 60429 7545 60485
rect 7601 60429 7687 60485
rect 7743 60429 7829 60485
rect 7885 60429 7971 60485
rect 8027 60429 8113 60485
rect 8169 60429 8255 60485
rect 8311 60429 8397 60485
rect 8453 60429 8539 60485
rect 8595 60429 8681 60485
rect 8737 60429 8823 60485
rect 8879 60429 8965 60485
rect 9021 60429 9107 60485
rect 9163 60429 9249 60485
rect 9305 60429 9391 60485
rect 9447 60429 9533 60485
rect 9589 60429 9675 60485
rect 9731 60429 9817 60485
rect 9873 60429 9959 60485
rect 10015 60429 10101 60485
rect 10157 60429 10243 60485
rect 10299 60429 10385 60485
rect 10441 60429 10527 60485
rect 10583 60429 10669 60485
rect 10725 60429 10811 60485
rect 10867 60429 10953 60485
rect 11009 60429 11095 60485
rect 11151 60429 11237 60485
rect 11293 60429 11379 60485
rect 11435 60429 11521 60485
rect 11577 60429 11663 60485
rect 11719 60429 11805 60485
rect 11861 60429 11947 60485
rect 12003 60429 12089 60485
rect 12145 60429 12231 60485
rect 12287 60429 12373 60485
rect 12429 60429 12515 60485
rect 12571 60429 12657 60485
rect 12713 60429 12799 60485
rect 12855 60429 12941 60485
rect 12997 60429 13083 60485
rect 13139 60429 13225 60485
rect 13281 60429 13367 60485
rect 13423 60429 13509 60485
rect 13565 60429 13651 60485
rect 13707 60429 13793 60485
rect 13849 60429 13935 60485
rect 13991 60429 14077 60485
rect 14133 60429 14219 60485
rect 14275 60429 14361 60485
rect 14417 60429 14503 60485
rect 14559 60429 14645 60485
rect 14701 60429 14787 60485
rect 14843 60429 15000 60485
rect 0 60400 15000 60429
rect 0 60171 15000 60200
rect 0 60115 161 60171
rect 217 60115 303 60171
rect 359 60115 445 60171
rect 501 60115 587 60171
rect 643 60115 729 60171
rect 785 60115 871 60171
rect 927 60115 1013 60171
rect 1069 60115 1155 60171
rect 1211 60115 1297 60171
rect 1353 60115 1439 60171
rect 1495 60115 1581 60171
rect 1637 60115 1723 60171
rect 1779 60115 1865 60171
rect 1921 60115 2007 60171
rect 2063 60115 2149 60171
rect 2205 60115 2291 60171
rect 2347 60115 2433 60171
rect 2489 60115 2575 60171
rect 2631 60115 2717 60171
rect 2773 60115 2859 60171
rect 2915 60115 3001 60171
rect 3057 60115 3143 60171
rect 3199 60115 3285 60171
rect 3341 60115 3427 60171
rect 3483 60115 3569 60171
rect 3625 60115 3711 60171
rect 3767 60115 3853 60171
rect 3909 60115 3995 60171
rect 4051 60115 4137 60171
rect 4193 60115 4279 60171
rect 4335 60115 4421 60171
rect 4477 60115 4563 60171
rect 4619 60115 4705 60171
rect 4761 60115 4847 60171
rect 4903 60115 4989 60171
rect 5045 60115 5131 60171
rect 5187 60115 5273 60171
rect 5329 60115 5415 60171
rect 5471 60115 5557 60171
rect 5613 60115 5699 60171
rect 5755 60115 5841 60171
rect 5897 60115 5983 60171
rect 6039 60115 6125 60171
rect 6181 60115 6267 60171
rect 6323 60115 6409 60171
rect 6465 60115 6551 60171
rect 6607 60115 6693 60171
rect 6749 60115 6835 60171
rect 6891 60115 6977 60171
rect 7033 60115 7119 60171
rect 7175 60115 7261 60171
rect 7317 60115 7403 60171
rect 7459 60115 7545 60171
rect 7601 60115 7687 60171
rect 7743 60115 7829 60171
rect 7885 60115 7971 60171
rect 8027 60115 8113 60171
rect 8169 60115 8255 60171
rect 8311 60115 8397 60171
rect 8453 60115 8539 60171
rect 8595 60115 8681 60171
rect 8737 60115 8823 60171
rect 8879 60115 8965 60171
rect 9021 60115 9107 60171
rect 9163 60115 9249 60171
rect 9305 60115 9391 60171
rect 9447 60115 9533 60171
rect 9589 60115 9675 60171
rect 9731 60115 9817 60171
rect 9873 60115 9959 60171
rect 10015 60115 10101 60171
rect 10157 60115 10243 60171
rect 10299 60115 10385 60171
rect 10441 60115 10527 60171
rect 10583 60115 10669 60171
rect 10725 60115 10811 60171
rect 10867 60115 10953 60171
rect 11009 60115 11095 60171
rect 11151 60115 11237 60171
rect 11293 60115 11379 60171
rect 11435 60115 11521 60171
rect 11577 60115 11663 60171
rect 11719 60115 11805 60171
rect 11861 60115 11947 60171
rect 12003 60115 12089 60171
rect 12145 60115 12231 60171
rect 12287 60115 12373 60171
rect 12429 60115 12515 60171
rect 12571 60115 12657 60171
rect 12713 60115 12799 60171
rect 12855 60115 12941 60171
rect 12997 60115 13083 60171
rect 13139 60115 13225 60171
rect 13281 60115 13367 60171
rect 13423 60115 13509 60171
rect 13565 60115 13651 60171
rect 13707 60115 13793 60171
rect 13849 60115 13935 60171
rect 13991 60115 14077 60171
rect 14133 60115 14219 60171
rect 14275 60115 14361 60171
rect 14417 60115 14503 60171
rect 14559 60115 14645 60171
rect 14701 60115 14787 60171
rect 14843 60115 15000 60171
rect 0 60029 15000 60115
rect 0 59973 161 60029
rect 217 59973 303 60029
rect 359 59973 445 60029
rect 501 59973 587 60029
rect 643 59973 729 60029
rect 785 59973 871 60029
rect 927 59973 1013 60029
rect 1069 59973 1155 60029
rect 1211 59973 1297 60029
rect 1353 59973 1439 60029
rect 1495 59973 1581 60029
rect 1637 59973 1723 60029
rect 1779 59973 1865 60029
rect 1921 59973 2007 60029
rect 2063 59973 2149 60029
rect 2205 59973 2291 60029
rect 2347 59973 2433 60029
rect 2489 59973 2575 60029
rect 2631 59973 2717 60029
rect 2773 59973 2859 60029
rect 2915 59973 3001 60029
rect 3057 59973 3143 60029
rect 3199 59973 3285 60029
rect 3341 59973 3427 60029
rect 3483 59973 3569 60029
rect 3625 59973 3711 60029
rect 3767 59973 3853 60029
rect 3909 59973 3995 60029
rect 4051 59973 4137 60029
rect 4193 59973 4279 60029
rect 4335 59973 4421 60029
rect 4477 59973 4563 60029
rect 4619 59973 4705 60029
rect 4761 59973 4847 60029
rect 4903 59973 4989 60029
rect 5045 59973 5131 60029
rect 5187 59973 5273 60029
rect 5329 59973 5415 60029
rect 5471 59973 5557 60029
rect 5613 59973 5699 60029
rect 5755 59973 5841 60029
rect 5897 59973 5983 60029
rect 6039 59973 6125 60029
rect 6181 59973 6267 60029
rect 6323 59973 6409 60029
rect 6465 59973 6551 60029
rect 6607 59973 6693 60029
rect 6749 59973 6835 60029
rect 6891 59973 6977 60029
rect 7033 59973 7119 60029
rect 7175 59973 7261 60029
rect 7317 59973 7403 60029
rect 7459 59973 7545 60029
rect 7601 59973 7687 60029
rect 7743 59973 7829 60029
rect 7885 59973 7971 60029
rect 8027 59973 8113 60029
rect 8169 59973 8255 60029
rect 8311 59973 8397 60029
rect 8453 59973 8539 60029
rect 8595 59973 8681 60029
rect 8737 59973 8823 60029
rect 8879 59973 8965 60029
rect 9021 59973 9107 60029
rect 9163 59973 9249 60029
rect 9305 59973 9391 60029
rect 9447 59973 9533 60029
rect 9589 59973 9675 60029
rect 9731 59973 9817 60029
rect 9873 59973 9959 60029
rect 10015 59973 10101 60029
rect 10157 59973 10243 60029
rect 10299 59973 10385 60029
rect 10441 59973 10527 60029
rect 10583 59973 10669 60029
rect 10725 59973 10811 60029
rect 10867 59973 10953 60029
rect 11009 59973 11095 60029
rect 11151 59973 11237 60029
rect 11293 59973 11379 60029
rect 11435 59973 11521 60029
rect 11577 59973 11663 60029
rect 11719 59973 11805 60029
rect 11861 59973 11947 60029
rect 12003 59973 12089 60029
rect 12145 59973 12231 60029
rect 12287 59973 12373 60029
rect 12429 59973 12515 60029
rect 12571 59973 12657 60029
rect 12713 59973 12799 60029
rect 12855 59973 12941 60029
rect 12997 59973 13083 60029
rect 13139 59973 13225 60029
rect 13281 59973 13367 60029
rect 13423 59973 13509 60029
rect 13565 59973 13651 60029
rect 13707 59973 13793 60029
rect 13849 59973 13935 60029
rect 13991 59973 14077 60029
rect 14133 59973 14219 60029
rect 14275 59973 14361 60029
rect 14417 59973 14503 60029
rect 14559 59973 14645 60029
rect 14701 59973 14787 60029
rect 14843 59973 15000 60029
rect 0 59887 15000 59973
rect 0 59831 161 59887
rect 217 59831 303 59887
rect 359 59831 445 59887
rect 501 59831 587 59887
rect 643 59831 729 59887
rect 785 59831 871 59887
rect 927 59831 1013 59887
rect 1069 59831 1155 59887
rect 1211 59831 1297 59887
rect 1353 59831 1439 59887
rect 1495 59831 1581 59887
rect 1637 59831 1723 59887
rect 1779 59831 1865 59887
rect 1921 59831 2007 59887
rect 2063 59831 2149 59887
rect 2205 59831 2291 59887
rect 2347 59831 2433 59887
rect 2489 59831 2575 59887
rect 2631 59831 2717 59887
rect 2773 59831 2859 59887
rect 2915 59831 3001 59887
rect 3057 59831 3143 59887
rect 3199 59831 3285 59887
rect 3341 59831 3427 59887
rect 3483 59831 3569 59887
rect 3625 59831 3711 59887
rect 3767 59831 3853 59887
rect 3909 59831 3995 59887
rect 4051 59831 4137 59887
rect 4193 59831 4279 59887
rect 4335 59831 4421 59887
rect 4477 59831 4563 59887
rect 4619 59831 4705 59887
rect 4761 59831 4847 59887
rect 4903 59831 4989 59887
rect 5045 59831 5131 59887
rect 5187 59831 5273 59887
rect 5329 59831 5415 59887
rect 5471 59831 5557 59887
rect 5613 59831 5699 59887
rect 5755 59831 5841 59887
rect 5897 59831 5983 59887
rect 6039 59831 6125 59887
rect 6181 59831 6267 59887
rect 6323 59831 6409 59887
rect 6465 59831 6551 59887
rect 6607 59831 6693 59887
rect 6749 59831 6835 59887
rect 6891 59831 6977 59887
rect 7033 59831 7119 59887
rect 7175 59831 7261 59887
rect 7317 59831 7403 59887
rect 7459 59831 7545 59887
rect 7601 59831 7687 59887
rect 7743 59831 7829 59887
rect 7885 59831 7971 59887
rect 8027 59831 8113 59887
rect 8169 59831 8255 59887
rect 8311 59831 8397 59887
rect 8453 59831 8539 59887
rect 8595 59831 8681 59887
rect 8737 59831 8823 59887
rect 8879 59831 8965 59887
rect 9021 59831 9107 59887
rect 9163 59831 9249 59887
rect 9305 59831 9391 59887
rect 9447 59831 9533 59887
rect 9589 59831 9675 59887
rect 9731 59831 9817 59887
rect 9873 59831 9959 59887
rect 10015 59831 10101 59887
rect 10157 59831 10243 59887
rect 10299 59831 10385 59887
rect 10441 59831 10527 59887
rect 10583 59831 10669 59887
rect 10725 59831 10811 59887
rect 10867 59831 10953 59887
rect 11009 59831 11095 59887
rect 11151 59831 11237 59887
rect 11293 59831 11379 59887
rect 11435 59831 11521 59887
rect 11577 59831 11663 59887
rect 11719 59831 11805 59887
rect 11861 59831 11947 59887
rect 12003 59831 12089 59887
rect 12145 59831 12231 59887
rect 12287 59831 12373 59887
rect 12429 59831 12515 59887
rect 12571 59831 12657 59887
rect 12713 59831 12799 59887
rect 12855 59831 12941 59887
rect 12997 59831 13083 59887
rect 13139 59831 13225 59887
rect 13281 59831 13367 59887
rect 13423 59831 13509 59887
rect 13565 59831 13651 59887
rect 13707 59831 13793 59887
rect 13849 59831 13935 59887
rect 13991 59831 14077 59887
rect 14133 59831 14219 59887
rect 14275 59831 14361 59887
rect 14417 59831 14503 59887
rect 14559 59831 14645 59887
rect 14701 59831 14787 59887
rect 14843 59831 15000 59887
rect 0 59745 15000 59831
rect 0 59689 161 59745
rect 217 59689 303 59745
rect 359 59689 445 59745
rect 501 59689 587 59745
rect 643 59689 729 59745
rect 785 59689 871 59745
rect 927 59689 1013 59745
rect 1069 59689 1155 59745
rect 1211 59689 1297 59745
rect 1353 59689 1439 59745
rect 1495 59689 1581 59745
rect 1637 59689 1723 59745
rect 1779 59689 1865 59745
rect 1921 59689 2007 59745
rect 2063 59689 2149 59745
rect 2205 59689 2291 59745
rect 2347 59689 2433 59745
rect 2489 59689 2575 59745
rect 2631 59689 2717 59745
rect 2773 59689 2859 59745
rect 2915 59689 3001 59745
rect 3057 59689 3143 59745
rect 3199 59689 3285 59745
rect 3341 59689 3427 59745
rect 3483 59689 3569 59745
rect 3625 59689 3711 59745
rect 3767 59689 3853 59745
rect 3909 59689 3995 59745
rect 4051 59689 4137 59745
rect 4193 59689 4279 59745
rect 4335 59689 4421 59745
rect 4477 59689 4563 59745
rect 4619 59689 4705 59745
rect 4761 59689 4847 59745
rect 4903 59689 4989 59745
rect 5045 59689 5131 59745
rect 5187 59689 5273 59745
rect 5329 59689 5415 59745
rect 5471 59689 5557 59745
rect 5613 59689 5699 59745
rect 5755 59689 5841 59745
rect 5897 59689 5983 59745
rect 6039 59689 6125 59745
rect 6181 59689 6267 59745
rect 6323 59689 6409 59745
rect 6465 59689 6551 59745
rect 6607 59689 6693 59745
rect 6749 59689 6835 59745
rect 6891 59689 6977 59745
rect 7033 59689 7119 59745
rect 7175 59689 7261 59745
rect 7317 59689 7403 59745
rect 7459 59689 7545 59745
rect 7601 59689 7687 59745
rect 7743 59689 7829 59745
rect 7885 59689 7971 59745
rect 8027 59689 8113 59745
rect 8169 59689 8255 59745
rect 8311 59689 8397 59745
rect 8453 59689 8539 59745
rect 8595 59689 8681 59745
rect 8737 59689 8823 59745
rect 8879 59689 8965 59745
rect 9021 59689 9107 59745
rect 9163 59689 9249 59745
rect 9305 59689 9391 59745
rect 9447 59689 9533 59745
rect 9589 59689 9675 59745
rect 9731 59689 9817 59745
rect 9873 59689 9959 59745
rect 10015 59689 10101 59745
rect 10157 59689 10243 59745
rect 10299 59689 10385 59745
rect 10441 59689 10527 59745
rect 10583 59689 10669 59745
rect 10725 59689 10811 59745
rect 10867 59689 10953 59745
rect 11009 59689 11095 59745
rect 11151 59689 11237 59745
rect 11293 59689 11379 59745
rect 11435 59689 11521 59745
rect 11577 59689 11663 59745
rect 11719 59689 11805 59745
rect 11861 59689 11947 59745
rect 12003 59689 12089 59745
rect 12145 59689 12231 59745
rect 12287 59689 12373 59745
rect 12429 59689 12515 59745
rect 12571 59689 12657 59745
rect 12713 59689 12799 59745
rect 12855 59689 12941 59745
rect 12997 59689 13083 59745
rect 13139 59689 13225 59745
rect 13281 59689 13367 59745
rect 13423 59689 13509 59745
rect 13565 59689 13651 59745
rect 13707 59689 13793 59745
rect 13849 59689 13935 59745
rect 13991 59689 14077 59745
rect 14133 59689 14219 59745
rect 14275 59689 14361 59745
rect 14417 59689 14503 59745
rect 14559 59689 14645 59745
rect 14701 59689 14787 59745
rect 14843 59689 15000 59745
rect 0 59603 15000 59689
rect 0 59547 161 59603
rect 217 59547 303 59603
rect 359 59547 445 59603
rect 501 59547 587 59603
rect 643 59547 729 59603
rect 785 59547 871 59603
rect 927 59547 1013 59603
rect 1069 59547 1155 59603
rect 1211 59547 1297 59603
rect 1353 59547 1439 59603
rect 1495 59547 1581 59603
rect 1637 59547 1723 59603
rect 1779 59547 1865 59603
rect 1921 59547 2007 59603
rect 2063 59547 2149 59603
rect 2205 59547 2291 59603
rect 2347 59547 2433 59603
rect 2489 59547 2575 59603
rect 2631 59547 2717 59603
rect 2773 59547 2859 59603
rect 2915 59547 3001 59603
rect 3057 59547 3143 59603
rect 3199 59547 3285 59603
rect 3341 59547 3427 59603
rect 3483 59547 3569 59603
rect 3625 59547 3711 59603
rect 3767 59547 3853 59603
rect 3909 59547 3995 59603
rect 4051 59547 4137 59603
rect 4193 59547 4279 59603
rect 4335 59547 4421 59603
rect 4477 59547 4563 59603
rect 4619 59547 4705 59603
rect 4761 59547 4847 59603
rect 4903 59547 4989 59603
rect 5045 59547 5131 59603
rect 5187 59547 5273 59603
rect 5329 59547 5415 59603
rect 5471 59547 5557 59603
rect 5613 59547 5699 59603
rect 5755 59547 5841 59603
rect 5897 59547 5983 59603
rect 6039 59547 6125 59603
rect 6181 59547 6267 59603
rect 6323 59547 6409 59603
rect 6465 59547 6551 59603
rect 6607 59547 6693 59603
rect 6749 59547 6835 59603
rect 6891 59547 6977 59603
rect 7033 59547 7119 59603
rect 7175 59547 7261 59603
rect 7317 59547 7403 59603
rect 7459 59547 7545 59603
rect 7601 59547 7687 59603
rect 7743 59547 7829 59603
rect 7885 59547 7971 59603
rect 8027 59547 8113 59603
rect 8169 59547 8255 59603
rect 8311 59547 8397 59603
rect 8453 59547 8539 59603
rect 8595 59547 8681 59603
rect 8737 59547 8823 59603
rect 8879 59547 8965 59603
rect 9021 59547 9107 59603
rect 9163 59547 9249 59603
rect 9305 59547 9391 59603
rect 9447 59547 9533 59603
rect 9589 59547 9675 59603
rect 9731 59547 9817 59603
rect 9873 59547 9959 59603
rect 10015 59547 10101 59603
rect 10157 59547 10243 59603
rect 10299 59547 10385 59603
rect 10441 59547 10527 59603
rect 10583 59547 10669 59603
rect 10725 59547 10811 59603
rect 10867 59547 10953 59603
rect 11009 59547 11095 59603
rect 11151 59547 11237 59603
rect 11293 59547 11379 59603
rect 11435 59547 11521 59603
rect 11577 59547 11663 59603
rect 11719 59547 11805 59603
rect 11861 59547 11947 59603
rect 12003 59547 12089 59603
rect 12145 59547 12231 59603
rect 12287 59547 12373 59603
rect 12429 59547 12515 59603
rect 12571 59547 12657 59603
rect 12713 59547 12799 59603
rect 12855 59547 12941 59603
rect 12997 59547 13083 59603
rect 13139 59547 13225 59603
rect 13281 59547 13367 59603
rect 13423 59547 13509 59603
rect 13565 59547 13651 59603
rect 13707 59547 13793 59603
rect 13849 59547 13935 59603
rect 13991 59547 14077 59603
rect 14133 59547 14219 59603
rect 14275 59547 14361 59603
rect 14417 59547 14503 59603
rect 14559 59547 14645 59603
rect 14701 59547 14787 59603
rect 14843 59547 15000 59603
rect 0 59461 15000 59547
rect 0 59405 161 59461
rect 217 59405 303 59461
rect 359 59405 445 59461
rect 501 59405 587 59461
rect 643 59405 729 59461
rect 785 59405 871 59461
rect 927 59405 1013 59461
rect 1069 59405 1155 59461
rect 1211 59405 1297 59461
rect 1353 59405 1439 59461
rect 1495 59405 1581 59461
rect 1637 59405 1723 59461
rect 1779 59405 1865 59461
rect 1921 59405 2007 59461
rect 2063 59405 2149 59461
rect 2205 59405 2291 59461
rect 2347 59405 2433 59461
rect 2489 59405 2575 59461
rect 2631 59405 2717 59461
rect 2773 59405 2859 59461
rect 2915 59405 3001 59461
rect 3057 59405 3143 59461
rect 3199 59405 3285 59461
rect 3341 59405 3427 59461
rect 3483 59405 3569 59461
rect 3625 59405 3711 59461
rect 3767 59405 3853 59461
rect 3909 59405 3995 59461
rect 4051 59405 4137 59461
rect 4193 59405 4279 59461
rect 4335 59405 4421 59461
rect 4477 59405 4563 59461
rect 4619 59405 4705 59461
rect 4761 59405 4847 59461
rect 4903 59405 4989 59461
rect 5045 59405 5131 59461
rect 5187 59405 5273 59461
rect 5329 59405 5415 59461
rect 5471 59405 5557 59461
rect 5613 59405 5699 59461
rect 5755 59405 5841 59461
rect 5897 59405 5983 59461
rect 6039 59405 6125 59461
rect 6181 59405 6267 59461
rect 6323 59405 6409 59461
rect 6465 59405 6551 59461
rect 6607 59405 6693 59461
rect 6749 59405 6835 59461
rect 6891 59405 6977 59461
rect 7033 59405 7119 59461
rect 7175 59405 7261 59461
rect 7317 59405 7403 59461
rect 7459 59405 7545 59461
rect 7601 59405 7687 59461
rect 7743 59405 7829 59461
rect 7885 59405 7971 59461
rect 8027 59405 8113 59461
rect 8169 59405 8255 59461
rect 8311 59405 8397 59461
rect 8453 59405 8539 59461
rect 8595 59405 8681 59461
rect 8737 59405 8823 59461
rect 8879 59405 8965 59461
rect 9021 59405 9107 59461
rect 9163 59405 9249 59461
rect 9305 59405 9391 59461
rect 9447 59405 9533 59461
rect 9589 59405 9675 59461
rect 9731 59405 9817 59461
rect 9873 59405 9959 59461
rect 10015 59405 10101 59461
rect 10157 59405 10243 59461
rect 10299 59405 10385 59461
rect 10441 59405 10527 59461
rect 10583 59405 10669 59461
rect 10725 59405 10811 59461
rect 10867 59405 10953 59461
rect 11009 59405 11095 59461
rect 11151 59405 11237 59461
rect 11293 59405 11379 59461
rect 11435 59405 11521 59461
rect 11577 59405 11663 59461
rect 11719 59405 11805 59461
rect 11861 59405 11947 59461
rect 12003 59405 12089 59461
rect 12145 59405 12231 59461
rect 12287 59405 12373 59461
rect 12429 59405 12515 59461
rect 12571 59405 12657 59461
rect 12713 59405 12799 59461
rect 12855 59405 12941 59461
rect 12997 59405 13083 59461
rect 13139 59405 13225 59461
rect 13281 59405 13367 59461
rect 13423 59405 13509 59461
rect 13565 59405 13651 59461
rect 13707 59405 13793 59461
rect 13849 59405 13935 59461
rect 13991 59405 14077 59461
rect 14133 59405 14219 59461
rect 14275 59405 14361 59461
rect 14417 59405 14503 59461
rect 14559 59405 14645 59461
rect 14701 59405 14787 59461
rect 14843 59405 15000 59461
rect 0 59319 15000 59405
rect 0 59263 161 59319
rect 217 59263 303 59319
rect 359 59263 445 59319
rect 501 59263 587 59319
rect 643 59263 729 59319
rect 785 59263 871 59319
rect 927 59263 1013 59319
rect 1069 59263 1155 59319
rect 1211 59263 1297 59319
rect 1353 59263 1439 59319
rect 1495 59263 1581 59319
rect 1637 59263 1723 59319
rect 1779 59263 1865 59319
rect 1921 59263 2007 59319
rect 2063 59263 2149 59319
rect 2205 59263 2291 59319
rect 2347 59263 2433 59319
rect 2489 59263 2575 59319
rect 2631 59263 2717 59319
rect 2773 59263 2859 59319
rect 2915 59263 3001 59319
rect 3057 59263 3143 59319
rect 3199 59263 3285 59319
rect 3341 59263 3427 59319
rect 3483 59263 3569 59319
rect 3625 59263 3711 59319
rect 3767 59263 3853 59319
rect 3909 59263 3995 59319
rect 4051 59263 4137 59319
rect 4193 59263 4279 59319
rect 4335 59263 4421 59319
rect 4477 59263 4563 59319
rect 4619 59263 4705 59319
rect 4761 59263 4847 59319
rect 4903 59263 4989 59319
rect 5045 59263 5131 59319
rect 5187 59263 5273 59319
rect 5329 59263 5415 59319
rect 5471 59263 5557 59319
rect 5613 59263 5699 59319
rect 5755 59263 5841 59319
rect 5897 59263 5983 59319
rect 6039 59263 6125 59319
rect 6181 59263 6267 59319
rect 6323 59263 6409 59319
rect 6465 59263 6551 59319
rect 6607 59263 6693 59319
rect 6749 59263 6835 59319
rect 6891 59263 6977 59319
rect 7033 59263 7119 59319
rect 7175 59263 7261 59319
rect 7317 59263 7403 59319
rect 7459 59263 7545 59319
rect 7601 59263 7687 59319
rect 7743 59263 7829 59319
rect 7885 59263 7971 59319
rect 8027 59263 8113 59319
rect 8169 59263 8255 59319
rect 8311 59263 8397 59319
rect 8453 59263 8539 59319
rect 8595 59263 8681 59319
rect 8737 59263 8823 59319
rect 8879 59263 8965 59319
rect 9021 59263 9107 59319
rect 9163 59263 9249 59319
rect 9305 59263 9391 59319
rect 9447 59263 9533 59319
rect 9589 59263 9675 59319
rect 9731 59263 9817 59319
rect 9873 59263 9959 59319
rect 10015 59263 10101 59319
rect 10157 59263 10243 59319
rect 10299 59263 10385 59319
rect 10441 59263 10527 59319
rect 10583 59263 10669 59319
rect 10725 59263 10811 59319
rect 10867 59263 10953 59319
rect 11009 59263 11095 59319
rect 11151 59263 11237 59319
rect 11293 59263 11379 59319
rect 11435 59263 11521 59319
rect 11577 59263 11663 59319
rect 11719 59263 11805 59319
rect 11861 59263 11947 59319
rect 12003 59263 12089 59319
rect 12145 59263 12231 59319
rect 12287 59263 12373 59319
rect 12429 59263 12515 59319
rect 12571 59263 12657 59319
rect 12713 59263 12799 59319
rect 12855 59263 12941 59319
rect 12997 59263 13083 59319
rect 13139 59263 13225 59319
rect 13281 59263 13367 59319
rect 13423 59263 13509 59319
rect 13565 59263 13651 59319
rect 13707 59263 13793 59319
rect 13849 59263 13935 59319
rect 13991 59263 14077 59319
rect 14133 59263 14219 59319
rect 14275 59263 14361 59319
rect 14417 59263 14503 59319
rect 14559 59263 14645 59319
rect 14701 59263 14787 59319
rect 14843 59263 15000 59319
rect 0 59177 15000 59263
rect 0 59121 161 59177
rect 217 59121 303 59177
rect 359 59121 445 59177
rect 501 59121 587 59177
rect 643 59121 729 59177
rect 785 59121 871 59177
rect 927 59121 1013 59177
rect 1069 59121 1155 59177
rect 1211 59121 1297 59177
rect 1353 59121 1439 59177
rect 1495 59121 1581 59177
rect 1637 59121 1723 59177
rect 1779 59121 1865 59177
rect 1921 59121 2007 59177
rect 2063 59121 2149 59177
rect 2205 59121 2291 59177
rect 2347 59121 2433 59177
rect 2489 59121 2575 59177
rect 2631 59121 2717 59177
rect 2773 59121 2859 59177
rect 2915 59121 3001 59177
rect 3057 59121 3143 59177
rect 3199 59121 3285 59177
rect 3341 59121 3427 59177
rect 3483 59121 3569 59177
rect 3625 59121 3711 59177
rect 3767 59121 3853 59177
rect 3909 59121 3995 59177
rect 4051 59121 4137 59177
rect 4193 59121 4279 59177
rect 4335 59121 4421 59177
rect 4477 59121 4563 59177
rect 4619 59121 4705 59177
rect 4761 59121 4847 59177
rect 4903 59121 4989 59177
rect 5045 59121 5131 59177
rect 5187 59121 5273 59177
rect 5329 59121 5415 59177
rect 5471 59121 5557 59177
rect 5613 59121 5699 59177
rect 5755 59121 5841 59177
rect 5897 59121 5983 59177
rect 6039 59121 6125 59177
rect 6181 59121 6267 59177
rect 6323 59121 6409 59177
rect 6465 59121 6551 59177
rect 6607 59121 6693 59177
rect 6749 59121 6835 59177
rect 6891 59121 6977 59177
rect 7033 59121 7119 59177
rect 7175 59121 7261 59177
rect 7317 59121 7403 59177
rect 7459 59121 7545 59177
rect 7601 59121 7687 59177
rect 7743 59121 7829 59177
rect 7885 59121 7971 59177
rect 8027 59121 8113 59177
rect 8169 59121 8255 59177
rect 8311 59121 8397 59177
rect 8453 59121 8539 59177
rect 8595 59121 8681 59177
rect 8737 59121 8823 59177
rect 8879 59121 8965 59177
rect 9021 59121 9107 59177
rect 9163 59121 9249 59177
rect 9305 59121 9391 59177
rect 9447 59121 9533 59177
rect 9589 59121 9675 59177
rect 9731 59121 9817 59177
rect 9873 59121 9959 59177
rect 10015 59121 10101 59177
rect 10157 59121 10243 59177
rect 10299 59121 10385 59177
rect 10441 59121 10527 59177
rect 10583 59121 10669 59177
rect 10725 59121 10811 59177
rect 10867 59121 10953 59177
rect 11009 59121 11095 59177
rect 11151 59121 11237 59177
rect 11293 59121 11379 59177
rect 11435 59121 11521 59177
rect 11577 59121 11663 59177
rect 11719 59121 11805 59177
rect 11861 59121 11947 59177
rect 12003 59121 12089 59177
rect 12145 59121 12231 59177
rect 12287 59121 12373 59177
rect 12429 59121 12515 59177
rect 12571 59121 12657 59177
rect 12713 59121 12799 59177
rect 12855 59121 12941 59177
rect 12997 59121 13083 59177
rect 13139 59121 13225 59177
rect 13281 59121 13367 59177
rect 13423 59121 13509 59177
rect 13565 59121 13651 59177
rect 13707 59121 13793 59177
rect 13849 59121 13935 59177
rect 13991 59121 14077 59177
rect 14133 59121 14219 59177
rect 14275 59121 14361 59177
rect 14417 59121 14503 59177
rect 14559 59121 14645 59177
rect 14701 59121 14787 59177
rect 14843 59121 15000 59177
rect 0 59035 15000 59121
rect 0 58979 161 59035
rect 217 58979 303 59035
rect 359 58979 445 59035
rect 501 58979 587 59035
rect 643 58979 729 59035
rect 785 58979 871 59035
rect 927 58979 1013 59035
rect 1069 58979 1155 59035
rect 1211 58979 1297 59035
rect 1353 58979 1439 59035
rect 1495 58979 1581 59035
rect 1637 58979 1723 59035
rect 1779 58979 1865 59035
rect 1921 58979 2007 59035
rect 2063 58979 2149 59035
rect 2205 58979 2291 59035
rect 2347 58979 2433 59035
rect 2489 58979 2575 59035
rect 2631 58979 2717 59035
rect 2773 58979 2859 59035
rect 2915 58979 3001 59035
rect 3057 58979 3143 59035
rect 3199 58979 3285 59035
rect 3341 58979 3427 59035
rect 3483 58979 3569 59035
rect 3625 58979 3711 59035
rect 3767 58979 3853 59035
rect 3909 58979 3995 59035
rect 4051 58979 4137 59035
rect 4193 58979 4279 59035
rect 4335 58979 4421 59035
rect 4477 58979 4563 59035
rect 4619 58979 4705 59035
rect 4761 58979 4847 59035
rect 4903 58979 4989 59035
rect 5045 58979 5131 59035
rect 5187 58979 5273 59035
rect 5329 58979 5415 59035
rect 5471 58979 5557 59035
rect 5613 58979 5699 59035
rect 5755 58979 5841 59035
rect 5897 58979 5983 59035
rect 6039 58979 6125 59035
rect 6181 58979 6267 59035
rect 6323 58979 6409 59035
rect 6465 58979 6551 59035
rect 6607 58979 6693 59035
rect 6749 58979 6835 59035
rect 6891 58979 6977 59035
rect 7033 58979 7119 59035
rect 7175 58979 7261 59035
rect 7317 58979 7403 59035
rect 7459 58979 7545 59035
rect 7601 58979 7687 59035
rect 7743 58979 7829 59035
rect 7885 58979 7971 59035
rect 8027 58979 8113 59035
rect 8169 58979 8255 59035
rect 8311 58979 8397 59035
rect 8453 58979 8539 59035
rect 8595 58979 8681 59035
rect 8737 58979 8823 59035
rect 8879 58979 8965 59035
rect 9021 58979 9107 59035
rect 9163 58979 9249 59035
rect 9305 58979 9391 59035
rect 9447 58979 9533 59035
rect 9589 58979 9675 59035
rect 9731 58979 9817 59035
rect 9873 58979 9959 59035
rect 10015 58979 10101 59035
rect 10157 58979 10243 59035
rect 10299 58979 10385 59035
rect 10441 58979 10527 59035
rect 10583 58979 10669 59035
rect 10725 58979 10811 59035
rect 10867 58979 10953 59035
rect 11009 58979 11095 59035
rect 11151 58979 11237 59035
rect 11293 58979 11379 59035
rect 11435 58979 11521 59035
rect 11577 58979 11663 59035
rect 11719 58979 11805 59035
rect 11861 58979 11947 59035
rect 12003 58979 12089 59035
rect 12145 58979 12231 59035
rect 12287 58979 12373 59035
rect 12429 58979 12515 59035
rect 12571 58979 12657 59035
rect 12713 58979 12799 59035
rect 12855 58979 12941 59035
rect 12997 58979 13083 59035
rect 13139 58979 13225 59035
rect 13281 58979 13367 59035
rect 13423 58979 13509 59035
rect 13565 58979 13651 59035
rect 13707 58979 13793 59035
rect 13849 58979 13935 59035
rect 13991 58979 14077 59035
rect 14133 58979 14219 59035
rect 14275 58979 14361 59035
rect 14417 58979 14503 59035
rect 14559 58979 14645 59035
rect 14701 58979 14787 59035
rect 14843 58979 15000 59035
rect 0 58893 15000 58979
rect 0 58837 161 58893
rect 217 58837 303 58893
rect 359 58837 445 58893
rect 501 58837 587 58893
rect 643 58837 729 58893
rect 785 58837 871 58893
rect 927 58837 1013 58893
rect 1069 58837 1155 58893
rect 1211 58837 1297 58893
rect 1353 58837 1439 58893
rect 1495 58837 1581 58893
rect 1637 58837 1723 58893
rect 1779 58837 1865 58893
rect 1921 58837 2007 58893
rect 2063 58837 2149 58893
rect 2205 58837 2291 58893
rect 2347 58837 2433 58893
rect 2489 58837 2575 58893
rect 2631 58837 2717 58893
rect 2773 58837 2859 58893
rect 2915 58837 3001 58893
rect 3057 58837 3143 58893
rect 3199 58837 3285 58893
rect 3341 58837 3427 58893
rect 3483 58837 3569 58893
rect 3625 58837 3711 58893
rect 3767 58837 3853 58893
rect 3909 58837 3995 58893
rect 4051 58837 4137 58893
rect 4193 58837 4279 58893
rect 4335 58837 4421 58893
rect 4477 58837 4563 58893
rect 4619 58837 4705 58893
rect 4761 58837 4847 58893
rect 4903 58837 4989 58893
rect 5045 58837 5131 58893
rect 5187 58837 5273 58893
rect 5329 58837 5415 58893
rect 5471 58837 5557 58893
rect 5613 58837 5699 58893
rect 5755 58837 5841 58893
rect 5897 58837 5983 58893
rect 6039 58837 6125 58893
rect 6181 58837 6267 58893
rect 6323 58837 6409 58893
rect 6465 58837 6551 58893
rect 6607 58837 6693 58893
rect 6749 58837 6835 58893
rect 6891 58837 6977 58893
rect 7033 58837 7119 58893
rect 7175 58837 7261 58893
rect 7317 58837 7403 58893
rect 7459 58837 7545 58893
rect 7601 58837 7687 58893
rect 7743 58837 7829 58893
rect 7885 58837 7971 58893
rect 8027 58837 8113 58893
rect 8169 58837 8255 58893
rect 8311 58837 8397 58893
rect 8453 58837 8539 58893
rect 8595 58837 8681 58893
rect 8737 58837 8823 58893
rect 8879 58837 8965 58893
rect 9021 58837 9107 58893
rect 9163 58837 9249 58893
rect 9305 58837 9391 58893
rect 9447 58837 9533 58893
rect 9589 58837 9675 58893
rect 9731 58837 9817 58893
rect 9873 58837 9959 58893
rect 10015 58837 10101 58893
rect 10157 58837 10243 58893
rect 10299 58837 10385 58893
rect 10441 58837 10527 58893
rect 10583 58837 10669 58893
rect 10725 58837 10811 58893
rect 10867 58837 10953 58893
rect 11009 58837 11095 58893
rect 11151 58837 11237 58893
rect 11293 58837 11379 58893
rect 11435 58837 11521 58893
rect 11577 58837 11663 58893
rect 11719 58837 11805 58893
rect 11861 58837 11947 58893
rect 12003 58837 12089 58893
rect 12145 58837 12231 58893
rect 12287 58837 12373 58893
rect 12429 58837 12515 58893
rect 12571 58837 12657 58893
rect 12713 58837 12799 58893
rect 12855 58837 12941 58893
rect 12997 58837 13083 58893
rect 13139 58837 13225 58893
rect 13281 58837 13367 58893
rect 13423 58837 13509 58893
rect 13565 58837 13651 58893
rect 13707 58837 13793 58893
rect 13849 58837 13935 58893
rect 13991 58837 14077 58893
rect 14133 58837 14219 58893
rect 14275 58837 14361 58893
rect 14417 58837 14503 58893
rect 14559 58837 14645 58893
rect 14701 58837 14787 58893
rect 14843 58837 15000 58893
rect 0 58800 15000 58837
rect 0 58563 15000 58600
rect 0 58507 161 58563
rect 217 58507 303 58563
rect 359 58507 445 58563
rect 501 58507 587 58563
rect 643 58507 729 58563
rect 785 58507 871 58563
rect 927 58507 1013 58563
rect 1069 58507 1155 58563
rect 1211 58507 1297 58563
rect 1353 58507 1439 58563
rect 1495 58507 1581 58563
rect 1637 58507 1723 58563
rect 1779 58507 1865 58563
rect 1921 58507 2007 58563
rect 2063 58507 2149 58563
rect 2205 58507 2291 58563
rect 2347 58507 2433 58563
rect 2489 58507 2575 58563
rect 2631 58507 2717 58563
rect 2773 58507 2859 58563
rect 2915 58507 3001 58563
rect 3057 58507 3143 58563
rect 3199 58507 3285 58563
rect 3341 58507 3427 58563
rect 3483 58507 3569 58563
rect 3625 58507 3711 58563
rect 3767 58507 3853 58563
rect 3909 58507 3995 58563
rect 4051 58507 4137 58563
rect 4193 58507 4279 58563
rect 4335 58507 4421 58563
rect 4477 58507 4563 58563
rect 4619 58507 4705 58563
rect 4761 58507 4847 58563
rect 4903 58507 4989 58563
rect 5045 58507 5131 58563
rect 5187 58507 5273 58563
rect 5329 58507 5415 58563
rect 5471 58507 5557 58563
rect 5613 58507 5699 58563
rect 5755 58507 5841 58563
rect 5897 58507 5983 58563
rect 6039 58507 6125 58563
rect 6181 58507 6267 58563
rect 6323 58507 6409 58563
rect 6465 58507 6551 58563
rect 6607 58507 6693 58563
rect 6749 58507 6835 58563
rect 6891 58507 6977 58563
rect 7033 58507 7119 58563
rect 7175 58507 7261 58563
rect 7317 58507 7403 58563
rect 7459 58507 7545 58563
rect 7601 58507 7687 58563
rect 7743 58507 7829 58563
rect 7885 58507 7971 58563
rect 8027 58507 8113 58563
rect 8169 58507 8255 58563
rect 8311 58507 8397 58563
rect 8453 58507 8539 58563
rect 8595 58507 8681 58563
rect 8737 58507 8823 58563
rect 8879 58507 8965 58563
rect 9021 58507 9107 58563
rect 9163 58507 9249 58563
rect 9305 58507 9391 58563
rect 9447 58507 9533 58563
rect 9589 58507 9675 58563
rect 9731 58507 9817 58563
rect 9873 58507 9959 58563
rect 10015 58507 10101 58563
rect 10157 58507 10243 58563
rect 10299 58507 10385 58563
rect 10441 58507 10527 58563
rect 10583 58507 10669 58563
rect 10725 58507 10811 58563
rect 10867 58507 10953 58563
rect 11009 58507 11095 58563
rect 11151 58507 11237 58563
rect 11293 58507 11379 58563
rect 11435 58507 11521 58563
rect 11577 58507 11663 58563
rect 11719 58507 11805 58563
rect 11861 58507 11947 58563
rect 12003 58507 12089 58563
rect 12145 58507 12231 58563
rect 12287 58507 12373 58563
rect 12429 58507 12515 58563
rect 12571 58507 12657 58563
rect 12713 58507 12799 58563
rect 12855 58507 12941 58563
rect 12997 58507 13083 58563
rect 13139 58507 13225 58563
rect 13281 58507 13367 58563
rect 13423 58507 13509 58563
rect 13565 58507 13651 58563
rect 13707 58507 13793 58563
rect 13849 58507 13935 58563
rect 13991 58507 14077 58563
rect 14133 58507 14219 58563
rect 14275 58507 14361 58563
rect 14417 58507 14503 58563
rect 14559 58507 14645 58563
rect 14701 58507 14787 58563
rect 14843 58507 15000 58563
rect 0 58421 15000 58507
rect 0 58365 161 58421
rect 217 58365 303 58421
rect 359 58365 445 58421
rect 501 58365 587 58421
rect 643 58365 729 58421
rect 785 58365 871 58421
rect 927 58365 1013 58421
rect 1069 58365 1155 58421
rect 1211 58365 1297 58421
rect 1353 58365 1439 58421
rect 1495 58365 1581 58421
rect 1637 58365 1723 58421
rect 1779 58365 1865 58421
rect 1921 58365 2007 58421
rect 2063 58365 2149 58421
rect 2205 58365 2291 58421
rect 2347 58365 2433 58421
rect 2489 58365 2575 58421
rect 2631 58365 2717 58421
rect 2773 58365 2859 58421
rect 2915 58365 3001 58421
rect 3057 58365 3143 58421
rect 3199 58365 3285 58421
rect 3341 58365 3427 58421
rect 3483 58365 3569 58421
rect 3625 58365 3711 58421
rect 3767 58365 3853 58421
rect 3909 58365 3995 58421
rect 4051 58365 4137 58421
rect 4193 58365 4279 58421
rect 4335 58365 4421 58421
rect 4477 58365 4563 58421
rect 4619 58365 4705 58421
rect 4761 58365 4847 58421
rect 4903 58365 4989 58421
rect 5045 58365 5131 58421
rect 5187 58365 5273 58421
rect 5329 58365 5415 58421
rect 5471 58365 5557 58421
rect 5613 58365 5699 58421
rect 5755 58365 5841 58421
rect 5897 58365 5983 58421
rect 6039 58365 6125 58421
rect 6181 58365 6267 58421
rect 6323 58365 6409 58421
rect 6465 58365 6551 58421
rect 6607 58365 6693 58421
rect 6749 58365 6835 58421
rect 6891 58365 6977 58421
rect 7033 58365 7119 58421
rect 7175 58365 7261 58421
rect 7317 58365 7403 58421
rect 7459 58365 7545 58421
rect 7601 58365 7687 58421
rect 7743 58365 7829 58421
rect 7885 58365 7971 58421
rect 8027 58365 8113 58421
rect 8169 58365 8255 58421
rect 8311 58365 8397 58421
rect 8453 58365 8539 58421
rect 8595 58365 8681 58421
rect 8737 58365 8823 58421
rect 8879 58365 8965 58421
rect 9021 58365 9107 58421
rect 9163 58365 9249 58421
rect 9305 58365 9391 58421
rect 9447 58365 9533 58421
rect 9589 58365 9675 58421
rect 9731 58365 9817 58421
rect 9873 58365 9959 58421
rect 10015 58365 10101 58421
rect 10157 58365 10243 58421
rect 10299 58365 10385 58421
rect 10441 58365 10527 58421
rect 10583 58365 10669 58421
rect 10725 58365 10811 58421
rect 10867 58365 10953 58421
rect 11009 58365 11095 58421
rect 11151 58365 11237 58421
rect 11293 58365 11379 58421
rect 11435 58365 11521 58421
rect 11577 58365 11663 58421
rect 11719 58365 11805 58421
rect 11861 58365 11947 58421
rect 12003 58365 12089 58421
rect 12145 58365 12231 58421
rect 12287 58365 12373 58421
rect 12429 58365 12515 58421
rect 12571 58365 12657 58421
rect 12713 58365 12799 58421
rect 12855 58365 12941 58421
rect 12997 58365 13083 58421
rect 13139 58365 13225 58421
rect 13281 58365 13367 58421
rect 13423 58365 13509 58421
rect 13565 58365 13651 58421
rect 13707 58365 13793 58421
rect 13849 58365 13935 58421
rect 13991 58365 14077 58421
rect 14133 58365 14219 58421
rect 14275 58365 14361 58421
rect 14417 58365 14503 58421
rect 14559 58365 14645 58421
rect 14701 58365 14787 58421
rect 14843 58365 15000 58421
rect 0 58279 15000 58365
rect 0 58223 161 58279
rect 217 58223 303 58279
rect 359 58223 445 58279
rect 501 58223 587 58279
rect 643 58223 729 58279
rect 785 58223 871 58279
rect 927 58223 1013 58279
rect 1069 58223 1155 58279
rect 1211 58223 1297 58279
rect 1353 58223 1439 58279
rect 1495 58223 1581 58279
rect 1637 58223 1723 58279
rect 1779 58223 1865 58279
rect 1921 58223 2007 58279
rect 2063 58223 2149 58279
rect 2205 58223 2291 58279
rect 2347 58223 2433 58279
rect 2489 58223 2575 58279
rect 2631 58223 2717 58279
rect 2773 58223 2859 58279
rect 2915 58223 3001 58279
rect 3057 58223 3143 58279
rect 3199 58223 3285 58279
rect 3341 58223 3427 58279
rect 3483 58223 3569 58279
rect 3625 58223 3711 58279
rect 3767 58223 3853 58279
rect 3909 58223 3995 58279
rect 4051 58223 4137 58279
rect 4193 58223 4279 58279
rect 4335 58223 4421 58279
rect 4477 58223 4563 58279
rect 4619 58223 4705 58279
rect 4761 58223 4847 58279
rect 4903 58223 4989 58279
rect 5045 58223 5131 58279
rect 5187 58223 5273 58279
rect 5329 58223 5415 58279
rect 5471 58223 5557 58279
rect 5613 58223 5699 58279
rect 5755 58223 5841 58279
rect 5897 58223 5983 58279
rect 6039 58223 6125 58279
rect 6181 58223 6267 58279
rect 6323 58223 6409 58279
rect 6465 58223 6551 58279
rect 6607 58223 6693 58279
rect 6749 58223 6835 58279
rect 6891 58223 6977 58279
rect 7033 58223 7119 58279
rect 7175 58223 7261 58279
rect 7317 58223 7403 58279
rect 7459 58223 7545 58279
rect 7601 58223 7687 58279
rect 7743 58223 7829 58279
rect 7885 58223 7971 58279
rect 8027 58223 8113 58279
rect 8169 58223 8255 58279
rect 8311 58223 8397 58279
rect 8453 58223 8539 58279
rect 8595 58223 8681 58279
rect 8737 58223 8823 58279
rect 8879 58223 8965 58279
rect 9021 58223 9107 58279
rect 9163 58223 9249 58279
rect 9305 58223 9391 58279
rect 9447 58223 9533 58279
rect 9589 58223 9675 58279
rect 9731 58223 9817 58279
rect 9873 58223 9959 58279
rect 10015 58223 10101 58279
rect 10157 58223 10243 58279
rect 10299 58223 10385 58279
rect 10441 58223 10527 58279
rect 10583 58223 10669 58279
rect 10725 58223 10811 58279
rect 10867 58223 10953 58279
rect 11009 58223 11095 58279
rect 11151 58223 11237 58279
rect 11293 58223 11379 58279
rect 11435 58223 11521 58279
rect 11577 58223 11663 58279
rect 11719 58223 11805 58279
rect 11861 58223 11947 58279
rect 12003 58223 12089 58279
rect 12145 58223 12231 58279
rect 12287 58223 12373 58279
rect 12429 58223 12515 58279
rect 12571 58223 12657 58279
rect 12713 58223 12799 58279
rect 12855 58223 12941 58279
rect 12997 58223 13083 58279
rect 13139 58223 13225 58279
rect 13281 58223 13367 58279
rect 13423 58223 13509 58279
rect 13565 58223 13651 58279
rect 13707 58223 13793 58279
rect 13849 58223 13935 58279
rect 13991 58223 14077 58279
rect 14133 58223 14219 58279
rect 14275 58223 14361 58279
rect 14417 58223 14503 58279
rect 14559 58223 14645 58279
rect 14701 58223 14787 58279
rect 14843 58223 15000 58279
rect 0 58137 15000 58223
rect 0 58081 161 58137
rect 217 58081 303 58137
rect 359 58081 445 58137
rect 501 58081 587 58137
rect 643 58081 729 58137
rect 785 58081 871 58137
rect 927 58081 1013 58137
rect 1069 58081 1155 58137
rect 1211 58081 1297 58137
rect 1353 58081 1439 58137
rect 1495 58081 1581 58137
rect 1637 58081 1723 58137
rect 1779 58081 1865 58137
rect 1921 58081 2007 58137
rect 2063 58081 2149 58137
rect 2205 58081 2291 58137
rect 2347 58081 2433 58137
rect 2489 58081 2575 58137
rect 2631 58081 2717 58137
rect 2773 58081 2859 58137
rect 2915 58081 3001 58137
rect 3057 58081 3143 58137
rect 3199 58081 3285 58137
rect 3341 58081 3427 58137
rect 3483 58081 3569 58137
rect 3625 58081 3711 58137
rect 3767 58081 3853 58137
rect 3909 58081 3995 58137
rect 4051 58081 4137 58137
rect 4193 58081 4279 58137
rect 4335 58081 4421 58137
rect 4477 58081 4563 58137
rect 4619 58081 4705 58137
rect 4761 58081 4847 58137
rect 4903 58081 4989 58137
rect 5045 58081 5131 58137
rect 5187 58081 5273 58137
rect 5329 58081 5415 58137
rect 5471 58081 5557 58137
rect 5613 58081 5699 58137
rect 5755 58081 5841 58137
rect 5897 58081 5983 58137
rect 6039 58081 6125 58137
rect 6181 58081 6267 58137
rect 6323 58081 6409 58137
rect 6465 58081 6551 58137
rect 6607 58081 6693 58137
rect 6749 58081 6835 58137
rect 6891 58081 6977 58137
rect 7033 58081 7119 58137
rect 7175 58081 7261 58137
rect 7317 58081 7403 58137
rect 7459 58081 7545 58137
rect 7601 58081 7687 58137
rect 7743 58081 7829 58137
rect 7885 58081 7971 58137
rect 8027 58081 8113 58137
rect 8169 58081 8255 58137
rect 8311 58081 8397 58137
rect 8453 58081 8539 58137
rect 8595 58081 8681 58137
rect 8737 58081 8823 58137
rect 8879 58081 8965 58137
rect 9021 58081 9107 58137
rect 9163 58081 9249 58137
rect 9305 58081 9391 58137
rect 9447 58081 9533 58137
rect 9589 58081 9675 58137
rect 9731 58081 9817 58137
rect 9873 58081 9959 58137
rect 10015 58081 10101 58137
rect 10157 58081 10243 58137
rect 10299 58081 10385 58137
rect 10441 58081 10527 58137
rect 10583 58081 10669 58137
rect 10725 58081 10811 58137
rect 10867 58081 10953 58137
rect 11009 58081 11095 58137
rect 11151 58081 11237 58137
rect 11293 58081 11379 58137
rect 11435 58081 11521 58137
rect 11577 58081 11663 58137
rect 11719 58081 11805 58137
rect 11861 58081 11947 58137
rect 12003 58081 12089 58137
rect 12145 58081 12231 58137
rect 12287 58081 12373 58137
rect 12429 58081 12515 58137
rect 12571 58081 12657 58137
rect 12713 58081 12799 58137
rect 12855 58081 12941 58137
rect 12997 58081 13083 58137
rect 13139 58081 13225 58137
rect 13281 58081 13367 58137
rect 13423 58081 13509 58137
rect 13565 58081 13651 58137
rect 13707 58081 13793 58137
rect 13849 58081 13935 58137
rect 13991 58081 14077 58137
rect 14133 58081 14219 58137
rect 14275 58081 14361 58137
rect 14417 58081 14503 58137
rect 14559 58081 14645 58137
rect 14701 58081 14787 58137
rect 14843 58081 15000 58137
rect 0 57995 15000 58081
rect 0 57939 161 57995
rect 217 57939 303 57995
rect 359 57939 445 57995
rect 501 57939 587 57995
rect 643 57939 729 57995
rect 785 57939 871 57995
rect 927 57939 1013 57995
rect 1069 57939 1155 57995
rect 1211 57939 1297 57995
rect 1353 57939 1439 57995
rect 1495 57939 1581 57995
rect 1637 57939 1723 57995
rect 1779 57939 1865 57995
rect 1921 57939 2007 57995
rect 2063 57939 2149 57995
rect 2205 57939 2291 57995
rect 2347 57939 2433 57995
rect 2489 57939 2575 57995
rect 2631 57939 2717 57995
rect 2773 57939 2859 57995
rect 2915 57939 3001 57995
rect 3057 57939 3143 57995
rect 3199 57939 3285 57995
rect 3341 57939 3427 57995
rect 3483 57939 3569 57995
rect 3625 57939 3711 57995
rect 3767 57939 3853 57995
rect 3909 57939 3995 57995
rect 4051 57939 4137 57995
rect 4193 57939 4279 57995
rect 4335 57939 4421 57995
rect 4477 57939 4563 57995
rect 4619 57939 4705 57995
rect 4761 57939 4847 57995
rect 4903 57939 4989 57995
rect 5045 57939 5131 57995
rect 5187 57939 5273 57995
rect 5329 57939 5415 57995
rect 5471 57939 5557 57995
rect 5613 57939 5699 57995
rect 5755 57939 5841 57995
rect 5897 57939 5983 57995
rect 6039 57939 6125 57995
rect 6181 57939 6267 57995
rect 6323 57939 6409 57995
rect 6465 57939 6551 57995
rect 6607 57939 6693 57995
rect 6749 57939 6835 57995
rect 6891 57939 6977 57995
rect 7033 57939 7119 57995
rect 7175 57939 7261 57995
rect 7317 57939 7403 57995
rect 7459 57939 7545 57995
rect 7601 57939 7687 57995
rect 7743 57939 7829 57995
rect 7885 57939 7971 57995
rect 8027 57939 8113 57995
rect 8169 57939 8255 57995
rect 8311 57939 8397 57995
rect 8453 57939 8539 57995
rect 8595 57939 8681 57995
rect 8737 57939 8823 57995
rect 8879 57939 8965 57995
rect 9021 57939 9107 57995
rect 9163 57939 9249 57995
rect 9305 57939 9391 57995
rect 9447 57939 9533 57995
rect 9589 57939 9675 57995
rect 9731 57939 9817 57995
rect 9873 57939 9959 57995
rect 10015 57939 10101 57995
rect 10157 57939 10243 57995
rect 10299 57939 10385 57995
rect 10441 57939 10527 57995
rect 10583 57939 10669 57995
rect 10725 57939 10811 57995
rect 10867 57939 10953 57995
rect 11009 57939 11095 57995
rect 11151 57939 11237 57995
rect 11293 57939 11379 57995
rect 11435 57939 11521 57995
rect 11577 57939 11663 57995
rect 11719 57939 11805 57995
rect 11861 57939 11947 57995
rect 12003 57939 12089 57995
rect 12145 57939 12231 57995
rect 12287 57939 12373 57995
rect 12429 57939 12515 57995
rect 12571 57939 12657 57995
rect 12713 57939 12799 57995
rect 12855 57939 12941 57995
rect 12997 57939 13083 57995
rect 13139 57939 13225 57995
rect 13281 57939 13367 57995
rect 13423 57939 13509 57995
rect 13565 57939 13651 57995
rect 13707 57939 13793 57995
rect 13849 57939 13935 57995
rect 13991 57939 14077 57995
rect 14133 57939 14219 57995
rect 14275 57939 14361 57995
rect 14417 57939 14503 57995
rect 14559 57939 14645 57995
rect 14701 57939 14787 57995
rect 14843 57939 15000 57995
rect 0 57853 15000 57939
rect 0 57797 161 57853
rect 217 57797 303 57853
rect 359 57797 445 57853
rect 501 57797 587 57853
rect 643 57797 729 57853
rect 785 57797 871 57853
rect 927 57797 1013 57853
rect 1069 57797 1155 57853
rect 1211 57797 1297 57853
rect 1353 57797 1439 57853
rect 1495 57797 1581 57853
rect 1637 57797 1723 57853
rect 1779 57797 1865 57853
rect 1921 57797 2007 57853
rect 2063 57797 2149 57853
rect 2205 57797 2291 57853
rect 2347 57797 2433 57853
rect 2489 57797 2575 57853
rect 2631 57797 2717 57853
rect 2773 57797 2859 57853
rect 2915 57797 3001 57853
rect 3057 57797 3143 57853
rect 3199 57797 3285 57853
rect 3341 57797 3427 57853
rect 3483 57797 3569 57853
rect 3625 57797 3711 57853
rect 3767 57797 3853 57853
rect 3909 57797 3995 57853
rect 4051 57797 4137 57853
rect 4193 57797 4279 57853
rect 4335 57797 4421 57853
rect 4477 57797 4563 57853
rect 4619 57797 4705 57853
rect 4761 57797 4847 57853
rect 4903 57797 4989 57853
rect 5045 57797 5131 57853
rect 5187 57797 5273 57853
rect 5329 57797 5415 57853
rect 5471 57797 5557 57853
rect 5613 57797 5699 57853
rect 5755 57797 5841 57853
rect 5897 57797 5983 57853
rect 6039 57797 6125 57853
rect 6181 57797 6267 57853
rect 6323 57797 6409 57853
rect 6465 57797 6551 57853
rect 6607 57797 6693 57853
rect 6749 57797 6835 57853
rect 6891 57797 6977 57853
rect 7033 57797 7119 57853
rect 7175 57797 7261 57853
rect 7317 57797 7403 57853
rect 7459 57797 7545 57853
rect 7601 57797 7687 57853
rect 7743 57797 7829 57853
rect 7885 57797 7971 57853
rect 8027 57797 8113 57853
rect 8169 57797 8255 57853
rect 8311 57797 8397 57853
rect 8453 57797 8539 57853
rect 8595 57797 8681 57853
rect 8737 57797 8823 57853
rect 8879 57797 8965 57853
rect 9021 57797 9107 57853
rect 9163 57797 9249 57853
rect 9305 57797 9391 57853
rect 9447 57797 9533 57853
rect 9589 57797 9675 57853
rect 9731 57797 9817 57853
rect 9873 57797 9959 57853
rect 10015 57797 10101 57853
rect 10157 57797 10243 57853
rect 10299 57797 10385 57853
rect 10441 57797 10527 57853
rect 10583 57797 10669 57853
rect 10725 57797 10811 57853
rect 10867 57797 10953 57853
rect 11009 57797 11095 57853
rect 11151 57797 11237 57853
rect 11293 57797 11379 57853
rect 11435 57797 11521 57853
rect 11577 57797 11663 57853
rect 11719 57797 11805 57853
rect 11861 57797 11947 57853
rect 12003 57797 12089 57853
rect 12145 57797 12231 57853
rect 12287 57797 12373 57853
rect 12429 57797 12515 57853
rect 12571 57797 12657 57853
rect 12713 57797 12799 57853
rect 12855 57797 12941 57853
rect 12997 57797 13083 57853
rect 13139 57797 13225 57853
rect 13281 57797 13367 57853
rect 13423 57797 13509 57853
rect 13565 57797 13651 57853
rect 13707 57797 13793 57853
rect 13849 57797 13935 57853
rect 13991 57797 14077 57853
rect 14133 57797 14219 57853
rect 14275 57797 14361 57853
rect 14417 57797 14503 57853
rect 14559 57797 14645 57853
rect 14701 57797 14787 57853
rect 14843 57797 15000 57853
rect 0 57711 15000 57797
rect 0 57655 161 57711
rect 217 57655 303 57711
rect 359 57655 445 57711
rect 501 57655 587 57711
rect 643 57655 729 57711
rect 785 57655 871 57711
rect 927 57655 1013 57711
rect 1069 57655 1155 57711
rect 1211 57655 1297 57711
rect 1353 57655 1439 57711
rect 1495 57655 1581 57711
rect 1637 57655 1723 57711
rect 1779 57655 1865 57711
rect 1921 57655 2007 57711
rect 2063 57655 2149 57711
rect 2205 57655 2291 57711
rect 2347 57655 2433 57711
rect 2489 57655 2575 57711
rect 2631 57655 2717 57711
rect 2773 57655 2859 57711
rect 2915 57655 3001 57711
rect 3057 57655 3143 57711
rect 3199 57655 3285 57711
rect 3341 57655 3427 57711
rect 3483 57655 3569 57711
rect 3625 57655 3711 57711
rect 3767 57655 3853 57711
rect 3909 57655 3995 57711
rect 4051 57655 4137 57711
rect 4193 57655 4279 57711
rect 4335 57655 4421 57711
rect 4477 57655 4563 57711
rect 4619 57655 4705 57711
rect 4761 57655 4847 57711
rect 4903 57655 4989 57711
rect 5045 57655 5131 57711
rect 5187 57655 5273 57711
rect 5329 57655 5415 57711
rect 5471 57655 5557 57711
rect 5613 57655 5699 57711
rect 5755 57655 5841 57711
rect 5897 57655 5983 57711
rect 6039 57655 6125 57711
rect 6181 57655 6267 57711
rect 6323 57655 6409 57711
rect 6465 57655 6551 57711
rect 6607 57655 6693 57711
rect 6749 57655 6835 57711
rect 6891 57655 6977 57711
rect 7033 57655 7119 57711
rect 7175 57655 7261 57711
rect 7317 57655 7403 57711
rect 7459 57655 7545 57711
rect 7601 57655 7687 57711
rect 7743 57655 7829 57711
rect 7885 57655 7971 57711
rect 8027 57655 8113 57711
rect 8169 57655 8255 57711
rect 8311 57655 8397 57711
rect 8453 57655 8539 57711
rect 8595 57655 8681 57711
rect 8737 57655 8823 57711
rect 8879 57655 8965 57711
rect 9021 57655 9107 57711
rect 9163 57655 9249 57711
rect 9305 57655 9391 57711
rect 9447 57655 9533 57711
rect 9589 57655 9675 57711
rect 9731 57655 9817 57711
rect 9873 57655 9959 57711
rect 10015 57655 10101 57711
rect 10157 57655 10243 57711
rect 10299 57655 10385 57711
rect 10441 57655 10527 57711
rect 10583 57655 10669 57711
rect 10725 57655 10811 57711
rect 10867 57655 10953 57711
rect 11009 57655 11095 57711
rect 11151 57655 11237 57711
rect 11293 57655 11379 57711
rect 11435 57655 11521 57711
rect 11577 57655 11663 57711
rect 11719 57655 11805 57711
rect 11861 57655 11947 57711
rect 12003 57655 12089 57711
rect 12145 57655 12231 57711
rect 12287 57655 12373 57711
rect 12429 57655 12515 57711
rect 12571 57655 12657 57711
rect 12713 57655 12799 57711
rect 12855 57655 12941 57711
rect 12997 57655 13083 57711
rect 13139 57655 13225 57711
rect 13281 57655 13367 57711
rect 13423 57655 13509 57711
rect 13565 57655 13651 57711
rect 13707 57655 13793 57711
rect 13849 57655 13935 57711
rect 13991 57655 14077 57711
rect 14133 57655 14219 57711
rect 14275 57655 14361 57711
rect 14417 57655 14503 57711
rect 14559 57655 14645 57711
rect 14701 57655 14787 57711
rect 14843 57655 15000 57711
rect 0 57569 15000 57655
rect 0 57513 161 57569
rect 217 57513 303 57569
rect 359 57513 445 57569
rect 501 57513 587 57569
rect 643 57513 729 57569
rect 785 57513 871 57569
rect 927 57513 1013 57569
rect 1069 57513 1155 57569
rect 1211 57513 1297 57569
rect 1353 57513 1439 57569
rect 1495 57513 1581 57569
rect 1637 57513 1723 57569
rect 1779 57513 1865 57569
rect 1921 57513 2007 57569
rect 2063 57513 2149 57569
rect 2205 57513 2291 57569
rect 2347 57513 2433 57569
rect 2489 57513 2575 57569
rect 2631 57513 2717 57569
rect 2773 57513 2859 57569
rect 2915 57513 3001 57569
rect 3057 57513 3143 57569
rect 3199 57513 3285 57569
rect 3341 57513 3427 57569
rect 3483 57513 3569 57569
rect 3625 57513 3711 57569
rect 3767 57513 3853 57569
rect 3909 57513 3995 57569
rect 4051 57513 4137 57569
rect 4193 57513 4279 57569
rect 4335 57513 4421 57569
rect 4477 57513 4563 57569
rect 4619 57513 4705 57569
rect 4761 57513 4847 57569
rect 4903 57513 4989 57569
rect 5045 57513 5131 57569
rect 5187 57513 5273 57569
rect 5329 57513 5415 57569
rect 5471 57513 5557 57569
rect 5613 57513 5699 57569
rect 5755 57513 5841 57569
rect 5897 57513 5983 57569
rect 6039 57513 6125 57569
rect 6181 57513 6267 57569
rect 6323 57513 6409 57569
rect 6465 57513 6551 57569
rect 6607 57513 6693 57569
rect 6749 57513 6835 57569
rect 6891 57513 6977 57569
rect 7033 57513 7119 57569
rect 7175 57513 7261 57569
rect 7317 57513 7403 57569
rect 7459 57513 7545 57569
rect 7601 57513 7687 57569
rect 7743 57513 7829 57569
rect 7885 57513 7971 57569
rect 8027 57513 8113 57569
rect 8169 57513 8255 57569
rect 8311 57513 8397 57569
rect 8453 57513 8539 57569
rect 8595 57513 8681 57569
rect 8737 57513 8823 57569
rect 8879 57513 8965 57569
rect 9021 57513 9107 57569
rect 9163 57513 9249 57569
rect 9305 57513 9391 57569
rect 9447 57513 9533 57569
rect 9589 57513 9675 57569
rect 9731 57513 9817 57569
rect 9873 57513 9959 57569
rect 10015 57513 10101 57569
rect 10157 57513 10243 57569
rect 10299 57513 10385 57569
rect 10441 57513 10527 57569
rect 10583 57513 10669 57569
rect 10725 57513 10811 57569
rect 10867 57513 10953 57569
rect 11009 57513 11095 57569
rect 11151 57513 11237 57569
rect 11293 57513 11379 57569
rect 11435 57513 11521 57569
rect 11577 57513 11663 57569
rect 11719 57513 11805 57569
rect 11861 57513 11947 57569
rect 12003 57513 12089 57569
rect 12145 57513 12231 57569
rect 12287 57513 12373 57569
rect 12429 57513 12515 57569
rect 12571 57513 12657 57569
rect 12713 57513 12799 57569
rect 12855 57513 12941 57569
rect 12997 57513 13083 57569
rect 13139 57513 13225 57569
rect 13281 57513 13367 57569
rect 13423 57513 13509 57569
rect 13565 57513 13651 57569
rect 13707 57513 13793 57569
rect 13849 57513 13935 57569
rect 13991 57513 14077 57569
rect 14133 57513 14219 57569
rect 14275 57513 14361 57569
rect 14417 57513 14503 57569
rect 14559 57513 14645 57569
rect 14701 57513 14787 57569
rect 14843 57513 15000 57569
rect 0 57427 15000 57513
rect 0 57371 161 57427
rect 217 57371 303 57427
rect 359 57371 445 57427
rect 501 57371 587 57427
rect 643 57371 729 57427
rect 785 57371 871 57427
rect 927 57371 1013 57427
rect 1069 57371 1155 57427
rect 1211 57371 1297 57427
rect 1353 57371 1439 57427
rect 1495 57371 1581 57427
rect 1637 57371 1723 57427
rect 1779 57371 1865 57427
rect 1921 57371 2007 57427
rect 2063 57371 2149 57427
rect 2205 57371 2291 57427
rect 2347 57371 2433 57427
rect 2489 57371 2575 57427
rect 2631 57371 2717 57427
rect 2773 57371 2859 57427
rect 2915 57371 3001 57427
rect 3057 57371 3143 57427
rect 3199 57371 3285 57427
rect 3341 57371 3427 57427
rect 3483 57371 3569 57427
rect 3625 57371 3711 57427
rect 3767 57371 3853 57427
rect 3909 57371 3995 57427
rect 4051 57371 4137 57427
rect 4193 57371 4279 57427
rect 4335 57371 4421 57427
rect 4477 57371 4563 57427
rect 4619 57371 4705 57427
rect 4761 57371 4847 57427
rect 4903 57371 4989 57427
rect 5045 57371 5131 57427
rect 5187 57371 5273 57427
rect 5329 57371 5415 57427
rect 5471 57371 5557 57427
rect 5613 57371 5699 57427
rect 5755 57371 5841 57427
rect 5897 57371 5983 57427
rect 6039 57371 6125 57427
rect 6181 57371 6267 57427
rect 6323 57371 6409 57427
rect 6465 57371 6551 57427
rect 6607 57371 6693 57427
rect 6749 57371 6835 57427
rect 6891 57371 6977 57427
rect 7033 57371 7119 57427
rect 7175 57371 7261 57427
rect 7317 57371 7403 57427
rect 7459 57371 7545 57427
rect 7601 57371 7687 57427
rect 7743 57371 7829 57427
rect 7885 57371 7971 57427
rect 8027 57371 8113 57427
rect 8169 57371 8255 57427
rect 8311 57371 8397 57427
rect 8453 57371 8539 57427
rect 8595 57371 8681 57427
rect 8737 57371 8823 57427
rect 8879 57371 8965 57427
rect 9021 57371 9107 57427
rect 9163 57371 9249 57427
rect 9305 57371 9391 57427
rect 9447 57371 9533 57427
rect 9589 57371 9675 57427
rect 9731 57371 9817 57427
rect 9873 57371 9959 57427
rect 10015 57371 10101 57427
rect 10157 57371 10243 57427
rect 10299 57371 10385 57427
rect 10441 57371 10527 57427
rect 10583 57371 10669 57427
rect 10725 57371 10811 57427
rect 10867 57371 10953 57427
rect 11009 57371 11095 57427
rect 11151 57371 11237 57427
rect 11293 57371 11379 57427
rect 11435 57371 11521 57427
rect 11577 57371 11663 57427
rect 11719 57371 11805 57427
rect 11861 57371 11947 57427
rect 12003 57371 12089 57427
rect 12145 57371 12231 57427
rect 12287 57371 12373 57427
rect 12429 57371 12515 57427
rect 12571 57371 12657 57427
rect 12713 57371 12799 57427
rect 12855 57371 12941 57427
rect 12997 57371 13083 57427
rect 13139 57371 13225 57427
rect 13281 57371 13367 57427
rect 13423 57371 13509 57427
rect 13565 57371 13651 57427
rect 13707 57371 13793 57427
rect 13849 57371 13935 57427
rect 13991 57371 14077 57427
rect 14133 57371 14219 57427
rect 14275 57371 14361 57427
rect 14417 57371 14503 57427
rect 14559 57371 14645 57427
rect 14701 57371 14787 57427
rect 14843 57371 15000 57427
rect 0 57285 15000 57371
rect 0 57229 161 57285
rect 217 57229 303 57285
rect 359 57229 445 57285
rect 501 57229 587 57285
rect 643 57229 729 57285
rect 785 57229 871 57285
rect 927 57229 1013 57285
rect 1069 57229 1155 57285
rect 1211 57229 1297 57285
rect 1353 57229 1439 57285
rect 1495 57229 1581 57285
rect 1637 57229 1723 57285
rect 1779 57229 1865 57285
rect 1921 57229 2007 57285
rect 2063 57229 2149 57285
rect 2205 57229 2291 57285
rect 2347 57229 2433 57285
rect 2489 57229 2575 57285
rect 2631 57229 2717 57285
rect 2773 57229 2859 57285
rect 2915 57229 3001 57285
rect 3057 57229 3143 57285
rect 3199 57229 3285 57285
rect 3341 57229 3427 57285
rect 3483 57229 3569 57285
rect 3625 57229 3711 57285
rect 3767 57229 3853 57285
rect 3909 57229 3995 57285
rect 4051 57229 4137 57285
rect 4193 57229 4279 57285
rect 4335 57229 4421 57285
rect 4477 57229 4563 57285
rect 4619 57229 4705 57285
rect 4761 57229 4847 57285
rect 4903 57229 4989 57285
rect 5045 57229 5131 57285
rect 5187 57229 5273 57285
rect 5329 57229 5415 57285
rect 5471 57229 5557 57285
rect 5613 57229 5699 57285
rect 5755 57229 5841 57285
rect 5897 57229 5983 57285
rect 6039 57229 6125 57285
rect 6181 57229 6267 57285
rect 6323 57229 6409 57285
rect 6465 57229 6551 57285
rect 6607 57229 6693 57285
rect 6749 57229 6835 57285
rect 6891 57229 6977 57285
rect 7033 57229 7119 57285
rect 7175 57229 7261 57285
rect 7317 57229 7403 57285
rect 7459 57229 7545 57285
rect 7601 57229 7687 57285
rect 7743 57229 7829 57285
rect 7885 57229 7971 57285
rect 8027 57229 8113 57285
rect 8169 57229 8255 57285
rect 8311 57229 8397 57285
rect 8453 57229 8539 57285
rect 8595 57229 8681 57285
rect 8737 57229 8823 57285
rect 8879 57229 8965 57285
rect 9021 57229 9107 57285
rect 9163 57229 9249 57285
rect 9305 57229 9391 57285
rect 9447 57229 9533 57285
rect 9589 57229 9675 57285
rect 9731 57229 9817 57285
rect 9873 57229 9959 57285
rect 10015 57229 10101 57285
rect 10157 57229 10243 57285
rect 10299 57229 10385 57285
rect 10441 57229 10527 57285
rect 10583 57229 10669 57285
rect 10725 57229 10811 57285
rect 10867 57229 10953 57285
rect 11009 57229 11095 57285
rect 11151 57229 11237 57285
rect 11293 57229 11379 57285
rect 11435 57229 11521 57285
rect 11577 57229 11663 57285
rect 11719 57229 11805 57285
rect 11861 57229 11947 57285
rect 12003 57229 12089 57285
rect 12145 57229 12231 57285
rect 12287 57229 12373 57285
rect 12429 57229 12515 57285
rect 12571 57229 12657 57285
rect 12713 57229 12799 57285
rect 12855 57229 12941 57285
rect 12997 57229 13083 57285
rect 13139 57229 13225 57285
rect 13281 57229 13367 57285
rect 13423 57229 13509 57285
rect 13565 57229 13651 57285
rect 13707 57229 13793 57285
rect 13849 57229 13935 57285
rect 13991 57229 14077 57285
rect 14133 57229 14219 57285
rect 14275 57229 14361 57285
rect 14417 57229 14503 57285
rect 14559 57229 14645 57285
rect 14701 57229 14787 57285
rect 14843 57229 15000 57285
rect 0 57200 15000 57229
rect 0 56971 15000 57000
rect 0 56915 161 56971
rect 217 56915 303 56971
rect 359 56915 445 56971
rect 501 56915 587 56971
rect 643 56915 729 56971
rect 785 56915 871 56971
rect 927 56915 1013 56971
rect 1069 56915 1155 56971
rect 1211 56915 1297 56971
rect 1353 56915 1439 56971
rect 1495 56915 1581 56971
rect 1637 56915 1723 56971
rect 1779 56915 1865 56971
rect 1921 56915 2007 56971
rect 2063 56915 2149 56971
rect 2205 56915 2291 56971
rect 2347 56915 2433 56971
rect 2489 56915 2575 56971
rect 2631 56915 2717 56971
rect 2773 56915 2859 56971
rect 2915 56915 3001 56971
rect 3057 56915 3143 56971
rect 3199 56915 3285 56971
rect 3341 56915 3427 56971
rect 3483 56915 3569 56971
rect 3625 56915 3711 56971
rect 3767 56915 3853 56971
rect 3909 56915 3995 56971
rect 4051 56915 4137 56971
rect 4193 56915 4279 56971
rect 4335 56915 4421 56971
rect 4477 56915 4563 56971
rect 4619 56915 4705 56971
rect 4761 56915 4847 56971
rect 4903 56915 4989 56971
rect 5045 56915 5131 56971
rect 5187 56915 5273 56971
rect 5329 56915 5415 56971
rect 5471 56915 5557 56971
rect 5613 56915 5699 56971
rect 5755 56915 5841 56971
rect 5897 56915 5983 56971
rect 6039 56915 6125 56971
rect 6181 56915 6267 56971
rect 6323 56915 6409 56971
rect 6465 56915 6551 56971
rect 6607 56915 6693 56971
rect 6749 56915 6835 56971
rect 6891 56915 6977 56971
rect 7033 56915 7119 56971
rect 7175 56915 7261 56971
rect 7317 56915 7403 56971
rect 7459 56915 7545 56971
rect 7601 56915 7687 56971
rect 7743 56915 7829 56971
rect 7885 56915 7971 56971
rect 8027 56915 8113 56971
rect 8169 56915 8255 56971
rect 8311 56915 8397 56971
rect 8453 56915 8539 56971
rect 8595 56915 8681 56971
rect 8737 56915 8823 56971
rect 8879 56915 8965 56971
rect 9021 56915 9107 56971
rect 9163 56915 9249 56971
rect 9305 56915 9391 56971
rect 9447 56915 9533 56971
rect 9589 56915 9675 56971
rect 9731 56915 9817 56971
rect 9873 56915 9959 56971
rect 10015 56915 10101 56971
rect 10157 56915 10243 56971
rect 10299 56915 10385 56971
rect 10441 56915 10527 56971
rect 10583 56915 10669 56971
rect 10725 56915 10811 56971
rect 10867 56915 10953 56971
rect 11009 56915 11095 56971
rect 11151 56915 11237 56971
rect 11293 56915 11379 56971
rect 11435 56915 11521 56971
rect 11577 56915 11663 56971
rect 11719 56915 11805 56971
rect 11861 56915 11947 56971
rect 12003 56915 12089 56971
rect 12145 56915 12231 56971
rect 12287 56915 12373 56971
rect 12429 56915 12515 56971
rect 12571 56915 12657 56971
rect 12713 56915 12799 56971
rect 12855 56915 12941 56971
rect 12997 56915 13083 56971
rect 13139 56915 13225 56971
rect 13281 56915 13367 56971
rect 13423 56915 13509 56971
rect 13565 56915 13651 56971
rect 13707 56915 13793 56971
rect 13849 56915 13935 56971
rect 13991 56915 14077 56971
rect 14133 56915 14219 56971
rect 14275 56915 14361 56971
rect 14417 56915 14503 56971
rect 14559 56915 14645 56971
rect 14701 56915 14787 56971
rect 14843 56915 15000 56971
rect 0 56829 15000 56915
rect 0 56773 161 56829
rect 217 56773 303 56829
rect 359 56773 445 56829
rect 501 56773 587 56829
rect 643 56773 729 56829
rect 785 56773 871 56829
rect 927 56773 1013 56829
rect 1069 56773 1155 56829
rect 1211 56773 1297 56829
rect 1353 56773 1439 56829
rect 1495 56773 1581 56829
rect 1637 56773 1723 56829
rect 1779 56773 1865 56829
rect 1921 56773 2007 56829
rect 2063 56773 2149 56829
rect 2205 56773 2291 56829
rect 2347 56773 2433 56829
rect 2489 56773 2575 56829
rect 2631 56773 2717 56829
rect 2773 56773 2859 56829
rect 2915 56773 3001 56829
rect 3057 56773 3143 56829
rect 3199 56773 3285 56829
rect 3341 56773 3427 56829
rect 3483 56773 3569 56829
rect 3625 56773 3711 56829
rect 3767 56773 3853 56829
rect 3909 56773 3995 56829
rect 4051 56773 4137 56829
rect 4193 56773 4279 56829
rect 4335 56773 4421 56829
rect 4477 56773 4563 56829
rect 4619 56773 4705 56829
rect 4761 56773 4847 56829
rect 4903 56773 4989 56829
rect 5045 56773 5131 56829
rect 5187 56773 5273 56829
rect 5329 56773 5415 56829
rect 5471 56773 5557 56829
rect 5613 56773 5699 56829
rect 5755 56773 5841 56829
rect 5897 56773 5983 56829
rect 6039 56773 6125 56829
rect 6181 56773 6267 56829
rect 6323 56773 6409 56829
rect 6465 56773 6551 56829
rect 6607 56773 6693 56829
rect 6749 56773 6835 56829
rect 6891 56773 6977 56829
rect 7033 56773 7119 56829
rect 7175 56773 7261 56829
rect 7317 56773 7403 56829
rect 7459 56773 7545 56829
rect 7601 56773 7687 56829
rect 7743 56773 7829 56829
rect 7885 56773 7971 56829
rect 8027 56773 8113 56829
rect 8169 56773 8255 56829
rect 8311 56773 8397 56829
rect 8453 56773 8539 56829
rect 8595 56773 8681 56829
rect 8737 56773 8823 56829
rect 8879 56773 8965 56829
rect 9021 56773 9107 56829
rect 9163 56773 9249 56829
rect 9305 56773 9391 56829
rect 9447 56773 9533 56829
rect 9589 56773 9675 56829
rect 9731 56773 9817 56829
rect 9873 56773 9959 56829
rect 10015 56773 10101 56829
rect 10157 56773 10243 56829
rect 10299 56773 10385 56829
rect 10441 56773 10527 56829
rect 10583 56773 10669 56829
rect 10725 56773 10811 56829
rect 10867 56773 10953 56829
rect 11009 56773 11095 56829
rect 11151 56773 11237 56829
rect 11293 56773 11379 56829
rect 11435 56773 11521 56829
rect 11577 56773 11663 56829
rect 11719 56773 11805 56829
rect 11861 56773 11947 56829
rect 12003 56773 12089 56829
rect 12145 56773 12231 56829
rect 12287 56773 12373 56829
rect 12429 56773 12515 56829
rect 12571 56773 12657 56829
rect 12713 56773 12799 56829
rect 12855 56773 12941 56829
rect 12997 56773 13083 56829
rect 13139 56773 13225 56829
rect 13281 56773 13367 56829
rect 13423 56773 13509 56829
rect 13565 56773 13651 56829
rect 13707 56773 13793 56829
rect 13849 56773 13935 56829
rect 13991 56773 14077 56829
rect 14133 56773 14219 56829
rect 14275 56773 14361 56829
rect 14417 56773 14503 56829
rect 14559 56773 14645 56829
rect 14701 56773 14787 56829
rect 14843 56773 15000 56829
rect 0 56687 15000 56773
rect 0 56631 161 56687
rect 217 56631 303 56687
rect 359 56631 445 56687
rect 501 56631 587 56687
rect 643 56631 729 56687
rect 785 56631 871 56687
rect 927 56631 1013 56687
rect 1069 56631 1155 56687
rect 1211 56631 1297 56687
rect 1353 56631 1439 56687
rect 1495 56631 1581 56687
rect 1637 56631 1723 56687
rect 1779 56631 1865 56687
rect 1921 56631 2007 56687
rect 2063 56631 2149 56687
rect 2205 56631 2291 56687
rect 2347 56631 2433 56687
rect 2489 56631 2575 56687
rect 2631 56631 2717 56687
rect 2773 56631 2859 56687
rect 2915 56631 3001 56687
rect 3057 56631 3143 56687
rect 3199 56631 3285 56687
rect 3341 56631 3427 56687
rect 3483 56631 3569 56687
rect 3625 56631 3711 56687
rect 3767 56631 3853 56687
rect 3909 56631 3995 56687
rect 4051 56631 4137 56687
rect 4193 56631 4279 56687
rect 4335 56631 4421 56687
rect 4477 56631 4563 56687
rect 4619 56631 4705 56687
rect 4761 56631 4847 56687
rect 4903 56631 4989 56687
rect 5045 56631 5131 56687
rect 5187 56631 5273 56687
rect 5329 56631 5415 56687
rect 5471 56631 5557 56687
rect 5613 56631 5699 56687
rect 5755 56631 5841 56687
rect 5897 56631 5983 56687
rect 6039 56631 6125 56687
rect 6181 56631 6267 56687
rect 6323 56631 6409 56687
rect 6465 56631 6551 56687
rect 6607 56631 6693 56687
rect 6749 56631 6835 56687
rect 6891 56631 6977 56687
rect 7033 56631 7119 56687
rect 7175 56631 7261 56687
rect 7317 56631 7403 56687
rect 7459 56631 7545 56687
rect 7601 56631 7687 56687
rect 7743 56631 7829 56687
rect 7885 56631 7971 56687
rect 8027 56631 8113 56687
rect 8169 56631 8255 56687
rect 8311 56631 8397 56687
rect 8453 56631 8539 56687
rect 8595 56631 8681 56687
rect 8737 56631 8823 56687
rect 8879 56631 8965 56687
rect 9021 56631 9107 56687
rect 9163 56631 9249 56687
rect 9305 56631 9391 56687
rect 9447 56631 9533 56687
rect 9589 56631 9675 56687
rect 9731 56631 9817 56687
rect 9873 56631 9959 56687
rect 10015 56631 10101 56687
rect 10157 56631 10243 56687
rect 10299 56631 10385 56687
rect 10441 56631 10527 56687
rect 10583 56631 10669 56687
rect 10725 56631 10811 56687
rect 10867 56631 10953 56687
rect 11009 56631 11095 56687
rect 11151 56631 11237 56687
rect 11293 56631 11379 56687
rect 11435 56631 11521 56687
rect 11577 56631 11663 56687
rect 11719 56631 11805 56687
rect 11861 56631 11947 56687
rect 12003 56631 12089 56687
rect 12145 56631 12231 56687
rect 12287 56631 12373 56687
rect 12429 56631 12515 56687
rect 12571 56631 12657 56687
rect 12713 56631 12799 56687
rect 12855 56631 12941 56687
rect 12997 56631 13083 56687
rect 13139 56631 13225 56687
rect 13281 56631 13367 56687
rect 13423 56631 13509 56687
rect 13565 56631 13651 56687
rect 13707 56631 13793 56687
rect 13849 56631 13935 56687
rect 13991 56631 14077 56687
rect 14133 56631 14219 56687
rect 14275 56631 14361 56687
rect 14417 56631 14503 56687
rect 14559 56631 14645 56687
rect 14701 56631 14787 56687
rect 14843 56631 15000 56687
rect 0 56545 15000 56631
rect 0 56489 161 56545
rect 217 56489 303 56545
rect 359 56489 445 56545
rect 501 56489 587 56545
rect 643 56489 729 56545
rect 785 56489 871 56545
rect 927 56489 1013 56545
rect 1069 56489 1155 56545
rect 1211 56489 1297 56545
rect 1353 56489 1439 56545
rect 1495 56489 1581 56545
rect 1637 56489 1723 56545
rect 1779 56489 1865 56545
rect 1921 56489 2007 56545
rect 2063 56489 2149 56545
rect 2205 56489 2291 56545
rect 2347 56489 2433 56545
rect 2489 56489 2575 56545
rect 2631 56489 2717 56545
rect 2773 56489 2859 56545
rect 2915 56489 3001 56545
rect 3057 56489 3143 56545
rect 3199 56489 3285 56545
rect 3341 56489 3427 56545
rect 3483 56489 3569 56545
rect 3625 56489 3711 56545
rect 3767 56489 3853 56545
rect 3909 56489 3995 56545
rect 4051 56489 4137 56545
rect 4193 56489 4279 56545
rect 4335 56489 4421 56545
rect 4477 56489 4563 56545
rect 4619 56489 4705 56545
rect 4761 56489 4847 56545
rect 4903 56489 4989 56545
rect 5045 56489 5131 56545
rect 5187 56489 5273 56545
rect 5329 56489 5415 56545
rect 5471 56489 5557 56545
rect 5613 56489 5699 56545
rect 5755 56489 5841 56545
rect 5897 56489 5983 56545
rect 6039 56489 6125 56545
rect 6181 56489 6267 56545
rect 6323 56489 6409 56545
rect 6465 56489 6551 56545
rect 6607 56489 6693 56545
rect 6749 56489 6835 56545
rect 6891 56489 6977 56545
rect 7033 56489 7119 56545
rect 7175 56489 7261 56545
rect 7317 56489 7403 56545
rect 7459 56489 7545 56545
rect 7601 56489 7687 56545
rect 7743 56489 7829 56545
rect 7885 56489 7971 56545
rect 8027 56489 8113 56545
rect 8169 56489 8255 56545
rect 8311 56489 8397 56545
rect 8453 56489 8539 56545
rect 8595 56489 8681 56545
rect 8737 56489 8823 56545
rect 8879 56489 8965 56545
rect 9021 56489 9107 56545
rect 9163 56489 9249 56545
rect 9305 56489 9391 56545
rect 9447 56489 9533 56545
rect 9589 56489 9675 56545
rect 9731 56489 9817 56545
rect 9873 56489 9959 56545
rect 10015 56489 10101 56545
rect 10157 56489 10243 56545
rect 10299 56489 10385 56545
rect 10441 56489 10527 56545
rect 10583 56489 10669 56545
rect 10725 56489 10811 56545
rect 10867 56489 10953 56545
rect 11009 56489 11095 56545
rect 11151 56489 11237 56545
rect 11293 56489 11379 56545
rect 11435 56489 11521 56545
rect 11577 56489 11663 56545
rect 11719 56489 11805 56545
rect 11861 56489 11947 56545
rect 12003 56489 12089 56545
rect 12145 56489 12231 56545
rect 12287 56489 12373 56545
rect 12429 56489 12515 56545
rect 12571 56489 12657 56545
rect 12713 56489 12799 56545
rect 12855 56489 12941 56545
rect 12997 56489 13083 56545
rect 13139 56489 13225 56545
rect 13281 56489 13367 56545
rect 13423 56489 13509 56545
rect 13565 56489 13651 56545
rect 13707 56489 13793 56545
rect 13849 56489 13935 56545
rect 13991 56489 14077 56545
rect 14133 56489 14219 56545
rect 14275 56489 14361 56545
rect 14417 56489 14503 56545
rect 14559 56489 14645 56545
rect 14701 56489 14787 56545
rect 14843 56489 15000 56545
rect 0 56403 15000 56489
rect 0 56347 161 56403
rect 217 56347 303 56403
rect 359 56347 445 56403
rect 501 56347 587 56403
rect 643 56347 729 56403
rect 785 56347 871 56403
rect 927 56347 1013 56403
rect 1069 56347 1155 56403
rect 1211 56347 1297 56403
rect 1353 56347 1439 56403
rect 1495 56347 1581 56403
rect 1637 56347 1723 56403
rect 1779 56347 1865 56403
rect 1921 56347 2007 56403
rect 2063 56347 2149 56403
rect 2205 56347 2291 56403
rect 2347 56347 2433 56403
rect 2489 56347 2575 56403
rect 2631 56347 2717 56403
rect 2773 56347 2859 56403
rect 2915 56347 3001 56403
rect 3057 56347 3143 56403
rect 3199 56347 3285 56403
rect 3341 56347 3427 56403
rect 3483 56347 3569 56403
rect 3625 56347 3711 56403
rect 3767 56347 3853 56403
rect 3909 56347 3995 56403
rect 4051 56347 4137 56403
rect 4193 56347 4279 56403
rect 4335 56347 4421 56403
rect 4477 56347 4563 56403
rect 4619 56347 4705 56403
rect 4761 56347 4847 56403
rect 4903 56347 4989 56403
rect 5045 56347 5131 56403
rect 5187 56347 5273 56403
rect 5329 56347 5415 56403
rect 5471 56347 5557 56403
rect 5613 56347 5699 56403
rect 5755 56347 5841 56403
rect 5897 56347 5983 56403
rect 6039 56347 6125 56403
rect 6181 56347 6267 56403
rect 6323 56347 6409 56403
rect 6465 56347 6551 56403
rect 6607 56347 6693 56403
rect 6749 56347 6835 56403
rect 6891 56347 6977 56403
rect 7033 56347 7119 56403
rect 7175 56347 7261 56403
rect 7317 56347 7403 56403
rect 7459 56347 7545 56403
rect 7601 56347 7687 56403
rect 7743 56347 7829 56403
rect 7885 56347 7971 56403
rect 8027 56347 8113 56403
rect 8169 56347 8255 56403
rect 8311 56347 8397 56403
rect 8453 56347 8539 56403
rect 8595 56347 8681 56403
rect 8737 56347 8823 56403
rect 8879 56347 8965 56403
rect 9021 56347 9107 56403
rect 9163 56347 9249 56403
rect 9305 56347 9391 56403
rect 9447 56347 9533 56403
rect 9589 56347 9675 56403
rect 9731 56347 9817 56403
rect 9873 56347 9959 56403
rect 10015 56347 10101 56403
rect 10157 56347 10243 56403
rect 10299 56347 10385 56403
rect 10441 56347 10527 56403
rect 10583 56347 10669 56403
rect 10725 56347 10811 56403
rect 10867 56347 10953 56403
rect 11009 56347 11095 56403
rect 11151 56347 11237 56403
rect 11293 56347 11379 56403
rect 11435 56347 11521 56403
rect 11577 56347 11663 56403
rect 11719 56347 11805 56403
rect 11861 56347 11947 56403
rect 12003 56347 12089 56403
rect 12145 56347 12231 56403
rect 12287 56347 12373 56403
rect 12429 56347 12515 56403
rect 12571 56347 12657 56403
rect 12713 56347 12799 56403
rect 12855 56347 12941 56403
rect 12997 56347 13083 56403
rect 13139 56347 13225 56403
rect 13281 56347 13367 56403
rect 13423 56347 13509 56403
rect 13565 56347 13651 56403
rect 13707 56347 13793 56403
rect 13849 56347 13935 56403
rect 13991 56347 14077 56403
rect 14133 56347 14219 56403
rect 14275 56347 14361 56403
rect 14417 56347 14503 56403
rect 14559 56347 14645 56403
rect 14701 56347 14787 56403
rect 14843 56347 15000 56403
rect 0 56261 15000 56347
rect 0 56205 161 56261
rect 217 56205 303 56261
rect 359 56205 445 56261
rect 501 56205 587 56261
rect 643 56205 729 56261
rect 785 56205 871 56261
rect 927 56205 1013 56261
rect 1069 56205 1155 56261
rect 1211 56205 1297 56261
rect 1353 56205 1439 56261
rect 1495 56205 1581 56261
rect 1637 56205 1723 56261
rect 1779 56205 1865 56261
rect 1921 56205 2007 56261
rect 2063 56205 2149 56261
rect 2205 56205 2291 56261
rect 2347 56205 2433 56261
rect 2489 56205 2575 56261
rect 2631 56205 2717 56261
rect 2773 56205 2859 56261
rect 2915 56205 3001 56261
rect 3057 56205 3143 56261
rect 3199 56205 3285 56261
rect 3341 56205 3427 56261
rect 3483 56205 3569 56261
rect 3625 56205 3711 56261
rect 3767 56205 3853 56261
rect 3909 56205 3995 56261
rect 4051 56205 4137 56261
rect 4193 56205 4279 56261
rect 4335 56205 4421 56261
rect 4477 56205 4563 56261
rect 4619 56205 4705 56261
rect 4761 56205 4847 56261
rect 4903 56205 4989 56261
rect 5045 56205 5131 56261
rect 5187 56205 5273 56261
rect 5329 56205 5415 56261
rect 5471 56205 5557 56261
rect 5613 56205 5699 56261
rect 5755 56205 5841 56261
rect 5897 56205 5983 56261
rect 6039 56205 6125 56261
rect 6181 56205 6267 56261
rect 6323 56205 6409 56261
rect 6465 56205 6551 56261
rect 6607 56205 6693 56261
rect 6749 56205 6835 56261
rect 6891 56205 6977 56261
rect 7033 56205 7119 56261
rect 7175 56205 7261 56261
rect 7317 56205 7403 56261
rect 7459 56205 7545 56261
rect 7601 56205 7687 56261
rect 7743 56205 7829 56261
rect 7885 56205 7971 56261
rect 8027 56205 8113 56261
rect 8169 56205 8255 56261
rect 8311 56205 8397 56261
rect 8453 56205 8539 56261
rect 8595 56205 8681 56261
rect 8737 56205 8823 56261
rect 8879 56205 8965 56261
rect 9021 56205 9107 56261
rect 9163 56205 9249 56261
rect 9305 56205 9391 56261
rect 9447 56205 9533 56261
rect 9589 56205 9675 56261
rect 9731 56205 9817 56261
rect 9873 56205 9959 56261
rect 10015 56205 10101 56261
rect 10157 56205 10243 56261
rect 10299 56205 10385 56261
rect 10441 56205 10527 56261
rect 10583 56205 10669 56261
rect 10725 56205 10811 56261
rect 10867 56205 10953 56261
rect 11009 56205 11095 56261
rect 11151 56205 11237 56261
rect 11293 56205 11379 56261
rect 11435 56205 11521 56261
rect 11577 56205 11663 56261
rect 11719 56205 11805 56261
rect 11861 56205 11947 56261
rect 12003 56205 12089 56261
rect 12145 56205 12231 56261
rect 12287 56205 12373 56261
rect 12429 56205 12515 56261
rect 12571 56205 12657 56261
rect 12713 56205 12799 56261
rect 12855 56205 12941 56261
rect 12997 56205 13083 56261
rect 13139 56205 13225 56261
rect 13281 56205 13367 56261
rect 13423 56205 13509 56261
rect 13565 56205 13651 56261
rect 13707 56205 13793 56261
rect 13849 56205 13935 56261
rect 13991 56205 14077 56261
rect 14133 56205 14219 56261
rect 14275 56205 14361 56261
rect 14417 56205 14503 56261
rect 14559 56205 14645 56261
rect 14701 56205 14787 56261
rect 14843 56205 15000 56261
rect 0 56119 15000 56205
rect 0 56063 161 56119
rect 217 56063 303 56119
rect 359 56063 445 56119
rect 501 56063 587 56119
rect 643 56063 729 56119
rect 785 56063 871 56119
rect 927 56063 1013 56119
rect 1069 56063 1155 56119
rect 1211 56063 1297 56119
rect 1353 56063 1439 56119
rect 1495 56063 1581 56119
rect 1637 56063 1723 56119
rect 1779 56063 1865 56119
rect 1921 56063 2007 56119
rect 2063 56063 2149 56119
rect 2205 56063 2291 56119
rect 2347 56063 2433 56119
rect 2489 56063 2575 56119
rect 2631 56063 2717 56119
rect 2773 56063 2859 56119
rect 2915 56063 3001 56119
rect 3057 56063 3143 56119
rect 3199 56063 3285 56119
rect 3341 56063 3427 56119
rect 3483 56063 3569 56119
rect 3625 56063 3711 56119
rect 3767 56063 3853 56119
rect 3909 56063 3995 56119
rect 4051 56063 4137 56119
rect 4193 56063 4279 56119
rect 4335 56063 4421 56119
rect 4477 56063 4563 56119
rect 4619 56063 4705 56119
rect 4761 56063 4847 56119
rect 4903 56063 4989 56119
rect 5045 56063 5131 56119
rect 5187 56063 5273 56119
rect 5329 56063 5415 56119
rect 5471 56063 5557 56119
rect 5613 56063 5699 56119
rect 5755 56063 5841 56119
rect 5897 56063 5983 56119
rect 6039 56063 6125 56119
rect 6181 56063 6267 56119
rect 6323 56063 6409 56119
rect 6465 56063 6551 56119
rect 6607 56063 6693 56119
rect 6749 56063 6835 56119
rect 6891 56063 6977 56119
rect 7033 56063 7119 56119
rect 7175 56063 7261 56119
rect 7317 56063 7403 56119
rect 7459 56063 7545 56119
rect 7601 56063 7687 56119
rect 7743 56063 7829 56119
rect 7885 56063 7971 56119
rect 8027 56063 8113 56119
rect 8169 56063 8255 56119
rect 8311 56063 8397 56119
rect 8453 56063 8539 56119
rect 8595 56063 8681 56119
rect 8737 56063 8823 56119
rect 8879 56063 8965 56119
rect 9021 56063 9107 56119
rect 9163 56063 9249 56119
rect 9305 56063 9391 56119
rect 9447 56063 9533 56119
rect 9589 56063 9675 56119
rect 9731 56063 9817 56119
rect 9873 56063 9959 56119
rect 10015 56063 10101 56119
rect 10157 56063 10243 56119
rect 10299 56063 10385 56119
rect 10441 56063 10527 56119
rect 10583 56063 10669 56119
rect 10725 56063 10811 56119
rect 10867 56063 10953 56119
rect 11009 56063 11095 56119
rect 11151 56063 11237 56119
rect 11293 56063 11379 56119
rect 11435 56063 11521 56119
rect 11577 56063 11663 56119
rect 11719 56063 11805 56119
rect 11861 56063 11947 56119
rect 12003 56063 12089 56119
rect 12145 56063 12231 56119
rect 12287 56063 12373 56119
rect 12429 56063 12515 56119
rect 12571 56063 12657 56119
rect 12713 56063 12799 56119
rect 12855 56063 12941 56119
rect 12997 56063 13083 56119
rect 13139 56063 13225 56119
rect 13281 56063 13367 56119
rect 13423 56063 13509 56119
rect 13565 56063 13651 56119
rect 13707 56063 13793 56119
rect 13849 56063 13935 56119
rect 13991 56063 14077 56119
rect 14133 56063 14219 56119
rect 14275 56063 14361 56119
rect 14417 56063 14503 56119
rect 14559 56063 14645 56119
rect 14701 56063 14787 56119
rect 14843 56063 15000 56119
rect 0 55977 15000 56063
rect 0 55921 161 55977
rect 217 55921 303 55977
rect 359 55921 445 55977
rect 501 55921 587 55977
rect 643 55921 729 55977
rect 785 55921 871 55977
rect 927 55921 1013 55977
rect 1069 55921 1155 55977
rect 1211 55921 1297 55977
rect 1353 55921 1439 55977
rect 1495 55921 1581 55977
rect 1637 55921 1723 55977
rect 1779 55921 1865 55977
rect 1921 55921 2007 55977
rect 2063 55921 2149 55977
rect 2205 55921 2291 55977
rect 2347 55921 2433 55977
rect 2489 55921 2575 55977
rect 2631 55921 2717 55977
rect 2773 55921 2859 55977
rect 2915 55921 3001 55977
rect 3057 55921 3143 55977
rect 3199 55921 3285 55977
rect 3341 55921 3427 55977
rect 3483 55921 3569 55977
rect 3625 55921 3711 55977
rect 3767 55921 3853 55977
rect 3909 55921 3995 55977
rect 4051 55921 4137 55977
rect 4193 55921 4279 55977
rect 4335 55921 4421 55977
rect 4477 55921 4563 55977
rect 4619 55921 4705 55977
rect 4761 55921 4847 55977
rect 4903 55921 4989 55977
rect 5045 55921 5131 55977
rect 5187 55921 5273 55977
rect 5329 55921 5415 55977
rect 5471 55921 5557 55977
rect 5613 55921 5699 55977
rect 5755 55921 5841 55977
rect 5897 55921 5983 55977
rect 6039 55921 6125 55977
rect 6181 55921 6267 55977
rect 6323 55921 6409 55977
rect 6465 55921 6551 55977
rect 6607 55921 6693 55977
rect 6749 55921 6835 55977
rect 6891 55921 6977 55977
rect 7033 55921 7119 55977
rect 7175 55921 7261 55977
rect 7317 55921 7403 55977
rect 7459 55921 7545 55977
rect 7601 55921 7687 55977
rect 7743 55921 7829 55977
rect 7885 55921 7971 55977
rect 8027 55921 8113 55977
rect 8169 55921 8255 55977
rect 8311 55921 8397 55977
rect 8453 55921 8539 55977
rect 8595 55921 8681 55977
rect 8737 55921 8823 55977
rect 8879 55921 8965 55977
rect 9021 55921 9107 55977
rect 9163 55921 9249 55977
rect 9305 55921 9391 55977
rect 9447 55921 9533 55977
rect 9589 55921 9675 55977
rect 9731 55921 9817 55977
rect 9873 55921 9959 55977
rect 10015 55921 10101 55977
rect 10157 55921 10243 55977
rect 10299 55921 10385 55977
rect 10441 55921 10527 55977
rect 10583 55921 10669 55977
rect 10725 55921 10811 55977
rect 10867 55921 10953 55977
rect 11009 55921 11095 55977
rect 11151 55921 11237 55977
rect 11293 55921 11379 55977
rect 11435 55921 11521 55977
rect 11577 55921 11663 55977
rect 11719 55921 11805 55977
rect 11861 55921 11947 55977
rect 12003 55921 12089 55977
rect 12145 55921 12231 55977
rect 12287 55921 12373 55977
rect 12429 55921 12515 55977
rect 12571 55921 12657 55977
rect 12713 55921 12799 55977
rect 12855 55921 12941 55977
rect 12997 55921 13083 55977
rect 13139 55921 13225 55977
rect 13281 55921 13367 55977
rect 13423 55921 13509 55977
rect 13565 55921 13651 55977
rect 13707 55921 13793 55977
rect 13849 55921 13935 55977
rect 13991 55921 14077 55977
rect 14133 55921 14219 55977
rect 14275 55921 14361 55977
rect 14417 55921 14503 55977
rect 14559 55921 14645 55977
rect 14701 55921 14787 55977
rect 14843 55921 15000 55977
rect 0 55835 15000 55921
rect 0 55779 161 55835
rect 217 55779 303 55835
rect 359 55779 445 55835
rect 501 55779 587 55835
rect 643 55779 729 55835
rect 785 55779 871 55835
rect 927 55779 1013 55835
rect 1069 55779 1155 55835
rect 1211 55779 1297 55835
rect 1353 55779 1439 55835
rect 1495 55779 1581 55835
rect 1637 55779 1723 55835
rect 1779 55779 1865 55835
rect 1921 55779 2007 55835
rect 2063 55779 2149 55835
rect 2205 55779 2291 55835
rect 2347 55779 2433 55835
rect 2489 55779 2575 55835
rect 2631 55779 2717 55835
rect 2773 55779 2859 55835
rect 2915 55779 3001 55835
rect 3057 55779 3143 55835
rect 3199 55779 3285 55835
rect 3341 55779 3427 55835
rect 3483 55779 3569 55835
rect 3625 55779 3711 55835
rect 3767 55779 3853 55835
rect 3909 55779 3995 55835
rect 4051 55779 4137 55835
rect 4193 55779 4279 55835
rect 4335 55779 4421 55835
rect 4477 55779 4563 55835
rect 4619 55779 4705 55835
rect 4761 55779 4847 55835
rect 4903 55779 4989 55835
rect 5045 55779 5131 55835
rect 5187 55779 5273 55835
rect 5329 55779 5415 55835
rect 5471 55779 5557 55835
rect 5613 55779 5699 55835
rect 5755 55779 5841 55835
rect 5897 55779 5983 55835
rect 6039 55779 6125 55835
rect 6181 55779 6267 55835
rect 6323 55779 6409 55835
rect 6465 55779 6551 55835
rect 6607 55779 6693 55835
rect 6749 55779 6835 55835
rect 6891 55779 6977 55835
rect 7033 55779 7119 55835
rect 7175 55779 7261 55835
rect 7317 55779 7403 55835
rect 7459 55779 7545 55835
rect 7601 55779 7687 55835
rect 7743 55779 7829 55835
rect 7885 55779 7971 55835
rect 8027 55779 8113 55835
rect 8169 55779 8255 55835
rect 8311 55779 8397 55835
rect 8453 55779 8539 55835
rect 8595 55779 8681 55835
rect 8737 55779 8823 55835
rect 8879 55779 8965 55835
rect 9021 55779 9107 55835
rect 9163 55779 9249 55835
rect 9305 55779 9391 55835
rect 9447 55779 9533 55835
rect 9589 55779 9675 55835
rect 9731 55779 9817 55835
rect 9873 55779 9959 55835
rect 10015 55779 10101 55835
rect 10157 55779 10243 55835
rect 10299 55779 10385 55835
rect 10441 55779 10527 55835
rect 10583 55779 10669 55835
rect 10725 55779 10811 55835
rect 10867 55779 10953 55835
rect 11009 55779 11095 55835
rect 11151 55779 11237 55835
rect 11293 55779 11379 55835
rect 11435 55779 11521 55835
rect 11577 55779 11663 55835
rect 11719 55779 11805 55835
rect 11861 55779 11947 55835
rect 12003 55779 12089 55835
rect 12145 55779 12231 55835
rect 12287 55779 12373 55835
rect 12429 55779 12515 55835
rect 12571 55779 12657 55835
rect 12713 55779 12799 55835
rect 12855 55779 12941 55835
rect 12997 55779 13083 55835
rect 13139 55779 13225 55835
rect 13281 55779 13367 55835
rect 13423 55779 13509 55835
rect 13565 55779 13651 55835
rect 13707 55779 13793 55835
rect 13849 55779 13935 55835
rect 13991 55779 14077 55835
rect 14133 55779 14219 55835
rect 14275 55779 14361 55835
rect 14417 55779 14503 55835
rect 14559 55779 14645 55835
rect 14701 55779 14787 55835
rect 14843 55779 15000 55835
rect 0 55693 15000 55779
rect 0 55637 161 55693
rect 217 55637 303 55693
rect 359 55637 445 55693
rect 501 55637 587 55693
rect 643 55637 729 55693
rect 785 55637 871 55693
rect 927 55637 1013 55693
rect 1069 55637 1155 55693
rect 1211 55637 1297 55693
rect 1353 55637 1439 55693
rect 1495 55637 1581 55693
rect 1637 55637 1723 55693
rect 1779 55637 1865 55693
rect 1921 55637 2007 55693
rect 2063 55637 2149 55693
rect 2205 55637 2291 55693
rect 2347 55637 2433 55693
rect 2489 55637 2575 55693
rect 2631 55637 2717 55693
rect 2773 55637 2859 55693
rect 2915 55637 3001 55693
rect 3057 55637 3143 55693
rect 3199 55637 3285 55693
rect 3341 55637 3427 55693
rect 3483 55637 3569 55693
rect 3625 55637 3711 55693
rect 3767 55637 3853 55693
rect 3909 55637 3995 55693
rect 4051 55637 4137 55693
rect 4193 55637 4279 55693
rect 4335 55637 4421 55693
rect 4477 55637 4563 55693
rect 4619 55637 4705 55693
rect 4761 55637 4847 55693
rect 4903 55637 4989 55693
rect 5045 55637 5131 55693
rect 5187 55637 5273 55693
rect 5329 55637 5415 55693
rect 5471 55637 5557 55693
rect 5613 55637 5699 55693
rect 5755 55637 5841 55693
rect 5897 55637 5983 55693
rect 6039 55637 6125 55693
rect 6181 55637 6267 55693
rect 6323 55637 6409 55693
rect 6465 55637 6551 55693
rect 6607 55637 6693 55693
rect 6749 55637 6835 55693
rect 6891 55637 6977 55693
rect 7033 55637 7119 55693
rect 7175 55637 7261 55693
rect 7317 55637 7403 55693
rect 7459 55637 7545 55693
rect 7601 55637 7687 55693
rect 7743 55637 7829 55693
rect 7885 55637 7971 55693
rect 8027 55637 8113 55693
rect 8169 55637 8255 55693
rect 8311 55637 8397 55693
rect 8453 55637 8539 55693
rect 8595 55637 8681 55693
rect 8737 55637 8823 55693
rect 8879 55637 8965 55693
rect 9021 55637 9107 55693
rect 9163 55637 9249 55693
rect 9305 55637 9391 55693
rect 9447 55637 9533 55693
rect 9589 55637 9675 55693
rect 9731 55637 9817 55693
rect 9873 55637 9959 55693
rect 10015 55637 10101 55693
rect 10157 55637 10243 55693
rect 10299 55637 10385 55693
rect 10441 55637 10527 55693
rect 10583 55637 10669 55693
rect 10725 55637 10811 55693
rect 10867 55637 10953 55693
rect 11009 55637 11095 55693
rect 11151 55637 11237 55693
rect 11293 55637 11379 55693
rect 11435 55637 11521 55693
rect 11577 55637 11663 55693
rect 11719 55637 11805 55693
rect 11861 55637 11947 55693
rect 12003 55637 12089 55693
rect 12145 55637 12231 55693
rect 12287 55637 12373 55693
rect 12429 55637 12515 55693
rect 12571 55637 12657 55693
rect 12713 55637 12799 55693
rect 12855 55637 12941 55693
rect 12997 55637 13083 55693
rect 13139 55637 13225 55693
rect 13281 55637 13367 55693
rect 13423 55637 13509 55693
rect 13565 55637 13651 55693
rect 13707 55637 13793 55693
rect 13849 55637 13935 55693
rect 13991 55637 14077 55693
rect 14133 55637 14219 55693
rect 14275 55637 14361 55693
rect 14417 55637 14503 55693
rect 14559 55637 14645 55693
rect 14701 55637 14787 55693
rect 14843 55637 15000 55693
rect 0 55600 15000 55637
rect 937 55400 3937 55600
rect 4337 55400 7337 55600
rect 7737 55400 10737 55600
rect 11137 55400 14137 55600
rect 0 55363 15000 55400
rect 0 55307 161 55363
rect 217 55307 303 55363
rect 359 55307 445 55363
rect 501 55307 587 55363
rect 643 55307 729 55363
rect 785 55307 871 55363
rect 927 55307 1013 55363
rect 1069 55307 1155 55363
rect 1211 55307 1297 55363
rect 1353 55307 1439 55363
rect 1495 55307 1581 55363
rect 1637 55307 1723 55363
rect 1779 55307 1865 55363
rect 1921 55307 2007 55363
rect 2063 55307 2149 55363
rect 2205 55307 2291 55363
rect 2347 55307 2433 55363
rect 2489 55307 2575 55363
rect 2631 55307 2717 55363
rect 2773 55307 2859 55363
rect 2915 55307 3001 55363
rect 3057 55307 3143 55363
rect 3199 55307 3285 55363
rect 3341 55307 3427 55363
rect 3483 55307 3569 55363
rect 3625 55307 3711 55363
rect 3767 55307 3853 55363
rect 3909 55307 3995 55363
rect 4051 55307 4137 55363
rect 4193 55307 4279 55363
rect 4335 55307 4421 55363
rect 4477 55307 4563 55363
rect 4619 55307 4705 55363
rect 4761 55307 4847 55363
rect 4903 55307 4989 55363
rect 5045 55307 5131 55363
rect 5187 55307 5273 55363
rect 5329 55307 5415 55363
rect 5471 55307 5557 55363
rect 5613 55307 5699 55363
rect 5755 55307 5841 55363
rect 5897 55307 5983 55363
rect 6039 55307 6125 55363
rect 6181 55307 6267 55363
rect 6323 55307 6409 55363
rect 6465 55307 6551 55363
rect 6607 55307 6693 55363
rect 6749 55307 6835 55363
rect 6891 55307 6977 55363
rect 7033 55307 7119 55363
rect 7175 55307 7261 55363
rect 7317 55307 7403 55363
rect 7459 55307 7545 55363
rect 7601 55307 7687 55363
rect 7743 55307 7829 55363
rect 7885 55307 7971 55363
rect 8027 55307 8113 55363
rect 8169 55307 8255 55363
rect 8311 55307 8397 55363
rect 8453 55307 8539 55363
rect 8595 55307 8681 55363
rect 8737 55307 8823 55363
rect 8879 55307 8965 55363
rect 9021 55307 9107 55363
rect 9163 55307 9249 55363
rect 9305 55307 9391 55363
rect 9447 55307 9533 55363
rect 9589 55307 9675 55363
rect 9731 55307 9817 55363
rect 9873 55307 9959 55363
rect 10015 55307 10101 55363
rect 10157 55307 10243 55363
rect 10299 55307 10385 55363
rect 10441 55307 10527 55363
rect 10583 55307 10669 55363
rect 10725 55307 10811 55363
rect 10867 55307 10953 55363
rect 11009 55307 11095 55363
rect 11151 55307 11237 55363
rect 11293 55307 11379 55363
rect 11435 55307 11521 55363
rect 11577 55307 11663 55363
rect 11719 55307 11805 55363
rect 11861 55307 11947 55363
rect 12003 55307 12089 55363
rect 12145 55307 12231 55363
rect 12287 55307 12373 55363
rect 12429 55307 12515 55363
rect 12571 55307 12657 55363
rect 12713 55307 12799 55363
rect 12855 55307 12941 55363
rect 12997 55307 13083 55363
rect 13139 55307 13225 55363
rect 13281 55307 13367 55363
rect 13423 55307 13509 55363
rect 13565 55307 13651 55363
rect 13707 55307 13793 55363
rect 13849 55307 13935 55363
rect 13991 55307 14077 55363
rect 14133 55307 14219 55363
rect 14275 55307 14361 55363
rect 14417 55307 14503 55363
rect 14559 55307 14645 55363
rect 14701 55307 14787 55363
rect 14843 55307 15000 55363
rect 0 55221 15000 55307
rect 0 55165 161 55221
rect 217 55165 303 55221
rect 359 55165 445 55221
rect 501 55165 587 55221
rect 643 55165 729 55221
rect 785 55165 871 55221
rect 927 55165 1013 55221
rect 1069 55165 1155 55221
rect 1211 55165 1297 55221
rect 1353 55165 1439 55221
rect 1495 55165 1581 55221
rect 1637 55165 1723 55221
rect 1779 55165 1865 55221
rect 1921 55165 2007 55221
rect 2063 55165 2149 55221
rect 2205 55165 2291 55221
rect 2347 55165 2433 55221
rect 2489 55165 2575 55221
rect 2631 55165 2717 55221
rect 2773 55165 2859 55221
rect 2915 55165 3001 55221
rect 3057 55165 3143 55221
rect 3199 55165 3285 55221
rect 3341 55165 3427 55221
rect 3483 55165 3569 55221
rect 3625 55165 3711 55221
rect 3767 55165 3853 55221
rect 3909 55165 3995 55221
rect 4051 55165 4137 55221
rect 4193 55165 4279 55221
rect 4335 55165 4421 55221
rect 4477 55165 4563 55221
rect 4619 55165 4705 55221
rect 4761 55165 4847 55221
rect 4903 55165 4989 55221
rect 5045 55165 5131 55221
rect 5187 55165 5273 55221
rect 5329 55165 5415 55221
rect 5471 55165 5557 55221
rect 5613 55165 5699 55221
rect 5755 55165 5841 55221
rect 5897 55165 5983 55221
rect 6039 55165 6125 55221
rect 6181 55165 6267 55221
rect 6323 55165 6409 55221
rect 6465 55165 6551 55221
rect 6607 55165 6693 55221
rect 6749 55165 6835 55221
rect 6891 55165 6977 55221
rect 7033 55165 7119 55221
rect 7175 55165 7261 55221
rect 7317 55165 7403 55221
rect 7459 55165 7545 55221
rect 7601 55165 7687 55221
rect 7743 55165 7829 55221
rect 7885 55165 7971 55221
rect 8027 55165 8113 55221
rect 8169 55165 8255 55221
rect 8311 55165 8397 55221
rect 8453 55165 8539 55221
rect 8595 55165 8681 55221
rect 8737 55165 8823 55221
rect 8879 55165 8965 55221
rect 9021 55165 9107 55221
rect 9163 55165 9249 55221
rect 9305 55165 9391 55221
rect 9447 55165 9533 55221
rect 9589 55165 9675 55221
rect 9731 55165 9817 55221
rect 9873 55165 9959 55221
rect 10015 55165 10101 55221
rect 10157 55165 10243 55221
rect 10299 55165 10385 55221
rect 10441 55165 10527 55221
rect 10583 55165 10669 55221
rect 10725 55165 10811 55221
rect 10867 55165 10953 55221
rect 11009 55165 11095 55221
rect 11151 55165 11237 55221
rect 11293 55165 11379 55221
rect 11435 55165 11521 55221
rect 11577 55165 11663 55221
rect 11719 55165 11805 55221
rect 11861 55165 11947 55221
rect 12003 55165 12089 55221
rect 12145 55165 12231 55221
rect 12287 55165 12373 55221
rect 12429 55165 12515 55221
rect 12571 55165 12657 55221
rect 12713 55165 12799 55221
rect 12855 55165 12941 55221
rect 12997 55165 13083 55221
rect 13139 55165 13225 55221
rect 13281 55165 13367 55221
rect 13423 55165 13509 55221
rect 13565 55165 13651 55221
rect 13707 55165 13793 55221
rect 13849 55165 13935 55221
rect 13991 55165 14077 55221
rect 14133 55165 14219 55221
rect 14275 55165 14361 55221
rect 14417 55165 14503 55221
rect 14559 55165 14645 55221
rect 14701 55165 14787 55221
rect 14843 55165 15000 55221
rect 0 55079 15000 55165
rect 0 55023 161 55079
rect 217 55023 303 55079
rect 359 55023 445 55079
rect 501 55023 587 55079
rect 643 55023 729 55079
rect 785 55023 871 55079
rect 927 55023 1013 55079
rect 1069 55023 1155 55079
rect 1211 55023 1297 55079
rect 1353 55023 1439 55079
rect 1495 55023 1581 55079
rect 1637 55023 1723 55079
rect 1779 55023 1865 55079
rect 1921 55023 2007 55079
rect 2063 55023 2149 55079
rect 2205 55023 2291 55079
rect 2347 55023 2433 55079
rect 2489 55023 2575 55079
rect 2631 55023 2717 55079
rect 2773 55023 2859 55079
rect 2915 55023 3001 55079
rect 3057 55023 3143 55079
rect 3199 55023 3285 55079
rect 3341 55023 3427 55079
rect 3483 55023 3569 55079
rect 3625 55023 3711 55079
rect 3767 55023 3853 55079
rect 3909 55023 3995 55079
rect 4051 55023 4137 55079
rect 4193 55023 4279 55079
rect 4335 55023 4421 55079
rect 4477 55023 4563 55079
rect 4619 55023 4705 55079
rect 4761 55023 4847 55079
rect 4903 55023 4989 55079
rect 5045 55023 5131 55079
rect 5187 55023 5273 55079
rect 5329 55023 5415 55079
rect 5471 55023 5557 55079
rect 5613 55023 5699 55079
rect 5755 55023 5841 55079
rect 5897 55023 5983 55079
rect 6039 55023 6125 55079
rect 6181 55023 6267 55079
rect 6323 55023 6409 55079
rect 6465 55023 6551 55079
rect 6607 55023 6693 55079
rect 6749 55023 6835 55079
rect 6891 55023 6977 55079
rect 7033 55023 7119 55079
rect 7175 55023 7261 55079
rect 7317 55023 7403 55079
rect 7459 55023 7545 55079
rect 7601 55023 7687 55079
rect 7743 55023 7829 55079
rect 7885 55023 7971 55079
rect 8027 55023 8113 55079
rect 8169 55023 8255 55079
rect 8311 55023 8397 55079
rect 8453 55023 8539 55079
rect 8595 55023 8681 55079
rect 8737 55023 8823 55079
rect 8879 55023 8965 55079
rect 9021 55023 9107 55079
rect 9163 55023 9249 55079
rect 9305 55023 9391 55079
rect 9447 55023 9533 55079
rect 9589 55023 9675 55079
rect 9731 55023 9817 55079
rect 9873 55023 9959 55079
rect 10015 55023 10101 55079
rect 10157 55023 10243 55079
rect 10299 55023 10385 55079
rect 10441 55023 10527 55079
rect 10583 55023 10669 55079
rect 10725 55023 10811 55079
rect 10867 55023 10953 55079
rect 11009 55023 11095 55079
rect 11151 55023 11237 55079
rect 11293 55023 11379 55079
rect 11435 55023 11521 55079
rect 11577 55023 11663 55079
rect 11719 55023 11805 55079
rect 11861 55023 11947 55079
rect 12003 55023 12089 55079
rect 12145 55023 12231 55079
rect 12287 55023 12373 55079
rect 12429 55023 12515 55079
rect 12571 55023 12657 55079
rect 12713 55023 12799 55079
rect 12855 55023 12941 55079
rect 12997 55023 13083 55079
rect 13139 55023 13225 55079
rect 13281 55023 13367 55079
rect 13423 55023 13509 55079
rect 13565 55023 13651 55079
rect 13707 55023 13793 55079
rect 13849 55023 13935 55079
rect 13991 55023 14077 55079
rect 14133 55023 14219 55079
rect 14275 55023 14361 55079
rect 14417 55023 14503 55079
rect 14559 55023 14645 55079
rect 14701 55023 14787 55079
rect 14843 55023 15000 55079
rect 0 54937 15000 55023
rect 0 54881 161 54937
rect 217 54881 303 54937
rect 359 54881 445 54937
rect 501 54881 587 54937
rect 643 54881 729 54937
rect 785 54881 871 54937
rect 927 54881 1013 54937
rect 1069 54881 1155 54937
rect 1211 54881 1297 54937
rect 1353 54881 1439 54937
rect 1495 54881 1581 54937
rect 1637 54881 1723 54937
rect 1779 54881 1865 54937
rect 1921 54881 2007 54937
rect 2063 54881 2149 54937
rect 2205 54881 2291 54937
rect 2347 54881 2433 54937
rect 2489 54881 2575 54937
rect 2631 54881 2717 54937
rect 2773 54881 2859 54937
rect 2915 54881 3001 54937
rect 3057 54881 3143 54937
rect 3199 54881 3285 54937
rect 3341 54881 3427 54937
rect 3483 54881 3569 54937
rect 3625 54881 3711 54937
rect 3767 54881 3853 54937
rect 3909 54881 3995 54937
rect 4051 54881 4137 54937
rect 4193 54881 4279 54937
rect 4335 54881 4421 54937
rect 4477 54881 4563 54937
rect 4619 54881 4705 54937
rect 4761 54881 4847 54937
rect 4903 54881 4989 54937
rect 5045 54881 5131 54937
rect 5187 54881 5273 54937
rect 5329 54881 5415 54937
rect 5471 54881 5557 54937
rect 5613 54881 5699 54937
rect 5755 54881 5841 54937
rect 5897 54881 5983 54937
rect 6039 54881 6125 54937
rect 6181 54881 6267 54937
rect 6323 54881 6409 54937
rect 6465 54881 6551 54937
rect 6607 54881 6693 54937
rect 6749 54881 6835 54937
rect 6891 54881 6977 54937
rect 7033 54881 7119 54937
rect 7175 54881 7261 54937
rect 7317 54881 7403 54937
rect 7459 54881 7545 54937
rect 7601 54881 7687 54937
rect 7743 54881 7829 54937
rect 7885 54881 7971 54937
rect 8027 54881 8113 54937
rect 8169 54881 8255 54937
rect 8311 54881 8397 54937
rect 8453 54881 8539 54937
rect 8595 54881 8681 54937
rect 8737 54881 8823 54937
rect 8879 54881 8965 54937
rect 9021 54881 9107 54937
rect 9163 54881 9249 54937
rect 9305 54881 9391 54937
rect 9447 54881 9533 54937
rect 9589 54881 9675 54937
rect 9731 54881 9817 54937
rect 9873 54881 9959 54937
rect 10015 54881 10101 54937
rect 10157 54881 10243 54937
rect 10299 54881 10385 54937
rect 10441 54881 10527 54937
rect 10583 54881 10669 54937
rect 10725 54881 10811 54937
rect 10867 54881 10953 54937
rect 11009 54881 11095 54937
rect 11151 54881 11237 54937
rect 11293 54881 11379 54937
rect 11435 54881 11521 54937
rect 11577 54881 11663 54937
rect 11719 54881 11805 54937
rect 11861 54881 11947 54937
rect 12003 54881 12089 54937
rect 12145 54881 12231 54937
rect 12287 54881 12373 54937
rect 12429 54881 12515 54937
rect 12571 54881 12657 54937
rect 12713 54881 12799 54937
rect 12855 54881 12941 54937
rect 12997 54881 13083 54937
rect 13139 54881 13225 54937
rect 13281 54881 13367 54937
rect 13423 54881 13509 54937
rect 13565 54881 13651 54937
rect 13707 54881 13793 54937
rect 13849 54881 13935 54937
rect 13991 54881 14077 54937
rect 14133 54881 14219 54937
rect 14275 54881 14361 54937
rect 14417 54881 14503 54937
rect 14559 54881 14645 54937
rect 14701 54881 14787 54937
rect 14843 54881 15000 54937
rect 0 54795 15000 54881
rect 0 54739 161 54795
rect 217 54739 303 54795
rect 359 54739 445 54795
rect 501 54739 587 54795
rect 643 54739 729 54795
rect 785 54739 871 54795
rect 927 54739 1013 54795
rect 1069 54739 1155 54795
rect 1211 54739 1297 54795
rect 1353 54739 1439 54795
rect 1495 54739 1581 54795
rect 1637 54739 1723 54795
rect 1779 54739 1865 54795
rect 1921 54739 2007 54795
rect 2063 54739 2149 54795
rect 2205 54739 2291 54795
rect 2347 54739 2433 54795
rect 2489 54739 2575 54795
rect 2631 54739 2717 54795
rect 2773 54739 2859 54795
rect 2915 54739 3001 54795
rect 3057 54739 3143 54795
rect 3199 54739 3285 54795
rect 3341 54739 3427 54795
rect 3483 54739 3569 54795
rect 3625 54739 3711 54795
rect 3767 54739 3853 54795
rect 3909 54739 3995 54795
rect 4051 54739 4137 54795
rect 4193 54739 4279 54795
rect 4335 54739 4421 54795
rect 4477 54739 4563 54795
rect 4619 54739 4705 54795
rect 4761 54739 4847 54795
rect 4903 54739 4989 54795
rect 5045 54739 5131 54795
rect 5187 54739 5273 54795
rect 5329 54739 5415 54795
rect 5471 54739 5557 54795
rect 5613 54739 5699 54795
rect 5755 54739 5841 54795
rect 5897 54739 5983 54795
rect 6039 54739 6125 54795
rect 6181 54739 6267 54795
rect 6323 54739 6409 54795
rect 6465 54739 6551 54795
rect 6607 54739 6693 54795
rect 6749 54739 6835 54795
rect 6891 54739 6977 54795
rect 7033 54739 7119 54795
rect 7175 54739 7261 54795
rect 7317 54739 7403 54795
rect 7459 54739 7545 54795
rect 7601 54739 7687 54795
rect 7743 54739 7829 54795
rect 7885 54739 7971 54795
rect 8027 54739 8113 54795
rect 8169 54739 8255 54795
rect 8311 54739 8397 54795
rect 8453 54739 8539 54795
rect 8595 54739 8681 54795
rect 8737 54739 8823 54795
rect 8879 54739 8965 54795
rect 9021 54739 9107 54795
rect 9163 54739 9249 54795
rect 9305 54739 9391 54795
rect 9447 54739 9533 54795
rect 9589 54739 9675 54795
rect 9731 54739 9817 54795
rect 9873 54739 9959 54795
rect 10015 54739 10101 54795
rect 10157 54739 10243 54795
rect 10299 54739 10385 54795
rect 10441 54739 10527 54795
rect 10583 54739 10669 54795
rect 10725 54739 10811 54795
rect 10867 54739 10953 54795
rect 11009 54739 11095 54795
rect 11151 54739 11237 54795
rect 11293 54739 11379 54795
rect 11435 54739 11521 54795
rect 11577 54739 11663 54795
rect 11719 54739 11805 54795
rect 11861 54739 11947 54795
rect 12003 54739 12089 54795
rect 12145 54739 12231 54795
rect 12287 54739 12373 54795
rect 12429 54739 12515 54795
rect 12571 54739 12657 54795
rect 12713 54739 12799 54795
rect 12855 54739 12941 54795
rect 12997 54739 13083 54795
rect 13139 54739 13225 54795
rect 13281 54739 13367 54795
rect 13423 54739 13509 54795
rect 13565 54739 13651 54795
rect 13707 54739 13793 54795
rect 13849 54739 13935 54795
rect 13991 54739 14077 54795
rect 14133 54739 14219 54795
rect 14275 54739 14361 54795
rect 14417 54739 14503 54795
rect 14559 54739 14645 54795
rect 14701 54739 14787 54795
rect 14843 54739 15000 54795
rect 0 54653 15000 54739
rect 0 54597 161 54653
rect 217 54597 303 54653
rect 359 54597 445 54653
rect 501 54597 587 54653
rect 643 54597 729 54653
rect 785 54597 871 54653
rect 927 54597 1013 54653
rect 1069 54597 1155 54653
rect 1211 54597 1297 54653
rect 1353 54597 1439 54653
rect 1495 54597 1581 54653
rect 1637 54597 1723 54653
rect 1779 54597 1865 54653
rect 1921 54597 2007 54653
rect 2063 54597 2149 54653
rect 2205 54597 2291 54653
rect 2347 54597 2433 54653
rect 2489 54597 2575 54653
rect 2631 54597 2717 54653
rect 2773 54597 2859 54653
rect 2915 54597 3001 54653
rect 3057 54597 3143 54653
rect 3199 54597 3285 54653
rect 3341 54597 3427 54653
rect 3483 54597 3569 54653
rect 3625 54597 3711 54653
rect 3767 54597 3853 54653
rect 3909 54597 3995 54653
rect 4051 54597 4137 54653
rect 4193 54597 4279 54653
rect 4335 54597 4421 54653
rect 4477 54597 4563 54653
rect 4619 54597 4705 54653
rect 4761 54597 4847 54653
rect 4903 54597 4989 54653
rect 5045 54597 5131 54653
rect 5187 54597 5273 54653
rect 5329 54597 5415 54653
rect 5471 54597 5557 54653
rect 5613 54597 5699 54653
rect 5755 54597 5841 54653
rect 5897 54597 5983 54653
rect 6039 54597 6125 54653
rect 6181 54597 6267 54653
rect 6323 54597 6409 54653
rect 6465 54597 6551 54653
rect 6607 54597 6693 54653
rect 6749 54597 6835 54653
rect 6891 54597 6977 54653
rect 7033 54597 7119 54653
rect 7175 54597 7261 54653
rect 7317 54597 7403 54653
rect 7459 54597 7545 54653
rect 7601 54597 7687 54653
rect 7743 54597 7829 54653
rect 7885 54597 7971 54653
rect 8027 54597 8113 54653
rect 8169 54597 8255 54653
rect 8311 54597 8397 54653
rect 8453 54597 8539 54653
rect 8595 54597 8681 54653
rect 8737 54597 8823 54653
rect 8879 54597 8965 54653
rect 9021 54597 9107 54653
rect 9163 54597 9249 54653
rect 9305 54597 9391 54653
rect 9447 54597 9533 54653
rect 9589 54597 9675 54653
rect 9731 54597 9817 54653
rect 9873 54597 9959 54653
rect 10015 54597 10101 54653
rect 10157 54597 10243 54653
rect 10299 54597 10385 54653
rect 10441 54597 10527 54653
rect 10583 54597 10669 54653
rect 10725 54597 10811 54653
rect 10867 54597 10953 54653
rect 11009 54597 11095 54653
rect 11151 54597 11237 54653
rect 11293 54597 11379 54653
rect 11435 54597 11521 54653
rect 11577 54597 11663 54653
rect 11719 54597 11805 54653
rect 11861 54597 11947 54653
rect 12003 54597 12089 54653
rect 12145 54597 12231 54653
rect 12287 54597 12373 54653
rect 12429 54597 12515 54653
rect 12571 54597 12657 54653
rect 12713 54597 12799 54653
rect 12855 54597 12941 54653
rect 12997 54597 13083 54653
rect 13139 54597 13225 54653
rect 13281 54597 13367 54653
rect 13423 54597 13509 54653
rect 13565 54597 13651 54653
rect 13707 54597 13793 54653
rect 13849 54597 13935 54653
rect 13991 54597 14077 54653
rect 14133 54597 14219 54653
rect 14275 54597 14361 54653
rect 14417 54597 14503 54653
rect 14559 54597 14645 54653
rect 14701 54597 14787 54653
rect 14843 54597 15000 54653
rect 0 54511 15000 54597
rect 0 54455 161 54511
rect 217 54455 303 54511
rect 359 54455 445 54511
rect 501 54455 587 54511
rect 643 54455 729 54511
rect 785 54455 871 54511
rect 927 54455 1013 54511
rect 1069 54455 1155 54511
rect 1211 54455 1297 54511
rect 1353 54455 1439 54511
rect 1495 54455 1581 54511
rect 1637 54455 1723 54511
rect 1779 54455 1865 54511
rect 1921 54455 2007 54511
rect 2063 54455 2149 54511
rect 2205 54455 2291 54511
rect 2347 54455 2433 54511
rect 2489 54455 2575 54511
rect 2631 54455 2717 54511
rect 2773 54455 2859 54511
rect 2915 54455 3001 54511
rect 3057 54455 3143 54511
rect 3199 54455 3285 54511
rect 3341 54455 3427 54511
rect 3483 54455 3569 54511
rect 3625 54455 3711 54511
rect 3767 54455 3853 54511
rect 3909 54455 3995 54511
rect 4051 54455 4137 54511
rect 4193 54455 4279 54511
rect 4335 54455 4421 54511
rect 4477 54455 4563 54511
rect 4619 54455 4705 54511
rect 4761 54455 4847 54511
rect 4903 54455 4989 54511
rect 5045 54455 5131 54511
rect 5187 54455 5273 54511
rect 5329 54455 5415 54511
rect 5471 54455 5557 54511
rect 5613 54455 5699 54511
rect 5755 54455 5841 54511
rect 5897 54455 5983 54511
rect 6039 54455 6125 54511
rect 6181 54455 6267 54511
rect 6323 54455 6409 54511
rect 6465 54455 6551 54511
rect 6607 54455 6693 54511
rect 6749 54455 6835 54511
rect 6891 54455 6977 54511
rect 7033 54455 7119 54511
rect 7175 54455 7261 54511
rect 7317 54455 7403 54511
rect 7459 54455 7545 54511
rect 7601 54455 7687 54511
rect 7743 54455 7829 54511
rect 7885 54455 7971 54511
rect 8027 54455 8113 54511
rect 8169 54455 8255 54511
rect 8311 54455 8397 54511
rect 8453 54455 8539 54511
rect 8595 54455 8681 54511
rect 8737 54455 8823 54511
rect 8879 54455 8965 54511
rect 9021 54455 9107 54511
rect 9163 54455 9249 54511
rect 9305 54455 9391 54511
rect 9447 54455 9533 54511
rect 9589 54455 9675 54511
rect 9731 54455 9817 54511
rect 9873 54455 9959 54511
rect 10015 54455 10101 54511
rect 10157 54455 10243 54511
rect 10299 54455 10385 54511
rect 10441 54455 10527 54511
rect 10583 54455 10669 54511
rect 10725 54455 10811 54511
rect 10867 54455 10953 54511
rect 11009 54455 11095 54511
rect 11151 54455 11237 54511
rect 11293 54455 11379 54511
rect 11435 54455 11521 54511
rect 11577 54455 11663 54511
rect 11719 54455 11805 54511
rect 11861 54455 11947 54511
rect 12003 54455 12089 54511
rect 12145 54455 12231 54511
rect 12287 54455 12373 54511
rect 12429 54455 12515 54511
rect 12571 54455 12657 54511
rect 12713 54455 12799 54511
rect 12855 54455 12941 54511
rect 12997 54455 13083 54511
rect 13139 54455 13225 54511
rect 13281 54455 13367 54511
rect 13423 54455 13509 54511
rect 13565 54455 13651 54511
rect 13707 54455 13793 54511
rect 13849 54455 13935 54511
rect 13991 54455 14077 54511
rect 14133 54455 14219 54511
rect 14275 54455 14361 54511
rect 14417 54455 14503 54511
rect 14559 54455 14645 54511
rect 14701 54455 14787 54511
rect 14843 54455 15000 54511
rect 0 54369 15000 54455
rect 0 54313 161 54369
rect 217 54313 303 54369
rect 359 54313 445 54369
rect 501 54313 587 54369
rect 643 54313 729 54369
rect 785 54313 871 54369
rect 927 54313 1013 54369
rect 1069 54313 1155 54369
rect 1211 54313 1297 54369
rect 1353 54313 1439 54369
rect 1495 54313 1581 54369
rect 1637 54313 1723 54369
rect 1779 54313 1865 54369
rect 1921 54313 2007 54369
rect 2063 54313 2149 54369
rect 2205 54313 2291 54369
rect 2347 54313 2433 54369
rect 2489 54313 2575 54369
rect 2631 54313 2717 54369
rect 2773 54313 2859 54369
rect 2915 54313 3001 54369
rect 3057 54313 3143 54369
rect 3199 54313 3285 54369
rect 3341 54313 3427 54369
rect 3483 54313 3569 54369
rect 3625 54313 3711 54369
rect 3767 54313 3853 54369
rect 3909 54313 3995 54369
rect 4051 54313 4137 54369
rect 4193 54313 4279 54369
rect 4335 54313 4421 54369
rect 4477 54313 4563 54369
rect 4619 54313 4705 54369
rect 4761 54313 4847 54369
rect 4903 54313 4989 54369
rect 5045 54313 5131 54369
rect 5187 54313 5273 54369
rect 5329 54313 5415 54369
rect 5471 54313 5557 54369
rect 5613 54313 5699 54369
rect 5755 54313 5841 54369
rect 5897 54313 5983 54369
rect 6039 54313 6125 54369
rect 6181 54313 6267 54369
rect 6323 54313 6409 54369
rect 6465 54313 6551 54369
rect 6607 54313 6693 54369
rect 6749 54313 6835 54369
rect 6891 54313 6977 54369
rect 7033 54313 7119 54369
rect 7175 54313 7261 54369
rect 7317 54313 7403 54369
rect 7459 54313 7545 54369
rect 7601 54313 7687 54369
rect 7743 54313 7829 54369
rect 7885 54313 7971 54369
rect 8027 54313 8113 54369
rect 8169 54313 8255 54369
rect 8311 54313 8397 54369
rect 8453 54313 8539 54369
rect 8595 54313 8681 54369
rect 8737 54313 8823 54369
rect 8879 54313 8965 54369
rect 9021 54313 9107 54369
rect 9163 54313 9249 54369
rect 9305 54313 9391 54369
rect 9447 54313 9533 54369
rect 9589 54313 9675 54369
rect 9731 54313 9817 54369
rect 9873 54313 9959 54369
rect 10015 54313 10101 54369
rect 10157 54313 10243 54369
rect 10299 54313 10385 54369
rect 10441 54313 10527 54369
rect 10583 54313 10669 54369
rect 10725 54313 10811 54369
rect 10867 54313 10953 54369
rect 11009 54313 11095 54369
rect 11151 54313 11237 54369
rect 11293 54313 11379 54369
rect 11435 54313 11521 54369
rect 11577 54313 11663 54369
rect 11719 54313 11805 54369
rect 11861 54313 11947 54369
rect 12003 54313 12089 54369
rect 12145 54313 12231 54369
rect 12287 54313 12373 54369
rect 12429 54313 12515 54369
rect 12571 54313 12657 54369
rect 12713 54313 12799 54369
rect 12855 54313 12941 54369
rect 12997 54313 13083 54369
rect 13139 54313 13225 54369
rect 13281 54313 13367 54369
rect 13423 54313 13509 54369
rect 13565 54313 13651 54369
rect 13707 54313 13793 54369
rect 13849 54313 13935 54369
rect 13991 54313 14077 54369
rect 14133 54313 14219 54369
rect 14275 54313 14361 54369
rect 14417 54313 14503 54369
rect 14559 54313 14645 54369
rect 14701 54313 14787 54369
rect 14843 54313 15000 54369
rect 0 54227 15000 54313
rect 0 54171 161 54227
rect 217 54171 303 54227
rect 359 54171 445 54227
rect 501 54171 587 54227
rect 643 54171 729 54227
rect 785 54171 871 54227
rect 927 54171 1013 54227
rect 1069 54171 1155 54227
rect 1211 54171 1297 54227
rect 1353 54171 1439 54227
rect 1495 54171 1581 54227
rect 1637 54171 1723 54227
rect 1779 54171 1865 54227
rect 1921 54171 2007 54227
rect 2063 54171 2149 54227
rect 2205 54171 2291 54227
rect 2347 54171 2433 54227
rect 2489 54171 2575 54227
rect 2631 54171 2717 54227
rect 2773 54171 2859 54227
rect 2915 54171 3001 54227
rect 3057 54171 3143 54227
rect 3199 54171 3285 54227
rect 3341 54171 3427 54227
rect 3483 54171 3569 54227
rect 3625 54171 3711 54227
rect 3767 54171 3853 54227
rect 3909 54171 3995 54227
rect 4051 54171 4137 54227
rect 4193 54171 4279 54227
rect 4335 54171 4421 54227
rect 4477 54171 4563 54227
rect 4619 54171 4705 54227
rect 4761 54171 4847 54227
rect 4903 54171 4989 54227
rect 5045 54171 5131 54227
rect 5187 54171 5273 54227
rect 5329 54171 5415 54227
rect 5471 54171 5557 54227
rect 5613 54171 5699 54227
rect 5755 54171 5841 54227
rect 5897 54171 5983 54227
rect 6039 54171 6125 54227
rect 6181 54171 6267 54227
rect 6323 54171 6409 54227
rect 6465 54171 6551 54227
rect 6607 54171 6693 54227
rect 6749 54171 6835 54227
rect 6891 54171 6977 54227
rect 7033 54171 7119 54227
rect 7175 54171 7261 54227
rect 7317 54171 7403 54227
rect 7459 54171 7545 54227
rect 7601 54171 7687 54227
rect 7743 54171 7829 54227
rect 7885 54171 7971 54227
rect 8027 54171 8113 54227
rect 8169 54171 8255 54227
rect 8311 54171 8397 54227
rect 8453 54171 8539 54227
rect 8595 54171 8681 54227
rect 8737 54171 8823 54227
rect 8879 54171 8965 54227
rect 9021 54171 9107 54227
rect 9163 54171 9249 54227
rect 9305 54171 9391 54227
rect 9447 54171 9533 54227
rect 9589 54171 9675 54227
rect 9731 54171 9817 54227
rect 9873 54171 9959 54227
rect 10015 54171 10101 54227
rect 10157 54171 10243 54227
rect 10299 54171 10385 54227
rect 10441 54171 10527 54227
rect 10583 54171 10669 54227
rect 10725 54171 10811 54227
rect 10867 54171 10953 54227
rect 11009 54171 11095 54227
rect 11151 54171 11237 54227
rect 11293 54171 11379 54227
rect 11435 54171 11521 54227
rect 11577 54171 11663 54227
rect 11719 54171 11805 54227
rect 11861 54171 11947 54227
rect 12003 54171 12089 54227
rect 12145 54171 12231 54227
rect 12287 54171 12373 54227
rect 12429 54171 12515 54227
rect 12571 54171 12657 54227
rect 12713 54171 12799 54227
rect 12855 54171 12941 54227
rect 12997 54171 13083 54227
rect 13139 54171 13225 54227
rect 13281 54171 13367 54227
rect 13423 54171 13509 54227
rect 13565 54171 13651 54227
rect 13707 54171 13793 54227
rect 13849 54171 13935 54227
rect 13991 54171 14077 54227
rect 14133 54171 14219 54227
rect 14275 54171 14361 54227
rect 14417 54171 14503 54227
rect 14559 54171 14645 54227
rect 14701 54171 14787 54227
rect 14843 54171 15000 54227
rect 0 54085 15000 54171
rect 0 54029 161 54085
rect 217 54029 303 54085
rect 359 54029 445 54085
rect 501 54029 587 54085
rect 643 54029 729 54085
rect 785 54029 871 54085
rect 927 54029 1013 54085
rect 1069 54029 1155 54085
rect 1211 54029 1297 54085
rect 1353 54029 1439 54085
rect 1495 54029 1581 54085
rect 1637 54029 1723 54085
rect 1779 54029 1865 54085
rect 1921 54029 2007 54085
rect 2063 54029 2149 54085
rect 2205 54029 2291 54085
rect 2347 54029 2433 54085
rect 2489 54029 2575 54085
rect 2631 54029 2717 54085
rect 2773 54029 2859 54085
rect 2915 54029 3001 54085
rect 3057 54029 3143 54085
rect 3199 54029 3285 54085
rect 3341 54029 3427 54085
rect 3483 54029 3569 54085
rect 3625 54029 3711 54085
rect 3767 54029 3853 54085
rect 3909 54029 3995 54085
rect 4051 54029 4137 54085
rect 4193 54029 4279 54085
rect 4335 54029 4421 54085
rect 4477 54029 4563 54085
rect 4619 54029 4705 54085
rect 4761 54029 4847 54085
rect 4903 54029 4989 54085
rect 5045 54029 5131 54085
rect 5187 54029 5273 54085
rect 5329 54029 5415 54085
rect 5471 54029 5557 54085
rect 5613 54029 5699 54085
rect 5755 54029 5841 54085
rect 5897 54029 5983 54085
rect 6039 54029 6125 54085
rect 6181 54029 6267 54085
rect 6323 54029 6409 54085
rect 6465 54029 6551 54085
rect 6607 54029 6693 54085
rect 6749 54029 6835 54085
rect 6891 54029 6977 54085
rect 7033 54029 7119 54085
rect 7175 54029 7261 54085
rect 7317 54029 7403 54085
rect 7459 54029 7545 54085
rect 7601 54029 7687 54085
rect 7743 54029 7829 54085
rect 7885 54029 7971 54085
rect 8027 54029 8113 54085
rect 8169 54029 8255 54085
rect 8311 54029 8397 54085
rect 8453 54029 8539 54085
rect 8595 54029 8681 54085
rect 8737 54029 8823 54085
rect 8879 54029 8965 54085
rect 9021 54029 9107 54085
rect 9163 54029 9249 54085
rect 9305 54029 9391 54085
rect 9447 54029 9533 54085
rect 9589 54029 9675 54085
rect 9731 54029 9817 54085
rect 9873 54029 9959 54085
rect 10015 54029 10101 54085
rect 10157 54029 10243 54085
rect 10299 54029 10385 54085
rect 10441 54029 10527 54085
rect 10583 54029 10669 54085
rect 10725 54029 10811 54085
rect 10867 54029 10953 54085
rect 11009 54029 11095 54085
rect 11151 54029 11237 54085
rect 11293 54029 11379 54085
rect 11435 54029 11521 54085
rect 11577 54029 11663 54085
rect 11719 54029 11805 54085
rect 11861 54029 11947 54085
rect 12003 54029 12089 54085
rect 12145 54029 12231 54085
rect 12287 54029 12373 54085
rect 12429 54029 12515 54085
rect 12571 54029 12657 54085
rect 12713 54029 12799 54085
rect 12855 54029 12941 54085
rect 12997 54029 13083 54085
rect 13139 54029 13225 54085
rect 13281 54029 13367 54085
rect 13423 54029 13509 54085
rect 13565 54029 13651 54085
rect 13707 54029 13793 54085
rect 13849 54029 13935 54085
rect 13991 54029 14077 54085
rect 14133 54029 14219 54085
rect 14275 54029 14361 54085
rect 14417 54029 14503 54085
rect 14559 54029 14645 54085
rect 14701 54029 14787 54085
rect 14843 54029 15000 54085
rect 0 54000 15000 54029
rect 937 53800 3937 54000
rect 4337 53800 7337 54000
rect 7737 53800 10737 54000
rect 11137 53800 14137 54000
rect 0 53771 15000 53800
rect 0 53715 161 53771
rect 217 53715 303 53771
rect 359 53715 445 53771
rect 501 53715 587 53771
rect 643 53715 729 53771
rect 785 53715 871 53771
rect 927 53715 1013 53771
rect 1069 53715 1155 53771
rect 1211 53715 1297 53771
rect 1353 53715 1439 53771
rect 1495 53715 1581 53771
rect 1637 53715 1723 53771
rect 1779 53715 1865 53771
rect 1921 53715 2007 53771
rect 2063 53715 2149 53771
rect 2205 53715 2291 53771
rect 2347 53715 2433 53771
rect 2489 53715 2575 53771
rect 2631 53715 2717 53771
rect 2773 53715 2859 53771
rect 2915 53715 3001 53771
rect 3057 53715 3143 53771
rect 3199 53715 3285 53771
rect 3341 53715 3427 53771
rect 3483 53715 3569 53771
rect 3625 53715 3711 53771
rect 3767 53715 3853 53771
rect 3909 53715 3995 53771
rect 4051 53715 4137 53771
rect 4193 53715 4279 53771
rect 4335 53715 4421 53771
rect 4477 53715 4563 53771
rect 4619 53715 4705 53771
rect 4761 53715 4847 53771
rect 4903 53715 4989 53771
rect 5045 53715 5131 53771
rect 5187 53715 5273 53771
rect 5329 53715 5415 53771
rect 5471 53715 5557 53771
rect 5613 53715 5699 53771
rect 5755 53715 5841 53771
rect 5897 53715 5983 53771
rect 6039 53715 6125 53771
rect 6181 53715 6267 53771
rect 6323 53715 6409 53771
rect 6465 53715 6551 53771
rect 6607 53715 6693 53771
rect 6749 53715 6835 53771
rect 6891 53715 6977 53771
rect 7033 53715 7119 53771
rect 7175 53715 7261 53771
rect 7317 53715 7403 53771
rect 7459 53715 7545 53771
rect 7601 53715 7687 53771
rect 7743 53715 7829 53771
rect 7885 53715 7971 53771
rect 8027 53715 8113 53771
rect 8169 53715 8255 53771
rect 8311 53715 8397 53771
rect 8453 53715 8539 53771
rect 8595 53715 8681 53771
rect 8737 53715 8823 53771
rect 8879 53715 8965 53771
rect 9021 53715 9107 53771
rect 9163 53715 9249 53771
rect 9305 53715 9391 53771
rect 9447 53715 9533 53771
rect 9589 53715 9675 53771
rect 9731 53715 9817 53771
rect 9873 53715 9959 53771
rect 10015 53715 10101 53771
rect 10157 53715 10243 53771
rect 10299 53715 10385 53771
rect 10441 53715 10527 53771
rect 10583 53715 10669 53771
rect 10725 53715 10811 53771
rect 10867 53715 10953 53771
rect 11009 53715 11095 53771
rect 11151 53715 11237 53771
rect 11293 53715 11379 53771
rect 11435 53715 11521 53771
rect 11577 53715 11663 53771
rect 11719 53715 11805 53771
rect 11861 53715 11947 53771
rect 12003 53715 12089 53771
rect 12145 53715 12231 53771
rect 12287 53715 12373 53771
rect 12429 53715 12515 53771
rect 12571 53715 12657 53771
rect 12713 53715 12799 53771
rect 12855 53715 12941 53771
rect 12997 53715 13083 53771
rect 13139 53715 13225 53771
rect 13281 53715 13367 53771
rect 13423 53715 13509 53771
rect 13565 53715 13651 53771
rect 13707 53715 13793 53771
rect 13849 53715 13935 53771
rect 13991 53715 14077 53771
rect 14133 53715 14219 53771
rect 14275 53715 14361 53771
rect 14417 53715 14503 53771
rect 14559 53715 14645 53771
rect 14701 53715 14787 53771
rect 14843 53715 15000 53771
rect 0 53629 15000 53715
rect 0 53573 161 53629
rect 217 53573 303 53629
rect 359 53573 445 53629
rect 501 53573 587 53629
rect 643 53573 729 53629
rect 785 53573 871 53629
rect 927 53573 1013 53629
rect 1069 53573 1155 53629
rect 1211 53573 1297 53629
rect 1353 53573 1439 53629
rect 1495 53573 1581 53629
rect 1637 53573 1723 53629
rect 1779 53573 1865 53629
rect 1921 53573 2007 53629
rect 2063 53573 2149 53629
rect 2205 53573 2291 53629
rect 2347 53573 2433 53629
rect 2489 53573 2575 53629
rect 2631 53573 2717 53629
rect 2773 53573 2859 53629
rect 2915 53573 3001 53629
rect 3057 53573 3143 53629
rect 3199 53573 3285 53629
rect 3341 53573 3427 53629
rect 3483 53573 3569 53629
rect 3625 53573 3711 53629
rect 3767 53573 3853 53629
rect 3909 53573 3995 53629
rect 4051 53573 4137 53629
rect 4193 53573 4279 53629
rect 4335 53573 4421 53629
rect 4477 53573 4563 53629
rect 4619 53573 4705 53629
rect 4761 53573 4847 53629
rect 4903 53573 4989 53629
rect 5045 53573 5131 53629
rect 5187 53573 5273 53629
rect 5329 53573 5415 53629
rect 5471 53573 5557 53629
rect 5613 53573 5699 53629
rect 5755 53573 5841 53629
rect 5897 53573 5983 53629
rect 6039 53573 6125 53629
rect 6181 53573 6267 53629
rect 6323 53573 6409 53629
rect 6465 53573 6551 53629
rect 6607 53573 6693 53629
rect 6749 53573 6835 53629
rect 6891 53573 6977 53629
rect 7033 53573 7119 53629
rect 7175 53573 7261 53629
rect 7317 53573 7403 53629
rect 7459 53573 7545 53629
rect 7601 53573 7687 53629
rect 7743 53573 7829 53629
rect 7885 53573 7971 53629
rect 8027 53573 8113 53629
rect 8169 53573 8255 53629
rect 8311 53573 8397 53629
rect 8453 53573 8539 53629
rect 8595 53573 8681 53629
rect 8737 53573 8823 53629
rect 8879 53573 8965 53629
rect 9021 53573 9107 53629
rect 9163 53573 9249 53629
rect 9305 53573 9391 53629
rect 9447 53573 9533 53629
rect 9589 53573 9675 53629
rect 9731 53573 9817 53629
rect 9873 53573 9959 53629
rect 10015 53573 10101 53629
rect 10157 53573 10243 53629
rect 10299 53573 10385 53629
rect 10441 53573 10527 53629
rect 10583 53573 10669 53629
rect 10725 53573 10811 53629
rect 10867 53573 10953 53629
rect 11009 53573 11095 53629
rect 11151 53573 11237 53629
rect 11293 53573 11379 53629
rect 11435 53573 11521 53629
rect 11577 53573 11663 53629
rect 11719 53573 11805 53629
rect 11861 53573 11947 53629
rect 12003 53573 12089 53629
rect 12145 53573 12231 53629
rect 12287 53573 12373 53629
rect 12429 53573 12515 53629
rect 12571 53573 12657 53629
rect 12713 53573 12799 53629
rect 12855 53573 12941 53629
rect 12997 53573 13083 53629
rect 13139 53573 13225 53629
rect 13281 53573 13367 53629
rect 13423 53573 13509 53629
rect 13565 53573 13651 53629
rect 13707 53573 13793 53629
rect 13849 53573 13935 53629
rect 13991 53573 14077 53629
rect 14133 53573 14219 53629
rect 14275 53573 14361 53629
rect 14417 53573 14503 53629
rect 14559 53573 14645 53629
rect 14701 53573 14787 53629
rect 14843 53573 15000 53629
rect 0 53487 15000 53573
rect 0 53431 161 53487
rect 217 53431 303 53487
rect 359 53431 445 53487
rect 501 53431 587 53487
rect 643 53431 729 53487
rect 785 53431 871 53487
rect 927 53431 1013 53487
rect 1069 53431 1155 53487
rect 1211 53431 1297 53487
rect 1353 53431 1439 53487
rect 1495 53431 1581 53487
rect 1637 53431 1723 53487
rect 1779 53431 1865 53487
rect 1921 53431 2007 53487
rect 2063 53431 2149 53487
rect 2205 53431 2291 53487
rect 2347 53431 2433 53487
rect 2489 53431 2575 53487
rect 2631 53431 2717 53487
rect 2773 53431 2859 53487
rect 2915 53431 3001 53487
rect 3057 53431 3143 53487
rect 3199 53431 3285 53487
rect 3341 53431 3427 53487
rect 3483 53431 3569 53487
rect 3625 53431 3711 53487
rect 3767 53431 3853 53487
rect 3909 53431 3995 53487
rect 4051 53431 4137 53487
rect 4193 53431 4279 53487
rect 4335 53431 4421 53487
rect 4477 53431 4563 53487
rect 4619 53431 4705 53487
rect 4761 53431 4847 53487
rect 4903 53431 4989 53487
rect 5045 53431 5131 53487
rect 5187 53431 5273 53487
rect 5329 53431 5415 53487
rect 5471 53431 5557 53487
rect 5613 53431 5699 53487
rect 5755 53431 5841 53487
rect 5897 53431 5983 53487
rect 6039 53431 6125 53487
rect 6181 53431 6267 53487
rect 6323 53431 6409 53487
rect 6465 53431 6551 53487
rect 6607 53431 6693 53487
rect 6749 53431 6835 53487
rect 6891 53431 6977 53487
rect 7033 53431 7119 53487
rect 7175 53431 7261 53487
rect 7317 53431 7403 53487
rect 7459 53431 7545 53487
rect 7601 53431 7687 53487
rect 7743 53431 7829 53487
rect 7885 53431 7971 53487
rect 8027 53431 8113 53487
rect 8169 53431 8255 53487
rect 8311 53431 8397 53487
rect 8453 53431 8539 53487
rect 8595 53431 8681 53487
rect 8737 53431 8823 53487
rect 8879 53431 8965 53487
rect 9021 53431 9107 53487
rect 9163 53431 9249 53487
rect 9305 53431 9391 53487
rect 9447 53431 9533 53487
rect 9589 53431 9675 53487
rect 9731 53431 9817 53487
rect 9873 53431 9959 53487
rect 10015 53431 10101 53487
rect 10157 53431 10243 53487
rect 10299 53431 10385 53487
rect 10441 53431 10527 53487
rect 10583 53431 10669 53487
rect 10725 53431 10811 53487
rect 10867 53431 10953 53487
rect 11009 53431 11095 53487
rect 11151 53431 11237 53487
rect 11293 53431 11379 53487
rect 11435 53431 11521 53487
rect 11577 53431 11663 53487
rect 11719 53431 11805 53487
rect 11861 53431 11947 53487
rect 12003 53431 12089 53487
rect 12145 53431 12231 53487
rect 12287 53431 12373 53487
rect 12429 53431 12515 53487
rect 12571 53431 12657 53487
rect 12713 53431 12799 53487
rect 12855 53431 12941 53487
rect 12997 53431 13083 53487
rect 13139 53431 13225 53487
rect 13281 53431 13367 53487
rect 13423 53431 13509 53487
rect 13565 53431 13651 53487
rect 13707 53431 13793 53487
rect 13849 53431 13935 53487
rect 13991 53431 14077 53487
rect 14133 53431 14219 53487
rect 14275 53431 14361 53487
rect 14417 53431 14503 53487
rect 14559 53431 14645 53487
rect 14701 53431 14787 53487
rect 14843 53431 15000 53487
rect 0 53345 15000 53431
rect 0 53289 161 53345
rect 217 53289 303 53345
rect 359 53289 445 53345
rect 501 53289 587 53345
rect 643 53289 729 53345
rect 785 53289 871 53345
rect 927 53289 1013 53345
rect 1069 53289 1155 53345
rect 1211 53289 1297 53345
rect 1353 53289 1439 53345
rect 1495 53289 1581 53345
rect 1637 53289 1723 53345
rect 1779 53289 1865 53345
rect 1921 53289 2007 53345
rect 2063 53289 2149 53345
rect 2205 53289 2291 53345
rect 2347 53289 2433 53345
rect 2489 53289 2575 53345
rect 2631 53289 2717 53345
rect 2773 53289 2859 53345
rect 2915 53289 3001 53345
rect 3057 53289 3143 53345
rect 3199 53289 3285 53345
rect 3341 53289 3427 53345
rect 3483 53289 3569 53345
rect 3625 53289 3711 53345
rect 3767 53289 3853 53345
rect 3909 53289 3995 53345
rect 4051 53289 4137 53345
rect 4193 53289 4279 53345
rect 4335 53289 4421 53345
rect 4477 53289 4563 53345
rect 4619 53289 4705 53345
rect 4761 53289 4847 53345
rect 4903 53289 4989 53345
rect 5045 53289 5131 53345
rect 5187 53289 5273 53345
rect 5329 53289 5415 53345
rect 5471 53289 5557 53345
rect 5613 53289 5699 53345
rect 5755 53289 5841 53345
rect 5897 53289 5983 53345
rect 6039 53289 6125 53345
rect 6181 53289 6267 53345
rect 6323 53289 6409 53345
rect 6465 53289 6551 53345
rect 6607 53289 6693 53345
rect 6749 53289 6835 53345
rect 6891 53289 6977 53345
rect 7033 53289 7119 53345
rect 7175 53289 7261 53345
rect 7317 53289 7403 53345
rect 7459 53289 7545 53345
rect 7601 53289 7687 53345
rect 7743 53289 7829 53345
rect 7885 53289 7971 53345
rect 8027 53289 8113 53345
rect 8169 53289 8255 53345
rect 8311 53289 8397 53345
rect 8453 53289 8539 53345
rect 8595 53289 8681 53345
rect 8737 53289 8823 53345
rect 8879 53289 8965 53345
rect 9021 53289 9107 53345
rect 9163 53289 9249 53345
rect 9305 53289 9391 53345
rect 9447 53289 9533 53345
rect 9589 53289 9675 53345
rect 9731 53289 9817 53345
rect 9873 53289 9959 53345
rect 10015 53289 10101 53345
rect 10157 53289 10243 53345
rect 10299 53289 10385 53345
rect 10441 53289 10527 53345
rect 10583 53289 10669 53345
rect 10725 53289 10811 53345
rect 10867 53289 10953 53345
rect 11009 53289 11095 53345
rect 11151 53289 11237 53345
rect 11293 53289 11379 53345
rect 11435 53289 11521 53345
rect 11577 53289 11663 53345
rect 11719 53289 11805 53345
rect 11861 53289 11947 53345
rect 12003 53289 12089 53345
rect 12145 53289 12231 53345
rect 12287 53289 12373 53345
rect 12429 53289 12515 53345
rect 12571 53289 12657 53345
rect 12713 53289 12799 53345
rect 12855 53289 12941 53345
rect 12997 53289 13083 53345
rect 13139 53289 13225 53345
rect 13281 53289 13367 53345
rect 13423 53289 13509 53345
rect 13565 53289 13651 53345
rect 13707 53289 13793 53345
rect 13849 53289 13935 53345
rect 13991 53289 14077 53345
rect 14133 53289 14219 53345
rect 14275 53289 14361 53345
rect 14417 53289 14503 53345
rect 14559 53289 14645 53345
rect 14701 53289 14787 53345
rect 14843 53289 15000 53345
rect 0 53203 15000 53289
rect 0 53147 161 53203
rect 217 53147 303 53203
rect 359 53147 445 53203
rect 501 53147 587 53203
rect 643 53147 729 53203
rect 785 53147 871 53203
rect 927 53147 1013 53203
rect 1069 53147 1155 53203
rect 1211 53147 1297 53203
rect 1353 53147 1439 53203
rect 1495 53147 1581 53203
rect 1637 53147 1723 53203
rect 1779 53147 1865 53203
rect 1921 53147 2007 53203
rect 2063 53147 2149 53203
rect 2205 53147 2291 53203
rect 2347 53147 2433 53203
rect 2489 53147 2575 53203
rect 2631 53147 2717 53203
rect 2773 53147 2859 53203
rect 2915 53147 3001 53203
rect 3057 53147 3143 53203
rect 3199 53147 3285 53203
rect 3341 53147 3427 53203
rect 3483 53147 3569 53203
rect 3625 53147 3711 53203
rect 3767 53147 3853 53203
rect 3909 53147 3995 53203
rect 4051 53147 4137 53203
rect 4193 53147 4279 53203
rect 4335 53147 4421 53203
rect 4477 53147 4563 53203
rect 4619 53147 4705 53203
rect 4761 53147 4847 53203
rect 4903 53147 4989 53203
rect 5045 53147 5131 53203
rect 5187 53147 5273 53203
rect 5329 53147 5415 53203
rect 5471 53147 5557 53203
rect 5613 53147 5699 53203
rect 5755 53147 5841 53203
rect 5897 53147 5983 53203
rect 6039 53147 6125 53203
rect 6181 53147 6267 53203
rect 6323 53147 6409 53203
rect 6465 53147 6551 53203
rect 6607 53147 6693 53203
rect 6749 53147 6835 53203
rect 6891 53147 6977 53203
rect 7033 53147 7119 53203
rect 7175 53147 7261 53203
rect 7317 53147 7403 53203
rect 7459 53147 7545 53203
rect 7601 53147 7687 53203
rect 7743 53147 7829 53203
rect 7885 53147 7971 53203
rect 8027 53147 8113 53203
rect 8169 53147 8255 53203
rect 8311 53147 8397 53203
rect 8453 53147 8539 53203
rect 8595 53147 8681 53203
rect 8737 53147 8823 53203
rect 8879 53147 8965 53203
rect 9021 53147 9107 53203
rect 9163 53147 9249 53203
rect 9305 53147 9391 53203
rect 9447 53147 9533 53203
rect 9589 53147 9675 53203
rect 9731 53147 9817 53203
rect 9873 53147 9959 53203
rect 10015 53147 10101 53203
rect 10157 53147 10243 53203
rect 10299 53147 10385 53203
rect 10441 53147 10527 53203
rect 10583 53147 10669 53203
rect 10725 53147 10811 53203
rect 10867 53147 10953 53203
rect 11009 53147 11095 53203
rect 11151 53147 11237 53203
rect 11293 53147 11379 53203
rect 11435 53147 11521 53203
rect 11577 53147 11663 53203
rect 11719 53147 11805 53203
rect 11861 53147 11947 53203
rect 12003 53147 12089 53203
rect 12145 53147 12231 53203
rect 12287 53147 12373 53203
rect 12429 53147 12515 53203
rect 12571 53147 12657 53203
rect 12713 53147 12799 53203
rect 12855 53147 12941 53203
rect 12997 53147 13083 53203
rect 13139 53147 13225 53203
rect 13281 53147 13367 53203
rect 13423 53147 13509 53203
rect 13565 53147 13651 53203
rect 13707 53147 13793 53203
rect 13849 53147 13935 53203
rect 13991 53147 14077 53203
rect 14133 53147 14219 53203
rect 14275 53147 14361 53203
rect 14417 53147 14503 53203
rect 14559 53147 14645 53203
rect 14701 53147 14787 53203
rect 14843 53147 15000 53203
rect 0 53061 15000 53147
rect 0 53005 161 53061
rect 217 53005 303 53061
rect 359 53005 445 53061
rect 501 53005 587 53061
rect 643 53005 729 53061
rect 785 53005 871 53061
rect 927 53005 1013 53061
rect 1069 53005 1155 53061
rect 1211 53005 1297 53061
rect 1353 53005 1439 53061
rect 1495 53005 1581 53061
rect 1637 53005 1723 53061
rect 1779 53005 1865 53061
rect 1921 53005 2007 53061
rect 2063 53005 2149 53061
rect 2205 53005 2291 53061
rect 2347 53005 2433 53061
rect 2489 53005 2575 53061
rect 2631 53005 2717 53061
rect 2773 53005 2859 53061
rect 2915 53005 3001 53061
rect 3057 53005 3143 53061
rect 3199 53005 3285 53061
rect 3341 53005 3427 53061
rect 3483 53005 3569 53061
rect 3625 53005 3711 53061
rect 3767 53005 3853 53061
rect 3909 53005 3995 53061
rect 4051 53005 4137 53061
rect 4193 53005 4279 53061
rect 4335 53005 4421 53061
rect 4477 53005 4563 53061
rect 4619 53005 4705 53061
rect 4761 53005 4847 53061
rect 4903 53005 4989 53061
rect 5045 53005 5131 53061
rect 5187 53005 5273 53061
rect 5329 53005 5415 53061
rect 5471 53005 5557 53061
rect 5613 53005 5699 53061
rect 5755 53005 5841 53061
rect 5897 53005 5983 53061
rect 6039 53005 6125 53061
rect 6181 53005 6267 53061
rect 6323 53005 6409 53061
rect 6465 53005 6551 53061
rect 6607 53005 6693 53061
rect 6749 53005 6835 53061
rect 6891 53005 6977 53061
rect 7033 53005 7119 53061
rect 7175 53005 7261 53061
rect 7317 53005 7403 53061
rect 7459 53005 7545 53061
rect 7601 53005 7687 53061
rect 7743 53005 7829 53061
rect 7885 53005 7971 53061
rect 8027 53005 8113 53061
rect 8169 53005 8255 53061
rect 8311 53005 8397 53061
rect 8453 53005 8539 53061
rect 8595 53005 8681 53061
rect 8737 53005 8823 53061
rect 8879 53005 8965 53061
rect 9021 53005 9107 53061
rect 9163 53005 9249 53061
rect 9305 53005 9391 53061
rect 9447 53005 9533 53061
rect 9589 53005 9675 53061
rect 9731 53005 9817 53061
rect 9873 53005 9959 53061
rect 10015 53005 10101 53061
rect 10157 53005 10243 53061
rect 10299 53005 10385 53061
rect 10441 53005 10527 53061
rect 10583 53005 10669 53061
rect 10725 53005 10811 53061
rect 10867 53005 10953 53061
rect 11009 53005 11095 53061
rect 11151 53005 11237 53061
rect 11293 53005 11379 53061
rect 11435 53005 11521 53061
rect 11577 53005 11663 53061
rect 11719 53005 11805 53061
rect 11861 53005 11947 53061
rect 12003 53005 12089 53061
rect 12145 53005 12231 53061
rect 12287 53005 12373 53061
rect 12429 53005 12515 53061
rect 12571 53005 12657 53061
rect 12713 53005 12799 53061
rect 12855 53005 12941 53061
rect 12997 53005 13083 53061
rect 13139 53005 13225 53061
rect 13281 53005 13367 53061
rect 13423 53005 13509 53061
rect 13565 53005 13651 53061
rect 13707 53005 13793 53061
rect 13849 53005 13935 53061
rect 13991 53005 14077 53061
rect 14133 53005 14219 53061
rect 14275 53005 14361 53061
rect 14417 53005 14503 53061
rect 14559 53005 14645 53061
rect 14701 53005 14787 53061
rect 14843 53005 15000 53061
rect 0 52919 15000 53005
rect 0 52863 161 52919
rect 217 52863 303 52919
rect 359 52863 445 52919
rect 501 52863 587 52919
rect 643 52863 729 52919
rect 785 52863 871 52919
rect 927 52863 1013 52919
rect 1069 52863 1155 52919
rect 1211 52863 1297 52919
rect 1353 52863 1439 52919
rect 1495 52863 1581 52919
rect 1637 52863 1723 52919
rect 1779 52863 1865 52919
rect 1921 52863 2007 52919
rect 2063 52863 2149 52919
rect 2205 52863 2291 52919
rect 2347 52863 2433 52919
rect 2489 52863 2575 52919
rect 2631 52863 2717 52919
rect 2773 52863 2859 52919
rect 2915 52863 3001 52919
rect 3057 52863 3143 52919
rect 3199 52863 3285 52919
rect 3341 52863 3427 52919
rect 3483 52863 3569 52919
rect 3625 52863 3711 52919
rect 3767 52863 3853 52919
rect 3909 52863 3995 52919
rect 4051 52863 4137 52919
rect 4193 52863 4279 52919
rect 4335 52863 4421 52919
rect 4477 52863 4563 52919
rect 4619 52863 4705 52919
rect 4761 52863 4847 52919
rect 4903 52863 4989 52919
rect 5045 52863 5131 52919
rect 5187 52863 5273 52919
rect 5329 52863 5415 52919
rect 5471 52863 5557 52919
rect 5613 52863 5699 52919
rect 5755 52863 5841 52919
rect 5897 52863 5983 52919
rect 6039 52863 6125 52919
rect 6181 52863 6267 52919
rect 6323 52863 6409 52919
rect 6465 52863 6551 52919
rect 6607 52863 6693 52919
rect 6749 52863 6835 52919
rect 6891 52863 6977 52919
rect 7033 52863 7119 52919
rect 7175 52863 7261 52919
rect 7317 52863 7403 52919
rect 7459 52863 7545 52919
rect 7601 52863 7687 52919
rect 7743 52863 7829 52919
rect 7885 52863 7971 52919
rect 8027 52863 8113 52919
rect 8169 52863 8255 52919
rect 8311 52863 8397 52919
rect 8453 52863 8539 52919
rect 8595 52863 8681 52919
rect 8737 52863 8823 52919
rect 8879 52863 8965 52919
rect 9021 52863 9107 52919
rect 9163 52863 9249 52919
rect 9305 52863 9391 52919
rect 9447 52863 9533 52919
rect 9589 52863 9675 52919
rect 9731 52863 9817 52919
rect 9873 52863 9959 52919
rect 10015 52863 10101 52919
rect 10157 52863 10243 52919
rect 10299 52863 10385 52919
rect 10441 52863 10527 52919
rect 10583 52863 10669 52919
rect 10725 52863 10811 52919
rect 10867 52863 10953 52919
rect 11009 52863 11095 52919
rect 11151 52863 11237 52919
rect 11293 52863 11379 52919
rect 11435 52863 11521 52919
rect 11577 52863 11663 52919
rect 11719 52863 11805 52919
rect 11861 52863 11947 52919
rect 12003 52863 12089 52919
rect 12145 52863 12231 52919
rect 12287 52863 12373 52919
rect 12429 52863 12515 52919
rect 12571 52863 12657 52919
rect 12713 52863 12799 52919
rect 12855 52863 12941 52919
rect 12997 52863 13083 52919
rect 13139 52863 13225 52919
rect 13281 52863 13367 52919
rect 13423 52863 13509 52919
rect 13565 52863 13651 52919
rect 13707 52863 13793 52919
rect 13849 52863 13935 52919
rect 13991 52863 14077 52919
rect 14133 52863 14219 52919
rect 14275 52863 14361 52919
rect 14417 52863 14503 52919
rect 14559 52863 14645 52919
rect 14701 52863 14787 52919
rect 14843 52863 15000 52919
rect 0 52777 15000 52863
rect 0 52721 161 52777
rect 217 52721 303 52777
rect 359 52721 445 52777
rect 501 52721 587 52777
rect 643 52721 729 52777
rect 785 52721 871 52777
rect 927 52721 1013 52777
rect 1069 52721 1155 52777
rect 1211 52721 1297 52777
rect 1353 52721 1439 52777
rect 1495 52721 1581 52777
rect 1637 52721 1723 52777
rect 1779 52721 1865 52777
rect 1921 52721 2007 52777
rect 2063 52721 2149 52777
rect 2205 52721 2291 52777
rect 2347 52721 2433 52777
rect 2489 52721 2575 52777
rect 2631 52721 2717 52777
rect 2773 52721 2859 52777
rect 2915 52721 3001 52777
rect 3057 52721 3143 52777
rect 3199 52721 3285 52777
rect 3341 52721 3427 52777
rect 3483 52721 3569 52777
rect 3625 52721 3711 52777
rect 3767 52721 3853 52777
rect 3909 52721 3995 52777
rect 4051 52721 4137 52777
rect 4193 52721 4279 52777
rect 4335 52721 4421 52777
rect 4477 52721 4563 52777
rect 4619 52721 4705 52777
rect 4761 52721 4847 52777
rect 4903 52721 4989 52777
rect 5045 52721 5131 52777
rect 5187 52721 5273 52777
rect 5329 52721 5415 52777
rect 5471 52721 5557 52777
rect 5613 52721 5699 52777
rect 5755 52721 5841 52777
rect 5897 52721 5983 52777
rect 6039 52721 6125 52777
rect 6181 52721 6267 52777
rect 6323 52721 6409 52777
rect 6465 52721 6551 52777
rect 6607 52721 6693 52777
rect 6749 52721 6835 52777
rect 6891 52721 6977 52777
rect 7033 52721 7119 52777
rect 7175 52721 7261 52777
rect 7317 52721 7403 52777
rect 7459 52721 7545 52777
rect 7601 52721 7687 52777
rect 7743 52721 7829 52777
rect 7885 52721 7971 52777
rect 8027 52721 8113 52777
rect 8169 52721 8255 52777
rect 8311 52721 8397 52777
rect 8453 52721 8539 52777
rect 8595 52721 8681 52777
rect 8737 52721 8823 52777
rect 8879 52721 8965 52777
rect 9021 52721 9107 52777
rect 9163 52721 9249 52777
rect 9305 52721 9391 52777
rect 9447 52721 9533 52777
rect 9589 52721 9675 52777
rect 9731 52721 9817 52777
rect 9873 52721 9959 52777
rect 10015 52721 10101 52777
rect 10157 52721 10243 52777
rect 10299 52721 10385 52777
rect 10441 52721 10527 52777
rect 10583 52721 10669 52777
rect 10725 52721 10811 52777
rect 10867 52721 10953 52777
rect 11009 52721 11095 52777
rect 11151 52721 11237 52777
rect 11293 52721 11379 52777
rect 11435 52721 11521 52777
rect 11577 52721 11663 52777
rect 11719 52721 11805 52777
rect 11861 52721 11947 52777
rect 12003 52721 12089 52777
rect 12145 52721 12231 52777
rect 12287 52721 12373 52777
rect 12429 52721 12515 52777
rect 12571 52721 12657 52777
rect 12713 52721 12799 52777
rect 12855 52721 12941 52777
rect 12997 52721 13083 52777
rect 13139 52721 13225 52777
rect 13281 52721 13367 52777
rect 13423 52721 13509 52777
rect 13565 52721 13651 52777
rect 13707 52721 13793 52777
rect 13849 52721 13935 52777
rect 13991 52721 14077 52777
rect 14133 52721 14219 52777
rect 14275 52721 14361 52777
rect 14417 52721 14503 52777
rect 14559 52721 14645 52777
rect 14701 52721 14787 52777
rect 14843 52721 15000 52777
rect 0 52635 15000 52721
rect 0 52579 161 52635
rect 217 52579 303 52635
rect 359 52579 445 52635
rect 501 52579 587 52635
rect 643 52579 729 52635
rect 785 52579 871 52635
rect 927 52579 1013 52635
rect 1069 52579 1155 52635
rect 1211 52579 1297 52635
rect 1353 52579 1439 52635
rect 1495 52579 1581 52635
rect 1637 52579 1723 52635
rect 1779 52579 1865 52635
rect 1921 52579 2007 52635
rect 2063 52579 2149 52635
rect 2205 52579 2291 52635
rect 2347 52579 2433 52635
rect 2489 52579 2575 52635
rect 2631 52579 2717 52635
rect 2773 52579 2859 52635
rect 2915 52579 3001 52635
rect 3057 52579 3143 52635
rect 3199 52579 3285 52635
rect 3341 52579 3427 52635
rect 3483 52579 3569 52635
rect 3625 52579 3711 52635
rect 3767 52579 3853 52635
rect 3909 52579 3995 52635
rect 4051 52579 4137 52635
rect 4193 52579 4279 52635
rect 4335 52579 4421 52635
rect 4477 52579 4563 52635
rect 4619 52579 4705 52635
rect 4761 52579 4847 52635
rect 4903 52579 4989 52635
rect 5045 52579 5131 52635
rect 5187 52579 5273 52635
rect 5329 52579 5415 52635
rect 5471 52579 5557 52635
rect 5613 52579 5699 52635
rect 5755 52579 5841 52635
rect 5897 52579 5983 52635
rect 6039 52579 6125 52635
rect 6181 52579 6267 52635
rect 6323 52579 6409 52635
rect 6465 52579 6551 52635
rect 6607 52579 6693 52635
rect 6749 52579 6835 52635
rect 6891 52579 6977 52635
rect 7033 52579 7119 52635
rect 7175 52579 7261 52635
rect 7317 52579 7403 52635
rect 7459 52579 7545 52635
rect 7601 52579 7687 52635
rect 7743 52579 7829 52635
rect 7885 52579 7971 52635
rect 8027 52579 8113 52635
rect 8169 52579 8255 52635
rect 8311 52579 8397 52635
rect 8453 52579 8539 52635
rect 8595 52579 8681 52635
rect 8737 52579 8823 52635
rect 8879 52579 8965 52635
rect 9021 52579 9107 52635
rect 9163 52579 9249 52635
rect 9305 52579 9391 52635
rect 9447 52579 9533 52635
rect 9589 52579 9675 52635
rect 9731 52579 9817 52635
rect 9873 52579 9959 52635
rect 10015 52579 10101 52635
rect 10157 52579 10243 52635
rect 10299 52579 10385 52635
rect 10441 52579 10527 52635
rect 10583 52579 10669 52635
rect 10725 52579 10811 52635
rect 10867 52579 10953 52635
rect 11009 52579 11095 52635
rect 11151 52579 11237 52635
rect 11293 52579 11379 52635
rect 11435 52579 11521 52635
rect 11577 52579 11663 52635
rect 11719 52579 11805 52635
rect 11861 52579 11947 52635
rect 12003 52579 12089 52635
rect 12145 52579 12231 52635
rect 12287 52579 12373 52635
rect 12429 52579 12515 52635
rect 12571 52579 12657 52635
rect 12713 52579 12799 52635
rect 12855 52579 12941 52635
rect 12997 52579 13083 52635
rect 13139 52579 13225 52635
rect 13281 52579 13367 52635
rect 13423 52579 13509 52635
rect 13565 52579 13651 52635
rect 13707 52579 13793 52635
rect 13849 52579 13935 52635
rect 13991 52579 14077 52635
rect 14133 52579 14219 52635
rect 14275 52579 14361 52635
rect 14417 52579 14503 52635
rect 14559 52579 14645 52635
rect 14701 52579 14787 52635
rect 14843 52579 15000 52635
rect 0 52493 15000 52579
rect 0 52437 161 52493
rect 217 52437 303 52493
rect 359 52437 445 52493
rect 501 52437 587 52493
rect 643 52437 729 52493
rect 785 52437 871 52493
rect 927 52437 1013 52493
rect 1069 52437 1155 52493
rect 1211 52437 1297 52493
rect 1353 52437 1439 52493
rect 1495 52437 1581 52493
rect 1637 52437 1723 52493
rect 1779 52437 1865 52493
rect 1921 52437 2007 52493
rect 2063 52437 2149 52493
rect 2205 52437 2291 52493
rect 2347 52437 2433 52493
rect 2489 52437 2575 52493
rect 2631 52437 2717 52493
rect 2773 52437 2859 52493
rect 2915 52437 3001 52493
rect 3057 52437 3143 52493
rect 3199 52437 3285 52493
rect 3341 52437 3427 52493
rect 3483 52437 3569 52493
rect 3625 52437 3711 52493
rect 3767 52437 3853 52493
rect 3909 52437 3995 52493
rect 4051 52437 4137 52493
rect 4193 52437 4279 52493
rect 4335 52437 4421 52493
rect 4477 52437 4563 52493
rect 4619 52437 4705 52493
rect 4761 52437 4847 52493
rect 4903 52437 4989 52493
rect 5045 52437 5131 52493
rect 5187 52437 5273 52493
rect 5329 52437 5415 52493
rect 5471 52437 5557 52493
rect 5613 52437 5699 52493
rect 5755 52437 5841 52493
rect 5897 52437 5983 52493
rect 6039 52437 6125 52493
rect 6181 52437 6267 52493
rect 6323 52437 6409 52493
rect 6465 52437 6551 52493
rect 6607 52437 6693 52493
rect 6749 52437 6835 52493
rect 6891 52437 6977 52493
rect 7033 52437 7119 52493
rect 7175 52437 7261 52493
rect 7317 52437 7403 52493
rect 7459 52437 7545 52493
rect 7601 52437 7687 52493
rect 7743 52437 7829 52493
rect 7885 52437 7971 52493
rect 8027 52437 8113 52493
rect 8169 52437 8255 52493
rect 8311 52437 8397 52493
rect 8453 52437 8539 52493
rect 8595 52437 8681 52493
rect 8737 52437 8823 52493
rect 8879 52437 8965 52493
rect 9021 52437 9107 52493
rect 9163 52437 9249 52493
rect 9305 52437 9391 52493
rect 9447 52437 9533 52493
rect 9589 52437 9675 52493
rect 9731 52437 9817 52493
rect 9873 52437 9959 52493
rect 10015 52437 10101 52493
rect 10157 52437 10243 52493
rect 10299 52437 10385 52493
rect 10441 52437 10527 52493
rect 10583 52437 10669 52493
rect 10725 52437 10811 52493
rect 10867 52437 10953 52493
rect 11009 52437 11095 52493
rect 11151 52437 11237 52493
rect 11293 52437 11379 52493
rect 11435 52437 11521 52493
rect 11577 52437 11663 52493
rect 11719 52437 11805 52493
rect 11861 52437 11947 52493
rect 12003 52437 12089 52493
rect 12145 52437 12231 52493
rect 12287 52437 12373 52493
rect 12429 52437 12515 52493
rect 12571 52437 12657 52493
rect 12713 52437 12799 52493
rect 12855 52437 12941 52493
rect 12997 52437 13083 52493
rect 13139 52437 13225 52493
rect 13281 52437 13367 52493
rect 13423 52437 13509 52493
rect 13565 52437 13651 52493
rect 13707 52437 13793 52493
rect 13849 52437 13935 52493
rect 13991 52437 14077 52493
rect 14133 52437 14219 52493
rect 14275 52437 14361 52493
rect 14417 52437 14503 52493
rect 14559 52437 14645 52493
rect 14701 52437 14787 52493
rect 14843 52437 15000 52493
rect 0 52400 15000 52437
rect 0 52163 15000 52200
rect 0 52107 161 52163
rect 217 52107 303 52163
rect 359 52107 445 52163
rect 501 52107 587 52163
rect 643 52107 729 52163
rect 785 52107 871 52163
rect 927 52107 1013 52163
rect 1069 52107 1155 52163
rect 1211 52107 1297 52163
rect 1353 52107 1439 52163
rect 1495 52107 1581 52163
rect 1637 52107 1723 52163
rect 1779 52107 1865 52163
rect 1921 52107 2007 52163
rect 2063 52107 2149 52163
rect 2205 52107 2291 52163
rect 2347 52107 2433 52163
rect 2489 52107 2575 52163
rect 2631 52107 2717 52163
rect 2773 52107 2859 52163
rect 2915 52107 3001 52163
rect 3057 52107 3143 52163
rect 3199 52107 3285 52163
rect 3341 52107 3427 52163
rect 3483 52107 3569 52163
rect 3625 52107 3711 52163
rect 3767 52107 3853 52163
rect 3909 52107 3995 52163
rect 4051 52107 4137 52163
rect 4193 52107 4279 52163
rect 4335 52107 4421 52163
rect 4477 52107 4563 52163
rect 4619 52107 4705 52163
rect 4761 52107 4847 52163
rect 4903 52107 4989 52163
rect 5045 52107 5131 52163
rect 5187 52107 5273 52163
rect 5329 52107 5415 52163
rect 5471 52107 5557 52163
rect 5613 52107 5699 52163
rect 5755 52107 5841 52163
rect 5897 52107 5983 52163
rect 6039 52107 6125 52163
rect 6181 52107 6267 52163
rect 6323 52107 6409 52163
rect 6465 52107 6551 52163
rect 6607 52107 6693 52163
rect 6749 52107 6835 52163
rect 6891 52107 6977 52163
rect 7033 52107 7119 52163
rect 7175 52107 7261 52163
rect 7317 52107 7403 52163
rect 7459 52107 7545 52163
rect 7601 52107 7687 52163
rect 7743 52107 7829 52163
rect 7885 52107 7971 52163
rect 8027 52107 8113 52163
rect 8169 52107 8255 52163
rect 8311 52107 8397 52163
rect 8453 52107 8539 52163
rect 8595 52107 8681 52163
rect 8737 52107 8823 52163
rect 8879 52107 8965 52163
rect 9021 52107 9107 52163
rect 9163 52107 9249 52163
rect 9305 52107 9391 52163
rect 9447 52107 9533 52163
rect 9589 52107 9675 52163
rect 9731 52107 9817 52163
rect 9873 52107 9959 52163
rect 10015 52107 10101 52163
rect 10157 52107 10243 52163
rect 10299 52107 10385 52163
rect 10441 52107 10527 52163
rect 10583 52107 10669 52163
rect 10725 52107 10811 52163
rect 10867 52107 10953 52163
rect 11009 52107 11095 52163
rect 11151 52107 11237 52163
rect 11293 52107 11379 52163
rect 11435 52107 11521 52163
rect 11577 52107 11663 52163
rect 11719 52107 11805 52163
rect 11861 52107 11947 52163
rect 12003 52107 12089 52163
rect 12145 52107 12231 52163
rect 12287 52107 12373 52163
rect 12429 52107 12515 52163
rect 12571 52107 12657 52163
rect 12713 52107 12799 52163
rect 12855 52107 12941 52163
rect 12997 52107 13083 52163
rect 13139 52107 13225 52163
rect 13281 52107 13367 52163
rect 13423 52107 13509 52163
rect 13565 52107 13651 52163
rect 13707 52107 13793 52163
rect 13849 52107 13935 52163
rect 13991 52107 14077 52163
rect 14133 52107 14219 52163
rect 14275 52107 14361 52163
rect 14417 52107 14503 52163
rect 14559 52107 14645 52163
rect 14701 52107 14787 52163
rect 14843 52107 15000 52163
rect 0 52021 15000 52107
rect 0 51965 161 52021
rect 217 51965 303 52021
rect 359 51965 445 52021
rect 501 51965 587 52021
rect 643 51965 729 52021
rect 785 51965 871 52021
rect 927 51965 1013 52021
rect 1069 51965 1155 52021
rect 1211 51965 1297 52021
rect 1353 51965 1439 52021
rect 1495 51965 1581 52021
rect 1637 51965 1723 52021
rect 1779 51965 1865 52021
rect 1921 51965 2007 52021
rect 2063 51965 2149 52021
rect 2205 51965 2291 52021
rect 2347 51965 2433 52021
rect 2489 51965 2575 52021
rect 2631 51965 2717 52021
rect 2773 51965 2859 52021
rect 2915 51965 3001 52021
rect 3057 51965 3143 52021
rect 3199 51965 3285 52021
rect 3341 51965 3427 52021
rect 3483 51965 3569 52021
rect 3625 51965 3711 52021
rect 3767 51965 3853 52021
rect 3909 51965 3995 52021
rect 4051 51965 4137 52021
rect 4193 51965 4279 52021
rect 4335 51965 4421 52021
rect 4477 51965 4563 52021
rect 4619 51965 4705 52021
rect 4761 51965 4847 52021
rect 4903 51965 4989 52021
rect 5045 51965 5131 52021
rect 5187 51965 5273 52021
rect 5329 51965 5415 52021
rect 5471 51965 5557 52021
rect 5613 51965 5699 52021
rect 5755 51965 5841 52021
rect 5897 51965 5983 52021
rect 6039 51965 6125 52021
rect 6181 51965 6267 52021
rect 6323 51965 6409 52021
rect 6465 51965 6551 52021
rect 6607 51965 6693 52021
rect 6749 51965 6835 52021
rect 6891 51965 6977 52021
rect 7033 51965 7119 52021
rect 7175 51965 7261 52021
rect 7317 51965 7403 52021
rect 7459 51965 7545 52021
rect 7601 51965 7687 52021
rect 7743 51965 7829 52021
rect 7885 51965 7971 52021
rect 8027 51965 8113 52021
rect 8169 51965 8255 52021
rect 8311 51965 8397 52021
rect 8453 51965 8539 52021
rect 8595 51965 8681 52021
rect 8737 51965 8823 52021
rect 8879 51965 8965 52021
rect 9021 51965 9107 52021
rect 9163 51965 9249 52021
rect 9305 51965 9391 52021
rect 9447 51965 9533 52021
rect 9589 51965 9675 52021
rect 9731 51965 9817 52021
rect 9873 51965 9959 52021
rect 10015 51965 10101 52021
rect 10157 51965 10243 52021
rect 10299 51965 10385 52021
rect 10441 51965 10527 52021
rect 10583 51965 10669 52021
rect 10725 51965 10811 52021
rect 10867 51965 10953 52021
rect 11009 51965 11095 52021
rect 11151 51965 11237 52021
rect 11293 51965 11379 52021
rect 11435 51965 11521 52021
rect 11577 51965 11663 52021
rect 11719 51965 11805 52021
rect 11861 51965 11947 52021
rect 12003 51965 12089 52021
rect 12145 51965 12231 52021
rect 12287 51965 12373 52021
rect 12429 51965 12515 52021
rect 12571 51965 12657 52021
rect 12713 51965 12799 52021
rect 12855 51965 12941 52021
rect 12997 51965 13083 52021
rect 13139 51965 13225 52021
rect 13281 51965 13367 52021
rect 13423 51965 13509 52021
rect 13565 51965 13651 52021
rect 13707 51965 13793 52021
rect 13849 51965 13935 52021
rect 13991 51965 14077 52021
rect 14133 51965 14219 52021
rect 14275 51965 14361 52021
rect 14417 51965 14503 52021
rect 14559 51965 14645 52021
rect 14701 51965 14787 52021
rect 14843 51965 15000 52021
rect 0 51879 15000 51965
rect 0 51823 161 51879
rect 217 51823 303 51879
rect 359 51823 445 51879
rect 501 51823 587 51879
rect 643 51823 729 51879
rect 785 51823 871 51879
rect 927 51823 1013 51879
rect 1069 51823 1155 51879
rect 1211 51823 1297 51879
rect 1353 51823 1439 51879
rect 1495 51823 1581 51879
rect 1637 51823 1723 51879
rect 1779 51823 1865 51879
rect 1921 51823 2007 51879
rect 2063 51823 2149 51879
rect 2205 51823 2291 51879
rect 2347 51823 2433 51879
rect 2489 51823 2575 51879
rect 2631 51823 2717 51879
rect 2773 51823 2859 51879
rect 2915 51823 3001 51879
rect 3057 51823 3143 51879
rect 3199 51823 3285 51879
rect 3341 51823 3427 51879
rect 3483 51823 3569 51879
rect 3625 51823 3711 51879
rect 3767 51823 3853 51879
rect 3909 51823 3995 51879
rect 4051 51823 4137 51879
rect 4193 51823 4279 51879
rect 4335 51823 4421 51879
rect 4477 51823 4563 51879
rect 4619 51823 4705 51879
rect 4761 51823 4847 51879
rect 4903 51823 4989 51879
rect 5045 51823 5131 51879
rect 5187 51823 5273 51879
rect 5329 51823 5415 51879
rect 5471 51823 5557 51879
rect 5613 51823 5699 51879
rect 5755 51823 5841 51879
rect 5897 51823 5983 51879
rect 6039 51823 6125 51879
rect 6181 51823 6267 51879
rect 6323 51823 6409 51879
rect 6465 51823 6551 51879
rect 6607 51823 6693 51879
rect 6749 51823 6835 51879
rect 6891 51823 6977 51879
rect 7033 51823 7119 51879
rect 7175 51823 7261 51879
rect 7317 51823 7403 51879
rect 7459 51823 7545 51879
rect 7601 51823 7687 51879
rect 7743 51823 7829 51879
rect 7885 51823 7971 51879
rect 8027 51823 8113 51879
rect 8169 51823 8255 51879
rect 8311 51823 8397 51879
rect 8453 51823 8539 51879
rect 8595 51823 8681 51879
rect 8737 51823 8823 51879
rect 8879 51823 8965 51879
rect 9021 51823 9107 51879
rect 9163 51823 9249 51879
rect 9305 51823 9391 51879
rect 9447 51823 9533 51879
rect 9589 51823 9675 51879
rect 9731 51823 9817 51879
rect 9873 51823 9959 51879
rect 10015 51823 10101 51879
rect 10157 51823 10243 51879
rect 10299 51823 10385 51879
rect 10441 51823 10527 51879
rect 10583 51823 10669 51879
rect 10725 51823 10811 51879
rect 10867 51823 10953 51879
rect 11009 51823 11095 51879
rect 11151 51823 11237 51879
rect 11293 51823 11379 51879
rect 11435 51823 11521 51879
rect 11577 51823 11663 51879
rect 11719 51823 11805 51879
rect 11861 51823 11947 51879
rect 12003 51823 12089 51879
rect 12145 51823 12231 51879
rect 12287 51823 12373 51879
rect 12429 51823 12515 51879
rect 12571 51823 12657 51879
rect 12713 51823 12799 51879
rect 12855 51823 12941 51879
rect 12997 51823 13083 51879
rect 13139 51823 13225 51879
rect 13281 51823 13367 51879
rect 13423 51823 13509 51879
rect 13565 51823 13651 51879
rect 13707 51823 13793 51879
rect 13849 51823 13935 51879
rect 13991 51823 14077 51879
rect 14133 51823 14219 51879
rect 14275 51823 14361 51879
rect 14417 51823 14503 51879
rect 14559 51823 14645 51879
rect 14701 51823 14787 51879
rect 14843 51823 15000 51879
rect 0 51737 15000 51823
rect 0 51681 161 51737
rect 217 51681 303 51737
rect 359 51681 445 51737
rect 501 51681 587 51737
rect 643 51681 729 51737
rect 785 51681 871 51737
rect 927 51681 1013 51737
rect 1069 51681 1155 51737
rect 1211 51681 1297 51737
rect 1353 51681 1439 51737
rect 1495 51681 1581 51737
rect 1637 51681 1723 51737
rect 1779 51681 1865 51737
rect 1921 51681 2007 51737
rect 2063 51681 2149 51737
rect 2205 51681 2291 51737
rect 2347 51681 2433 51737
rect 2489 51681 2575 51737
rect 2631 51681 2717 51737
rect 2773 51681 2859 51737
rect 2915 51681 3001 51737
rect 3057 51681 3143 51737
rect 3199 51681 3285 51737
rect 3341 51681 3427 51737
rect 3483 51681 3569 51737
rect 3625 51681 3711 51737
rect 3767 51681 3853 51737
rect 3909 51681 3995 51737
rect 4051 51681 4137 51737
rect 4193 51681 4279 51737
rect 4335 51681 4421 51737
rect 4477 51681 4563 51737
rect 4619 51681 4705 51737
rect 4761 51681 4847 51737
rect 4903 51681 4989 51737
rect 5045 51681 5131 51737
rect 5187 51681 5273 51737
rect 5329 51681 5415 51737
rect 5471 51681 5557 51737
rect 5613 51681 5699 51737
rect 5755 51681 5841 51737
rect 5897 51681 5983 51737
rect 6039 51681 6125 51737
rect 6181 51681 6267 51737
rect 6323 51681 6409 51737
rect 6465 51681 6551 51737
rect 6607 51681 6693 51737
rect 6749 51681 6835 51737
rect 6891 51681 6977 51737
rect 7033 51681 7119 51737
rect 7175 51681 7261 51737
rect 7317 51681 7403 51737
rect 7459 51681 7545 51737
rect 7601 51681 7687 51737
rect 7743 51681 7829 51737
rect 7885 51681 7971 51737
rect 8027 51681 8113 51737
rect 8169 51681 8255 51737
rect 8311 51681 8397 51737
rect 8453 51681 8539 51737
rect 8595 51681 8681 51737
rect 8737 51681 8823 51737
rect 8879 51681 8965 51737
rect 9021 51681 9107 51737
rect 9163 51681 9249 51737
rect 9305 51681 9391 51737
rect 9447 51681 9533 51737
rect 9589 51681 9675 51737
rect 9731 51681 9817 51737
rect 9873 51681 9959 51737
rect 10015 51681 10101 51737
rect 10157 51681 10243 51737
rect 10299 51681 10385 51737
rect 10441 51681 10527 51737
rect 10583 51681 10669 51737
rect 10725 51681 10811 51737
rect 10867 51681 10953 51737
rect 11009 51681 11095 51737
rect 11151 51681 11237 51737
rect 11293 51681 11379 51737
rect 11435 51681 11521 51737
rect 11577 51681 11663 51737
rect 11719 51681 11805 51737
rect 11861 51681 11947 51737
rect 12003 51681 12089 51737
rect 12145 51681 12231 51737
rect 12287 51681 12373 51737
rect 12429 51681 12515 51737
rect 12571 51681 12657 51737
rect 12713 51681 12799 51737
rect 12855 51681 12941 51737
rect 12997 51681 13083 51737
rect 13139 51681 13225 51737
rect 13281 51681 13367 51737
rect 13423 51681 13509 51737
rect 13565 51681 13651 51737
rect 13707 51681 13793 51737
rect 13849 51681 13935 51737
rect 13991 51681 14077 51737
rect 14133 51681 14219 51737
rect 14275 51681 14361 51737
rect 14417 51681 14503 51737
rect 14559 51681 14645 51737
rect 14701 51681 14787 51737
rect 14843 51681 15000 51737
rect 0 51595 15000 51681
rect 0 51539 161 51595
rect 217 51539 303 51595
rect 359 51539 445 51595
rect 501 51539 587 51595
rect 643 51539 729 51595
rect 785 51539 871 51595
rect 927 51539 1013 51595
rect 1069 51539 1155 51595
rect 1211 51539 1297 51595
rect 1353 51539 1439 51595
rect 1495 51539 1581 51595
rect 1637 51539 1723 51595
rect 1779 51539 1865 51595
rect 1921 51539 2007 51595
rect 2063 51539 2149 51595
rect 2205 51539 2291 51595
rect 2347 51539 2433 51595
rect 2489 51539 2575 51595
rect 2631 51539 2717 51595
rect 2773 51539 2859 51595
rect 2915 51539 3001 51595
rect 3057 51539 3143 51595
rect 3199 51539 3285 51595
rect 3341 51539 3427 51595
rect 3483 51539 3569 51595
rect 3625 51539 3711 51595
rect 3767 51539 3853 51595
rect 3909 51539 3995 51595
rect 4051 51539 4137 51595
rect 4193 51539 4279 51595
rect 4335 51539 4421 51595
rect 4477 51539 4563 51595
rect 4619 51539 4705 51595
rect 4761 51539 4847 51595
rect 4903 51539 4989 51595
rect 5045 51539 5131 51595
rect 5187 51539 5273 51595
rect 5329 51539 5415 51595
rect 5471 51539 5557 51595
rect 5613 51539 5699 51595
rect 5755 51539 5841 51595
rect 5897 51539 5983 51595
rect 6039 51539 6125 51595
rect 6181 51539 6267 51595
rect 6323 51539 6409 51595
rect 6465 51539 6551 51595
rect 6607 51539 6693 51595
rect 6749 51539 6835 51595
rect 6891 51539 6977 51595
rect 7033 51539 7119 51595
rect 7175 51539 7261 51595
rect 7317 51539 7403 51595
rect 7459 51539 7545 51595
rect 7601 51539 7687 51595
rect 7743 51539 7829 51595
rect 7885 51539 7971 51595
rect 8027 51539 8113 51595
rect 8169 51539 8255 51595
rect 8311 51539 8397 51595
rect 8453 51539 8539 51595
rect 8595 51539 8681 51595
rect 8737 51539 8823 51595
rect 8879 51539 8965 51595
rect 9021 51539 9107 51595
rect 9163 51539 9249 51595
rect 9305 51539 9391 51595
rect 9447 51539 9533 51595
rect 9589 51539 9675 51595
rect 9731 51539 9817 51595
rect 9873 51539 9959 51595
rect 10015 51539 10101 51595
rect 10157 51539 10243 51595
rect 10299 51539 10385 51595
rect 10441 51539 10527 51595
rect 10583 51539 10669 51595
rect 10725 51539 10811 51595
rect 10867 51539 10953 51595
rect 11009 51539 11095 51595
rect 11151 51539 11237 51595
rect 11293 51539 11379 51595
rect 11435 51539 11521 51595
rect 11577 51539 11663 51595
rect 11719 51539 11805 51595
rect 11861 51539 11947 51595
rect 12003 51539 12089 51595
rect 12145 51539 12231 51595
rect 12287 51539 12373 51595
rect 12429 51539 12515 51595
rect 12571 51539 12657 51595
rect 12713 51539 12799 51595
rect 12855 51539 12941 51595
rect 12997 51539 13083 51595
rect 13139 51539 13225 51595
rect 13281 51539 13367 51595
rect 13423 51539 13509 51595
rect 13565 51539 13651 51595
rect 13707 51539 13793 51595
rect 13849 51539 13935 51595
rect 13991 51539 14077 51595
rect 14133 51539 14219 51595
rect 14275 51539 14361 51595
rect 14417 51539 14503 51595
rect 14559 51539 14645 51595
rect 14701 51539 14787 51595
rect 14843 51539 15000 51595
rect 0 51453 15000 51539
rect 0 51397 161 51453
rect 217 51397 303 51453
rect 359 51397 445 51453
rect 501 51397 587 51453
rect 643 51397 729 51453
rect 785 51397 871 51453
rect 927 51397 1013 51453
rect 1069 51397 1155 51453
rect 1211 51397 1297 51453
rect 1353 51397 1439 51453
rect 1495 51397 1581 51453
rect 1637 51397 1723 51453
rect 1779 51397 1865 51453
rect 1921 51397 2007 51453
rect 2063 51397 2149 51453
rect 2205 51397 2291 51453
rect 2347 51397 2433 51453
rect 2489 51397 2575 51453
rect 2631 51397 2717 51453
rect 2773 51397 2859 51453
rect 2915 51397 3001 51453
rect 3057 51397 3143 51453
rect 3199 51397 3285 51453
rect 3341 51397 3427 51453
rect 3483 51397 3569 51453
rect 3625 51397 3711 51453
rect 3767 51397 3853 51453
rect 3909 51397 3995 51453
rect 4051 51397 4137 51453
rect 4193 51397 4279 51453
rect 4335 51397 4421 51453
rect 4477 51397 4563 51453
rect 4619 51397 4705 51453
rect 4761 51397 4847 51453
rect 4903 51397 4989 51453
rect 5045 51397 5131 51453
rect 5187 51397 5273 51453
rect 5329 51397 5415 51453
rect 5471 51397 5557 51453
rect 5613 51397 5699 51453
rect 5755 51397 5841 51453
rect 5897 51397 5983 51453
rect 6039 51397 6125 51453
rect 6181 51397 6267 51453
rect 6323 51397 6409 51453
rect 6465 51397 6551 51453
rect 6607 51397 6693 51453
rect 6749 51397 6835 51453
rect 6891 51397 6977 51453
rect 7033 51397 7119 51453
rect 7175 51397 7261 51453
rect 7317 51397 7403 51453
rect 7459 51397 7545 51453
rect 7601 51397 7687 51453
rect 7743 51397 7829 51453
rect 7885 51397 7971 51453
rect 8027 51397 8113 51453
rect 8169 51397 8255 51453
rect 8311 51397 8397 51453
rect 8453 51397 8539 51453
rect 8595 51397 8681 51453
rect 8737 51397 8823 51453
rect 8879 51397 8965 51453
rect 9021 51397 9107 51453
rect 9163 51397 9249 51453
rect 9305 51397 9391 51453
rect 9447 51397 9533 51453
rect 9589 51397 9675 51453
rect 9731 51397 9817 51453
rect 9873 51397 9959 51453
rect 10015 51397 10101 51453
rect 10157 51397 10243 51453
rect 10299 51397 10385 51453
rect 10441 51397 10527 51453
rect 10583 51397 10669 51453
rect 10725 51397 10811 51453
rect 10867 51397 10953 51453
rect 11009 51397 11095 51453
rect 11151 51397 11237 51453
rect 11293 51397 11379 51453
rect 11435 51397 11521 51453
rect 11577 51397 11663 51453
rect 11719 51397 11805 51453
rect 11861 51397 11947 51453
rect 12003 51397 12089 51453
rect 12145 51397 12231 51453
rect 12287 51397 12373 51453
rect 12429 51397 12515 51453
rect 12571 51397 12657 51453
rect 12713 51397 12799 51453
rect 12855 51397 12941 51453
rect 12997 51397 13083 51453
rect 13139 51397 13225 51453
rect 13281 51397 13367 51453
rect 13423 51397 13509 51453
rect 13565 51397 13651 51453
rect 13707 51397 13793 51453
rect 13849 51397 13935 51453
rect 13991 51397 14077 51453
rect 14133 51397 14219 51453
rect 14275 51397 14361 51453
rect 14417 51397 14503 51453
rect 14559 51397 14645 51453
rect 14701 51397 14787 51453
rect 14843 51397 15000 51453
rect 0 51311 15000 51397
rect 0 51255 161 51311
rect 217 51255 303 51311
rect 359 51255 445 51311
rect 501 51255 587 51311
rect 643 51255 729 51311
rect 785 51255 871 51311
rect 927 51255 1013 51311
rect 1069 51255 1155 51311
rect 1211 51255 1297 51311
rect 1353 51255 1439 51311
rect 1495 51255 1581 51311
rect 1637 51255 1723 51311
rect 1779 51255 1865 51311
rect 1921 51255 2007 51311
rect 2063 51255 2149 51311
rect 2205 51255 2291 51311
rect 2347 51255 2433 51311
rect 2489 51255 2575 51311
rect 2631 51255 2717 51311
rect 2773 51255 2859 51311
rect 2915 51255 3001 51311
rect 3057 51255 3143 51311
rect 3199 51255 3285 51311
rect 3341 51255 3427 51311
rect 3483 51255 3569 51311
rect 3625 51255 3711 51311
rect 3767 51255 3853 51311
rect 3909 51255 3995 51311
rect 4051 51255 4137 51311
rect 4193 51255 4279 51311
rect 4335 51255 4421 51311
rect 4477 51255 4563 51311
rect 4619 51255 4705 51311
rect 4761 51255 4847 51311
rect 4903 51255 4989 51311
rect 5045 51255 5131 51311
rect 5187 51255 5273 51311
rect 5329 51255 5415 51311
rect 5471 51255 5557 51311
rect 5613 51255 5699 51311
rect 5755 51255 5841 51311
rect 5897 51255 5983 51311
rect 6039 51255 6125 51311
rect 6181 51255 6267 51311
rect 6323 51255 6409 51311
rect 6465 51255 6551 51311
rect 6607 51255 6693 51311
rect 6749 51255 6835 51311
rect 6891 51255 6977 51311
rect 7033 51255 7119 51311
rect 7175 51255 7261 51311
rect 7317 51255 7403 51311
rect 7459 51255 7545 51311
rect 7601 51255 7687 51311
rect 7743 51255 7829 51311
rect 7885 51255 7971 51311
rect 8027 51255 8113 51311
rect 8169 51255 8255 51311
rect 8311 51255 8397 51311
rect 8453 51255 8539 51311
rect 8595 51255 8681 51311
rect 8737 51255 8823 51311
rect 8879 51255 8965 51311
rect 9021 51255 9107 51311
rect 9163 51255 9249 51311
rect 9305 51255 9391 51311
rect 9447 51255 9533 51311
rect 9589 51255 9675 51311
rect 9731 51255 9817 51311
rect 9873 51255 9959 51311
rect 10015 51255 10101 51311
rect 10157 51255 10243 51311
rect 10299 51255 10385 51311
rect 10441 51255 10527 51311
rect 10583 51255 10669 51311
rect 10725 51255 10811 51311
rect 10867 51255 10953 51311
rect 11009 51255 11095 51311
rect 11151 51255 11237 51311
rect 11293 51255 11379 51311
rect 11435 51255 11521 51311
rect 11577 51255 11663 51311
rect 11719 51255 11805 51311
rect 11861 51255 11947 51311
rect 12003 51255 12089 51311
rect 12145 51255 12231 51311
rect 12287 51255 12373 51311
rect 12429 51255 12515 51311
rect 12571 51255 12657 51311
rect 12713 51255 12799 51311
rect 12855 51255 12941 51311
rect 12997 51255 13083 51311
rect 13139 51255 13225 51311
rect 13281 51255 13367 51311
rect 13423 51255 13509 51311
rect 13565 51255 13651 51311
rect 13707 51255 13793 51311
rect 13849 51255 13935 51311
rect 13991 51255 14077 51311
rect 14133 51255 14219 51311
rect 14275 51255 14361 51311
rect 14417 51255 14503 51311
rect 14559 51255 14645 51311
rect 14701 51255 14787 51311
rect 14843 51255 15000 51311
rect 0 51169 15000 51255
rect 0 51113 161 51169
rect 217 51113 303 51169
rect 359 51113 445 51169
rect 501 51113 587 51169
rect 643 51113 729 51169
rect 785 51113 871 51169
rect 927 51113 1013 51169
rect 1069 51113 1155 51169
rect 1211 51113 1297 51169
rect 1353 51113 1439 51169
rect 1495 51113 1581 51169
rect 1637 51113 1723 51169
rect 1779 51113 1865 51169
rect 1921 51113 2007 51169
rect 2063 51113 2149 51169
rect 2205 51113 2291 51169
rect 2347 51113 2433 51169
rect 2489 51113 2575 51169
rect 2631 51113 2717 51169
rect 2773 51113 2859 51169
rect 2915 51113 3001 51169
rect 3057 51113 3143 51169
rect 3199 51113 3285 51169
rect 3341 51113 3427 51169
rect 3483 51113 3569 51169
rect 3625 51113 3711 51169
rect 3767 51113 3853 51169
rect 3909 51113 3995 51169
rect 4051 51113 4137 51169
rect 4193 51113 4279 51169
rect 4335 51113 4421 51169
rect 4477 51113 4563 51169
rect 4619 51113 4705 51169
rect 4761 51113 4847 51169
rect 4903 51113 4989 51169
rect 5045 51113 5131 51169
rect 5187 51113 5273 51169
rect 5329 51113 5415 51169
rect 5471 51113 5557 51169
rect 5613 51113 5699 51169
rect 5755 51113 5841 51169
rect 5897 51113 5983 51169
rect 6039 51113 6125 51169
rect 6181 51113 6267 51169
rect 6323 51113 6409 51169
rect 6465 51113 6551 51169
rect 6607 51113 6693 51169
rect 6749 51113 6835 51169
rect 6891 51113 6977 51169
rect 7033 51113 7119 51169
rect 7175 51113 7261 51169
rect 7317 51113 7403 51169
rect 7459 51113 7545 51169
rect 7601 51113 7687 51169
rect 7743 51113 7829 51169
rect 7885 51113 7971 51169
rect 8027 51113 8113 51169
rect 8169 51113 8255 51169
rect 8311 51113 8397 51169
rect 8453 51113 8539 51169
rect 8595 51113 8681 51169
rect 8737 51113 8823 51169
rect 8879 51113 8965 51169
rect 9021 51113 9107 51169
rect 9163 51113 9249 51169
rect 9305 51113 9391 51169
rect 9447 51113 9533 51169
rect 9589 51113 9675 51169
rect 9731 51113 9817 51169
rect 9873 51113 9959 51169
rect 10015 51113 10101 51169
rect 10157 51113 10243 51169
rect 10299 51113 10385 51169
rect 10441 51113 10527 51169
rect 10583 51113 10669 51169
rect 10725 51113 10811 51169
rect 10867 51113 10953 51169
rect 11009 51113 11095 51169
rect 11151 51113 11237 51169
rect 11293 51113 11379 51169
rect 11435 51113 11521 51169
rect 11577 51113 11663 51169
rect 11719 51113 11805 51169
rect 11861 51113 11947 51169
rect 12003 51113 12089 51169
rect 12145 51113 12231 51169
rect 12287 51113 12373 51169
rect 12429 51113 12515 51169
rect 12571 51113 12657 51169
rect 12713 51113 12799 51169
rect 12855 51113 12941 51169
rect 12997 51113 13083 51169
rect 13139 51113 13225 51169
rect 13281 51113 13367 51169
rect 13423 51113 13509 51169
rect 13565 51113 13651 51169
rect 13707 51113 13793 51169
rect 13849 51113 13935 51169
rect 13991 51113 14077 51169
rect 14133 51113 14219 51169
rect 14275 51113 14361 51169
rect 14417 51113 14503 51169
rect 14559 51113 14645 51169
rect 14701 51113 14787 51169
rect 14843 51113 15000 51169
rect 0 51027 15000 51113
rect 0 50971 161 51027
rect 217 50971 303 51027
rect 359 50971 445 51027
rect 501 50971 587 51027
rect 643 50971 729 51027
rect 785 50971 871 51027
rect 927 50971 1013 51027
rect 1069 50971 1155 51027
rect 1211 50971 1297 51027
rect 1353 50971 1439 51027
rect 1495 50971 1581 51027
rect 1637 50971 1723 51027
rect 1779 50971 1865 51027
rect 1921 50971 2007 51027
rect 2063 50971 2149 51027
rect 2205 50971 2291 51027
rect 2347 50971 2433 51027
rect 2489 50971 2575 51027
rect 2631 50971 2717 51027
rect 2773 50971 2859 51027
rect 2915 50971 3001 51027
rect 3057 50971 3143 51027
rect 3199 50971 3285 51027
rect 3341 50971 3427 51027
rect 3483 50971 3569 51027
rect 3625 50971 3711 51027
rect 3767 50971 3853 51027
rect 3909 50971 3995 51027
rect 4051 50971 4137 51027
rect 4193 50971 4279 51027
rect 4335 50971 4421 51027
rect 4477 50971 4563 51027
rect 4619 50971 4705 51027
rect 4761 50971 4847 51027
rect 4903 50971 4989 51027
rect 5045 50971 5131 51027
rect 5187 50971 5273 51027
rect 5329 50971 5415 51027
rect 5471 50971 5557 51027
rect 5613 50971 5699 51027
rect 5755 50971 5841 51027
rect 5897 50971 5983 51027
rect 6039 50971 6125 51027
rect 6181 50971 6267 51027
rect 6323 50971 6409 51027
rect 6465 50971 6551 51027
rect 6607 50971 6693 51027
rect 6749 50971 6835 51027
rect 6891 50971 6977 51027
rect 7033 50971 7119 51027
rect 7175 50971 7261 51027
rect 7317 50971 7403 51027
rect 7459 50971 7545 51027
rect 7601 50971 7687 51027
rect 7743 50971 7829 51027
rect 7885 50971 7971 51027
rect 8027 50971 8113 51027
rect 8169 50971 8255 51027
rect 8311 50971 8397 51027
rect 8453 50971 8539 51027
rect 8595 50971 8681 51027
rect 8737 50971 8823 51027
rect 8879 50971 8965 51027
rect 9021 50971 9107 51027
rect 9163 50971 9249 51027
rect 9305 50971 9391 51027
rect 9447 50971 9533 51027
rect 9589 50971 9675 51027
rect 9731 50971 9817 51027
rect 9873 50971 9959 51027
rect 10015 50971 10101 51027
rect 10157 50971 10243 51027
rect 10299 50971 10385 51027
rect 10441 50971 10527 51027
rect 10583 50971 10669 51027
rect 10725 50971 10811 51027
rect 10867 50971 10953 51027
rect 11009 50971 11095 51027
rect 11151 50971 11237 51027
rect 11293 50971 11379 51027
rect 11435 50971 11521 51027
rect 11577 50971 11663 51027
rect 11719 50971 11805 51027
rect 11861 50971 11947 51027
rect 12003 50971 12089 51027
rect 12145 50971 12231 51027
rect 12287 50971 12373 51027
rect 12429 50971 12515 51027
rect 12571 50971 12657 51027
rect 12713 50971 12799 51027
rect 12855 50971 12941 51027
rect 12997 50971 13083 51027
rect 13139 50971 13225 51027
rect 13281 50971 13367 51027
rect 13423 50971 13509 51027
rect 13565 50971 13651 51027
rect 13707 50971 13793 51027
rect 13849 50971 13935 51027
rect 13991 50971 14077 51027
rect 14133 50971 14219 51027
rect 14275 50971 14361 51027
rect 14417 50971 14503 51027
rect 14559 50971 14645 51027
rect 14701 50971 14787 51027
rect 14843 50971 15000 51027
rect 0 50885 15000 50971
rect 0 50829 161 50885
rect 217 50829 303 50885
rect 359 50829 445 50885
rect 501 50829 587 50885
rect 643 50829 729 50885
rect 785 50829 871 50885
rect 927 50829 1013 50885
rect 1069 50829 1155 50885
rect 1211 50829 1297 50885
rect 1353 50829 1439 50885
rect 1495 50829 1581 50885
rect 1637 50829 1723 50885
rect 1779 50829 1865 50885
rect 1921 50829 2007 50885
rect 2063 50829 2149 50885
rect 2205 50829 2291 50885
rect 2347 50829 2433 50885
rect 2489 50829 2575 50885
rect 2631 50829 2717 50885
rect 2773 50829 2859 50885
rect 2915 50829 3001 50885
rect 3057 50829 3143 50885
rect 3199 50829 3285 50885
rect 3341 50829 3427 50885
rect 3483 50829 3569 50885
rect 3625 50829 3711 50885
rect 3767 50829 3853 50885
rect 3909 50829 3995 50885
rect 4051 50829 4137 50885
rect 4193 50829 4279 50885
rect 4335 50829 4421 50885
rect 4477 50829 4563 50885
rect 4619 50829 4705 50885
rect 4761 50829 4847 50885
rect 4903 50829 4989 50885
rect 5045 50829 5131 50885
rect 5187 50829 5273 50885
rect 5329 50829 5415 50885
rect 5471 50829 5557 50885
rect 5613 50829 5699 50885
rect 5755 50829 5841 50885
rect 5897 50829 5983 50885
rect 6039 50829 6125 50885
rect 6181 50829 6267 50885
rect 6323 50829 6409 50885
rect 6465 50829 6551 50885
rect 6607 50829 6693 50885
rect 6749 50829 6835 50885
rect 6891 50829 6977 50885
rect 7033 50829 7119 50885
rect 7175 50829 7261 50885
rect 7317 50829 7403 50885
rect 7459 50829 7545 50885
rect 7601 50829 7687 50885
rect 7743 50829 7829 50885
rect 7885 50829 7971 50885
rect 8027 50829 8113 50885
rect 8169 50829 8255 50885
rect 8311 50829 8397 50885
rect 8453 50829 8539 50885
rect 8595 50829 8681 50885
rect 8737 50829 8823 50885
rect 8879 50829 8965 50885
rect 9021 50829 9107 50885
rect 9163 50829 9249 50885
rect 9305 50829 9391 50885
rect 9447 50829 9533 50885
rect 9589 50829 9675 50885
rect 9731 50829 9817 50885
rect 9873 50829 9959 50885
rect 10015 50829 10101 50885
rect 10157 50829 10243 50885
rect 10299 50829 10385 50885
rect 10441 50829 10527 50885
rect 10583 50829 10669 50885
rect 10725 50829 10811 50885
rect 10867 50829 10953 50885
rect 11009 50829 11095 50885
rect 11151 50829 11237 50885
rect 11293 50829 11379 50885
rect 11435 50829 11521 50885
rect 11577 50829 11663 50885
rect 11719 50829 11805 50885
rect 11861 50829 11947 50885
rect 12003 50829 12089 50885
rect 12145 50829 12231 50885
rect 12287 50829 12373 50885
rect 12429 50829 12515 50885
rect 12571 50829 12657 50885
rect 12713 50829 12799 50885
rect 12855 50829 12941 50885
rect 12997 50829 13083 50885
rect 13139 50829 13225 50885
rect 13281 50829 13367 50885
rect 13423 50829 13509 50885
rect 13565 50829 13651 50885
rect 13707 50829 13793 50885
rect 13849 50829 13935 50885
rect 13991 50829 14077 50885
rect 14133 50829 14219 50885
rect 14275 50829 14361 50885
rect 14417 50829 14503 50885
rect 14559 50829 14645 50885
rect 14701 50829 14787 50885
rect 14843 50829 15000 50885
rect 0 50800 15000 50829
rect 0 50563 15000 50600
rect 0 50507 161 50563
rect 217 50507 303 50563
rect 359 50507 445 50563
rect 501 50507 587 50563
rect 643 50507 729 50563
rect 785 50507 871 50563
rect 927 50507 1013 50563
rect 1069 50507 1155 50563
rect 1211 50507 1297 50563
rect 1353 50507 1439 50563
rect 1495 50507 1581 50563
rect 1637 50507 1723 50563
rect 1779 50507 1865 50563
rect 1921 50507 2007 50563
rect 2063 50507 2149 50563
rect 2205 50507 2291 50563
rect 2347 50507 2433 50563
rect 2489 50507 2575 50563
rect 2631 50507 2717 50563
rect 2773 50507 2859 50563
rect 2915 50507 3001 50563
rect 3057 50507 3143 50563
rect 3199 50507 3285 50563
rect 3341 50507 3427 50563
rect 3483 50507 3569 50563
rect 3625 50507 3711 50563
rect 3767 50507 3853 50563
rect 3909 50507 3995 50563
rect 4051 50507 4137 50563
rect 4193 50507 4279 50563
rect 4335 50507 4421 50563
rect 4477 50507 4563 50563
rect 4619 50507 4705 50563
rect 4761 50507 4847 50563
rect 4903 50507 4989 50563
rect 5045 50507 5131 50563
rect 5187 50507 5273 50563
rect 5329 50507 5415 50563
rect 5471 50507 5557 50563
rect 5613 50507 5699 50563
rect 5755 50507 5841 50563
rect 5897 50507 5983 50563
rect 6039 50507 6125 50563
rect 6181 50507 6267 50563
rect 6323 50507 6409 50563
rect 6465 50507 6551 50563
rect 6607 50507 6693 50563
rect 6749 50507 6835 50563
rect 6891 50507 6977 50563
rect 7033 50507 7119 50563
rect 7175 50507 7261 50563
rect 7317 50507 7403 50563
rect 7459 50507 7545 50563
rect 7601 50507 7687 50563
rect 7743 50507 7829 50563
rect 7885 50507 7971 50563
rect 8027 50507 8113 50563
rect 8169 50507 8255 50563
rect 8311 50507 8397 50563
rect 8453 50507 8539 50563
rect 8595 50507 8681 50563
rect 8737 50507 8823 50563
rect 8879 50507 8965 50563
rect 9021 50507 9107 50563
rect 9163 50507 9249 50563
rect 9305 50507 9391 50563
rect 9447 50507 9533 50563
rect 9589 50507 9675 50563
rect 9731 50507 9817 50563
rect 9873 50507 9959 50563
rect 10015 50507 10101 50563
rect 10157 50507 10243 50563
rect 10299 50507 10385 50563
rect 10441 50507 10527 50563
rect 10583 50507 10669 50563
rect 10725 50507 10811 50563
rect 10867 50507 10953 50563
rect 11009 50507 11095 50563
rect 11151 50507 11237 50563
rect 11293 50507 11379 50563
rect 11435 50507 11521 50563
rect 11577 50507 11663 50563
rect 11719 50507 11805 50563
rect 11861 50507 11947 50563
rect 12003 50507 12089 50563
rect 12145 50507 12231 50563
rect 12287 50507 12373 50563
rect 12429 50507 12515 50563
rect 12571 50507 12657 50563
rect 12713 50507 12799 50563
rect 12855 50507 12941 50563
rect 12997 50507 13083 50563
rect 13139 50507 13225 50563
rect 13281 50507 13367 50563
rect 13423 50507 13509 50563
rect 13565 50507 13651 50563
rect 13707 50507 13793 50563
rect 13849 50507 13935 50563
rect 13991 50507 14077 50563
rect 14133 50507 14219 50563
rect 14275 50507 14361 50563
rect 14417 50507 14503 50563
rect 14559 50507 14645 50563
rect 14701 50507 14787 50563
rect 14843 50507 15000 50563
rect 0 50421 15000 50507
rect 0 50365 161 50421
rect 217 50365 303 50421
rect 359 50365 445 50421
rect 501 50365 587 50421
rect 643 50365 729 50421
rect 785 50365 871 50421
rect 927 50365 1013 50421
rect 1069 50365 1155 50421
rect 1211 50365 1297 50421
rect 1353 50365 1439 50421
rect 1495 50365 1581 50421
rect 1637 50365 1723 50421
rect 1779 50365 1865 50421
rect 1921 50365 2007 50421
rect 2063 50365 2149 50421
rect 2205 50365 2291 50421
rect 2347 50365 2433 50421
rect 2489 50365 2575 50421
rect 2631 50365 2717 50421
rect 2773 50365 2859 50421
rect 2915 50365 3001 50421
rect 3057 50365 3143 50421
rect 3199 50365 3285 50421
rect 3341 50365 3427 50421
rect 3483 50365 3569 50421
rect 3625 50365 3711 50421
rect 3767 50365 3853 50421
rect 3909 50365 3995 50421
rect 4051 50365 4137 50421
rect 4193 50365 4279 50421
rect 4335 50365 4421 50421
rect 4477 50365 4563 50421
rect 4619 50365 4705 50421
rect 4761 50365 4847 50421
rect 4903 50365 4989 50421
rect 5045 50365 5131 50421
rect 5187 50365 5273 50421
rect 5329 50365 5415 50421
rect 5471 50365 5557 50421
rect 5613 50365 5699 50421
rect 5755 50365 5841 50421
rect 5897 50365 5983 50421
rect 6039 50365 6125 50421
rect 6181 50365 6267 50421
rect 6323 50365 6409 50421
rect 6465 50365 6551 50421
rect 6607 50365 6693 50421
rect 6749 50365 6835 50421
rect 6891 50365 6977 50421
rect 7033 50365 7119 50421
rect 7175 50365 7261 50421
rect 7317 50365 7403 50421
rect 7459 50365 7545 50421
rect 7601 50365 7687 50421
rect 7743 50365 7829 50421
rect 7885 50365 7971 50421
rect 8027 50365 8113 50421
rect 8169 50365 8255 50421
rect 8311 50365 8397 50421
rect 8453 50365 8539 50421
rect 8595 50365 8681 50421
rect 8737 50365 8823 50421
rect 8879 50365 8965 50421
rect 9021 50365 9107 50421
rect 9163 50365 9249 50421
rect 9305 50365 9391 50421
rect 9447 50365 9533 50421
rect 9589 50365 9675 50421
rect 9731 50365 9817 50421
rect 9873 50365 9959 50421
rect 10015 50365 10101 50421
rect 10157 50365 10243 50421
rect 10299 50365 10385 50421
rect 10441 50365 10527 50421
rect 10583 50365 10669 50421
rect 10725 50365 10811 50421
rect 10867 50365 10953 50421
rect 11009 50365 11095 50421
rect 11151 50365 11237 50421
rect 11293 50365 11379 50421
rect 11435 50365 11521 50421
rect 11577 50365 11663 50421
rect 11719 50365 11805 50421
rect 11861 50365 11947 50421
rect 12003 50365 12089 50421
rect 12145 50365 12231 50421
rect 12287 50365 12373 50421
rect 12429 50365 12515 50421
rect 12571 50365 12657 50421
rect 12713 50365 12799 50421
rect 12855 50365 12941 50421
rect 12997 50365 13083 50421
rect 13139 50365 13225 50421
rect 13281 50365 13367 50421
rect 13423 50365 13509 50421
rect 13565 50365 13651 50421
rect 13707 50365 13793 50421
rect 13849 50365 13935 50421
rect 13991 50365 14077 50421
rect 14133 50365 14219 50421
rect 14275 50365 14361 50421
rect 14417 50365 14503 50421
rect 14559 50365 14645 50421
rect 14701 50365 14787 50421
rect 14843 50365 15000 50421
rect 0 50279 15000 50365
rect 0 50223 161 50279
rect 217 50223 303 50279
rect 359 50223 445 50279
rect 501 50223 587 50279
rect 643 50223 729 50279
rect 785 50223 871 50279
rect 927 50223 1013 50279
rect 1069 50223 1155 50279
rect 1211 50223 1297 50279
rect 1353 50223 1439 50279
rect 1495 50223 1581 50279
rect 1637 50223 1723 50279
rect 1779 50223 1865 50279
rect 1921 50223 2007 50279
rect 2063 50223 2149 50279
rect 2205 50223 2291 50279
rect 2347 50223 2433 50279
rect 2489 50223 2575 50279
rect 2631 50223 2717 50279
rect 2773 50223 2859 50279
rect 2915 50223 3001 50279
rect 3057 50223 3143 50279
rect 3199 50223 3285 50279
rect 3341 50223 3427 50279
rect 3483 50223 3569 50279
rect 3625 50223 3711 50279
rect 3767 50223 3853 50279
rect 3909 50223 3995 50279
rect 4051 50223 4137 50279
rect 4193 50223 4279 50279
rect 4335 50223 4421 50279
rect 4477 50223 4563 50279
rect 4619 50223 4705 50279
rect 4761 50223 4847 50279
rect 4903 50223 4989 50279
rect 5045 50223 5131 50279
rect 5187 50223 5273 50279
rect 5329 50223 5415 50279
rect 5471 50223 5557 50279
rect 5613 50223 5699 50279
rect 5755 50223 5841 50279
rect 5897 50223 5983 50279
rect 6039 50223 6125 50279
rect 6181 50223 6267 50279
rect 6323 50223 6409 50279
rect 6465 50223 6551 50279
rect 6607 50223 6693 50279
rect 6749 50223 6835 50279
rect 6891 50223 6977 50279
rect 7033 50223 7119 50279
rect 7175 50223 7261 50279
rect 7317 50223 7403 50279
rect 7459 50223 7545 50279
rect 7601 50223 7687 50279
rect 7743 50223 7829 50279
rect 7885 50223 7971 50279
rect 8027 50223 8113 50279
rect 8169 50223 8255 50279
rect 8311 50223 8397 50279
rect 8453 50223 8539 50279
rect 8595 50223 8681 50279
rect 8737 50223 8823 50279
rect 8879 50223 8965 50279
rect 9021 50223 9107 50279
rect 9163 50223 9249 50279
rect 9305 50223 9391 50279
rect 9447 50223 9533 50279
rect 9589 50223 9675 50279
rect 9731 50223 9817 50279
rect 9873 50223 9959 50279
rect 10015 50223 10101 50279
rect 10157 50223 10243 50279
rect 10299 50223 10385 50279
rect 10441 50223 10527 50279
rect 10583 50223 10669 50279
rect 10725 50223 10811 50279
rect 10867 50223 10953 50279
rect 11009 50223 11095 50279
rect 11151 50223 11237 50279
rect 11293 50223 11379 50279
rect 11435 50223 11521 50279
rect 11577 50223 11663 50279
rect 11719 50223 11805 50279
rect 11861 50223 11947 50279
rect 12003 50223 12089 50279
rect 12145 50223 12231 50279
rect 12287 50223 12373 50279
rect 12429 50223 12515 50279
rect 12571 50223 12657 50279
rect 12713 50223 12799 50279
rect 12855 50223 12941 50279
rect 12997 50223 13083 50279
rect 13139 50223 13225 50279
rect 13281 50223 13367 50279
rect 13423 50223 13509 50279
rect 13565 50223 13651 50279
rect 13707 50223 13793 50279
rect 13849 50223 13935 50279
rect 13991 50223 14077 50279
rect 14133 50223 14219 50279
rect 14275 50223 14361 50279
rect 14417 50223 14503 50279
rect 14559 50223 14645 50279
rect 14701 50223 14787 50279
rect 14843 50223 15000 50279
rect 0 50137 15000 50223
rect 0 50081 161 50137
rect 217 50081 303 50137
rect 359 50081 445 50137
rect 501 50081 587 50137
rect 643 50081 729 50137
rect 785 50081 871 50137
rect 927 50081 1013 50137
rect 1069 50081 1155 50137
rect 1211 50081 1297 50137
rect 1353 50081 1439 50137
rect 1495 50081 1581 50137
rect 1637 50081 1723 50137
rect 1779 50081 1865 50137
rect 1921 50081 2007 50137
rect 2063 50081 2149 50137
rect 2205 50081 2291 50137
rect 2347 50081 2433 50137
rect 2489 50081 2575 50137
rect 2631 50081 2717 50137
rect 2773 50081 2859 50137
rect 2915 50081 3001 50137
rect 3057 50081 3143 50137
rect 3199 50081 3285 50137
rect 3341 50081 3427 50137
rect 3483 50081 3569 50137
rect 3625 50081 3711 50137
rect 3767 50081 3853 50137
rect 3909 50081 3995 50137
rect 4051 50081 4137 50137
rect 4193 50081 4279 50137
rect 4335 50081 4421 50137
rect 4477 50081 4563 50137
rect 4619 50081 4705 50137
rect 4761 50081 4847 50137
rect 4903 50081 4989 50137
rect 5045 50081 5131 50137
rect 5187 50081 5273 50137
rect 5329 50081 5415 50137
rect 5471 50081 5557 50137
rect 5613 50081 5699 50137
rect 5755 50081 5841 50137
rect 5897 50081 5983 50137
rect 6039 50081 6125 50137
rect 6181 50081 6267 50137
rect 6323 50081 6409 50137
rect 6465 50081 6551 50137
rect 6607 50081 6693 50137
rect 6749 50081 6835 50137
rect 6891 50081 6977 50137
rect 7033 50081 7119 50137
rect 7175 50081 7261 50137
rect 7317 50081 7403 50137
rect 7459 50081 7545 50137
rect 7601 50081 7687 50137
rect 7743 50081 7829 50137
rect 7885 50081 7971 50137
rect 8027 50081 8113 50137
rect 8169 50081 8255 50137
rect 8311 50081 8397 50137
rect 8453 50081 8539 50137
rect 8595 50081 8681 50137
rect 8737 50081 8823 50137
rect 8879 50081 8965 50137
rect 9021 50081 9107 50137
rect 9163 50081 9249 50137
rect 9305 50081 9391 50137
rect 9447 50081 9533 50137
rect 9589 50081 9675 50137
rect 9731 50081 9817 50137
rect 9873 50081 9959 50137
rect 10015 50081 10101 50137
rect 10157 50081 10243 50137
rect 10299 50081 10385 50137
rect 10441 50081 10527 50137
rect 10583 50081 10669 50137
rect 10725 50081 10811 50137
rect 10867 50081 10953 50137
rect 11009 50081 11095 50137
rect 11151 50081 11237 50137
rect 11293 50081 11379 50137
rect 11435 50081 11521 50137
rect 11577 50081 11663 50137
rect 11719 50081 11805 50137
rect 11861 50081 11947 50137
rect 12003 50081 12089 50137
rect 12145 50081 12231 50137
rect 12287 50081 12373 50137
rect 12429 50081 12515 50137
rect 12571 50081 12657 50137
rect 12713 50081 12799 50137
rect 12855 50081 12941 50137
rect 12997 50081 13083 50137
rect 13139 50081 13225 50137
rect 13281 50081 13367 50137
rect 13423 50081 13509 50137
rect 13565 50081 13651 50137
rect 13707 50081 13793 50137
rect 13849 50081 13935 50137
rect 13991 50081 14077 50137
rect 14133 50081 14219 50137
rect 14275 50081 14361 50137
rect 14417 50081 14503 50137
rect 14559 50081 14645 50137
rect 14701 50081 14787 50137
rect 14843 50081 15000 50137
rect 0 49995 15000 50081
rect 0 49939 161 49995
rect 217 49939 303 49995
rect 359 49939 445 49995
rect 501 49939 587 49995
rect 643 49939 729 49995
rect 785 49939 871 49995
rect 927 49939 1013 49995
rect 1069 49939 1155 49995
rect 1211 49939 1297 49995
rect 1353 49939 1439 49995
rect 1495 49939 1581 49995
rect 1637 49939 1723 49995
rect 1779 49939 1865 49995
rect 1921 49939 2007 49995
rect 2063 49939 2149 49995
rect 2205 49939 2291 49995
rect 2347 49939 2433 49995
rect 2489 49939 2575 49995
rect 2631 49939 2717 49995
rect 2773 49939 2859 49995
rect 2915 49939 3001 49995
rect 3057 49939 3143 49995
rect 3199 49939 3285 49995
rect 3341 49939 3427 49995
rect 3483 49939 3569 49995
rect 3625 49939 3711 49995
rect 3767 49939 3853 49995
rect 3909 49939 3995 49995
rect 4051 49939 4137 49995
rect 4193 49939 4279 49995
rect 4335 49939 4421 49995
rect 4477 49939 4563 49995
rect 4619 49939 4705 49995
rect 4761 49939 4847 49995
rect 4903 49939 4989 49995
rect 5045 49939 5131 49995
rect 5187 49939 5273 49995
rect 5329 49939 5415 49995
rect 5471 49939 5557 49995
rect 5613 49939 5699 49995
rect 5755 49939 5841 49995
rect 5897 49939 5983 49995
rect 6039 49939 6125 49995
rect 6181 49939 6267 49995
rect 6323 49939 6409 49995
rect 6465 49939 6551 49995
rect 6607 49939 6693 49995
rect 6749 49939 6835 49995
rect 6891 49939 6977 49995
rect 7033 49939 7119 49995
rect 7175 49939 7261 49995
rect 7317 49939 7403 49995
rect 7459 49939 7545 49995
rect 7601 49939 7687 49995
rect 7743 49939 7829 49995
rect 7885 49939 7971 49995
rect 8027 49939 8113 49995
rect 8169 49939 8255 49995
rect 8311 49939 8397 49995
rect 8453 49939 8539 49995
rect 8595 49939 8681 49995
rect 8737 49939 8823 49995
rect 8879 49939 8965 49995
rect 9021 49939 9107 49995
rect 9163 49939 9249 49995
rect 9305 49939 9391 49995
rect 9447 49939 9533 49995
rect 9589 49939 9675 49995
rect 9731 49939 9817 49995
rect 9873 49939 9959 49995
rect 10015 49939 10101 49995
rect 10157 49939 10243 49995
rect 10299 49939 10385 49995
rect 10441 49939 10527 49995
rect 10583 49939 10669 49995
rect 10725 49939 10811 49995
rect 10867 49939 10953 49995
rect 11009 49939 11095 49995
rect 11151 49939 11237 49995
rect 11293 49939 11379 49995
rect 11435 49939 11521 49995
rect 11577 49939 11663 49995
rect 11719 49939 11805 49995
rect 11861 49939 11947 49995
rect 12003 49939 12089 49995
rect 12145 49939 12231 49995
rect 12287 49939 12373 49995
rect 12429 49939 12515 49995
rect 12571 49939 12657 49995
rect 12713 49939 12799 49995
rect 12855 49939 12941 49995
rect 12997 49939 13083 49995
rect 13139 49939 13225 49995
rect 13281 49939 13367 49995
rect 13423 49939 13509 49995
rect 13565 49939 13651 49995
rect 13707 49939 13793 49995
rect 13849 49939 13935 49995
rect 13991 49939 14077 49995
rect 14133 49939 14219 49995
rect 14275 49939 14361 49995
rect 14417 49939 14503 49995
rect 14559 49939 14645 49995
rect 14701 49939 14787 49995
rect 14843 49939 15000 49995
rect 0 49853 15000 49939
rect 0 49797 161 49853
rect 217 49797 303 49853
rect 359 49797 445 49853
rect 501 49797 587 49853
rect 643 49797 729 49853
rect 785 49797 871 49853
rect 927 49797 1013 49853
rect 1069 49797 1155 49853
rect 1211 49797 1297 49853
rect 1353 49797 1439 49853
rect 1495 49797 1581 49853
rect 1637 49797 1723 49853
rect 1779 49797 1865 49853
rect 1921 49797 2007 49853
rect 2063 49797 2149 49853
rect 2205 49797 2291 49853
rect 2347 49797 2433 49853
rect 2489 49797 2575 49853
rect 2631 49797 2717 49853
rect 2773 49797 2859 49853
rect 2915 49797 3001 49853
rect 3057 49797 3143 49853
rect 3199 49797 3285 49853
rect 3341 49797 3427 49853
rect 3483 49797 3569 49853
rect 3625 49797 3711 49853
rect 3767 49797 3853 49853
rect 3909 49797 3995 49853
rect 4051 49797 4137 49853
rect 4193 49797 4279 49853
rect 4335 49797 4421 49853
rect 4477 49797 4563 49853
rect 4619 49797 4705 49853
rect 4761 49797 4847 49853
rect 4903 49797 4989 49853
rect 5045 49797 5131 49853
rect 5187 49797 5273 49853
rect 5329 49797 5415 49853
rect 5471 49797 5557 49853
rect 5613 49797 5699 49853
rect 5755 49797 5841 49853
rect 5897 49797 5983 49853
rect 6039 49797 6125 49853
rect 6181 49797 6267 49853
rect 6323 49797 6409 49853
rect 6465 49797 6551 49853
rect 6607 49797 6693 49853
rect 6749 49797 6835 49853
rect 6891 49797 6977 49853
rect 7033 49797 7119 49853
rect 7175 49797 7261 49853
rect 7317 49797 7403 49853
rect 7459 49797 7545 49853
rect 7601 49797 7687 49853
rect 7743 49797 7829 49853
rect 7885 49797 7971 49853
rect 8027 49797 8113 49853
rect 8169 49797 8255 49853
rect 8311 49797 8397 49853
rect 8453 49797 8539 49853
rect 8595 49797 8681 49853
rect 8737 49797 8823 49853
rect 8879 49797 8965 49853
rect 9021 49797 9107 49853
rect 9163 49797 9249 49853
rect 9305 49797 9391 49853
rect 9447 49797 9533 49853
rect 9589 49797 9675 49853
rect 9731 49797 9817 49853
rect 9873 49797 9959 49853
rect 10015 49797 10101 49853
rect 10157 49797 10243 49853
rect 10299 49797 10385 49853
rect 10441 49797 10527 49853
rect 10583 49797 10669 49853
rect 10725 49797 10811 49853
rect 10867 49797 10953 49853
rect 11009 49797 11095 49853
rect 11151 49797 11237 49853
rect 11293 49797 11379 49853
rect 11435 49797 11521 49853
rect 11577 49797 11663 49853
rect 11719 49797 11805 49853
rect 11861 49797 11947 49853
rect 12003 49797 12089 49853
rect 12145 49797 12231 49853
rect 12287 49797 12373 49853
rect 12429 49797 12515 49853
rect 12571 49797 12657 49853
rect 12713 49797 12799 49853
rect 12855 49797 12941 49853
rect 12997 49797 13083 49853
rect 13139 49797 13225 49853
rect 13281 49797 13367 49853
rect 13423 49797 13509 49853
rect 13565 49797 13651 49853
rect 13707 49797 13793 49853
rect 13849 49797 13935 49853
rect 13991 49797 14077 49853
rect 14133 49797 14219 49853
rect 14275 49797 14361 49853
rect 14417 49797 14503 49853
rect 14559 49797 14645 49853
rect 14701 49797 14787 49853
rect 14843 49797 15000 49853
rect 0 49711 15000 49797
rect 0 49655 161 49711
rect 217 49655 303 49711
rect 359 49655 445 49711
rect 501 49655 587 49711
rect 643 49655 729 49711
rect 785 49655 871 49711
rect 927 49655 1013 49711
rect 1069 49655 1155 49711
rect 1211 49655 1297 49711
rect 1353 49655 1439 49711
rect 1495 49655 1581 49711
rect 1637 49655 1723 49711
rect 1779 49655 1865 49711
rect 1921 49655 2007 49711
rect 2063 49655 2149 49711
rect 2205 49655 2291 49711
rect 2347 49655 2433 49711
rect 2489 49655 2575 49711
rect 2631 49655 2717 49711
rect 2773 49655 2859 49711
rect 2915 49655 3001 49711
rect 3057 49655 3143 49711
rect 3199 49655 3285 49711
rect 3341 49655 3427 49711
rect 3483 49655 3569 49711
rect 3625 49655 3711 49711
rect 3767 49655 3853 49711
rect 3909 49655 3995 49711
rect 4051 49655 4137 49711
rect 4193 49655 4279 49711
rect 4335 49655 4421 49711
rect 4477 49655 4563 49711
rect 4619 49655 4705 49711
rect 4761 49655 4847 49711
rect 4903 49655 4989 49711
rect 5045 49655 5131 49711
rect 5187 49655 5273 49711
rect 5329 49655 5415 49711
rect 5471 49655 5557 49711
rect 5613 49655 5699 49711
rect 5755 49655 5841 49711
rect 5897 49655 5983 49711
rect 6039 49655 6125 49711
rect 6181 49655 6267 49711
rect 6323 49655 6409 49711
rect 6465 49655 6551 49711
rect 6607 49655 6693 49711
rect 6749 49655 6835 49711
rect 6891 49655 6977 49711
rect 7033 49655 7119 49711
rect 7175 49655 7261 49711
rect 7317 49655 7403 49711
rect 7459 49655 7545 49711
rect 7601 49655 7687 49711
rect 7743 49655 7829 49711
rect 7885 49655 7971 49711
rect 8027 49655 8113 49711
rect 8169 49655 8255 49711
rect 8311 49655 8397 49711
rect 8453 49655 8539 49711
rect 8595 49655 8681 49711
rect 8737 49655 8823 49711
rect 8879 49655 8965 49711
rect 9021 49655 9107 49711
rect 9163 49655 9249 49711
rect 9305 49655 9391 49711
rect 9447 49655 9533 49711
rect 9589 49655 9675 49711
rect 9731 49655 9817 49711
rect 9873 49655 9959 49711
rect 10015 49655 10101 49711
rect 10157 49655 10243 49711
rect 10299 49655 10385 49711
rect 10441 49655 10527 49711
rect 10583 49655 10669 49711
rect 10725 49655 10811 49711
rect 10867 49655 10953 49711
rect 11009 49655 11095 49711
rect 11151 49655 11237 49711
rect 11293 49655 11379 49711
rect 11435 49655 11521 49711
rect 11577 49655 11663 49711
rect 11719 49655 11805 49711
rect 11861 49655 11947 49711
rect 12003 49655 12089 49711
rect 12145 49655 12231 49711
rect 12287 49655 12373 49711
rect 12429 49655 12515 49711
rect 12571 49655 12657 49711
rect 12713 49655 12799 49711
rect 12855 49655 12941 49711
rect 12997 49655 13083 49711
rect 13139 49655 13225 49711
rect 13281 49655 13367 49711
rect 13423 49655 13509 49711
rect 13565 49655 13651 49711
rect 13707 49655 13793 49711
rect 13849 49655 13935 49711
rect 13991 49655 14077 49711
rect 14133 49655 14219 49711
rect 14275 49655 14361 49711
rect 14417 49655 14503 49711
rect 14559 49655 14645 49711
rect 14701 49655 14787 49711
rect 14843 49655 15000 49711
rect 0 49569 15000 49655
rect 0 49513 161 49569
rect 217 49513 303 49569
rect 359 49513 445 49569
rect 501 49513 587 49569
rect 643 49513 729 49569
rect 785 49513 871 49569
rect 927 49513 1013 49569
rect 1069 49513 1155 49569
rect 1211 49513 1297 49569
rect 1353 49513 1439 49569
rect 1495 49513 1581 49569
rect 1637 49513 1723 49569
rect 1779 49513 1865 49569
rect 1921 49513 2007 49569
rect 2063 49513 2149 49569
rect 2205 49513 2291 49569
rect 2347 49513 2433 49569
rect 2489 49513 2575 49569
rect 2631 49513 2717 49569
rect 2773 49513 2859 49569
rect 2915 49513 3001 49569
rect 3057 49513 3143 49569
rect 3199 49513 3285 49569
rect 3341 49513 3427 49569
rect 3483 49513 3569 49569
rect 3625 49513 3711 49569
rect 3767 49513 3853 49569
rect 3909 49513 3995 49569
rect 4051 49513 4137 49569
rect 4193 49513 4279 49569
rect 4335 49513 4421 49569
rect 4477 49513 4563 49569
rect 4619 49513 4705 49569
rect 4761 49513 4847 49569
rect 4903 49513 4989 49569
rect 5045 49513 5131 49569
rect 5187 49513 5273 49569
rect 5329 49513 5415 49569
rect 5471 49513 5557 49569
rect 5613 49513 5699 49569
rect 5755 49513 5841 49569
rect 5897 49513 5983 49569
rect 6039 49513 6125 49569
rect 6181 49513 6267 49569
rect 6323 49513 6409 49569
rect 6465 49513 6551 49569
rect 6607 49513 6693 49569
rect 6749 49513 6835 49569
rect 6891 49513 6977 49569
rect 7033 49513 7119 49569
rect 7175 49513 7261 49569
rect 7317 49513 7403 49569
rect 7459 49513 7545 49569
rect 7601 49513 7687 49569
rect 7743 49513 7829 49569
rect 7885 49513 7971 49569
rect 8027 49513 8113 49569
rect 8169 49513 8255 49569
rect 8311 49513 8397 49569
rect 8453 49513 8539 49569
rect 8595 49513 8681 49569
rect 8737 49513 8823 49569
rect 8879 49513 8965 49569
rect 9021 49513 9107 49569
rect 9163 49513 9249 49569
rect 9305 49513 9391 49569
rect 9447 49513 9533 49569
rect 9589 49513 9675 49569
rect 9731 49513 9817 49569
rect 9873 49513 9959 49569
rect 10015 49513 10101 49569
rect 10157 49513 10243 49569
rect 10299 49513 10385 49569
rect 10441 49513 10527 49569
rect 10583 49513 10669 49569
rect 10725 49513 10811 49569
rect 10867 49513 10953 49569
rect 11009 49513 11095 49569
rect 11151 49513 11237 49569
rect 11293 49513 11379 49569
rect 11435 49513 11521 49569
rect 11577 49513 11663 49569
rect 11719 49513 11805 49569
rect 11861 49513 11947 49569
rect 12003 49513 12089 49569
rect 12145 49513 12231 49569
rect 12287 49513 12373 49569
rect 12429 49513 12515 49569
rect 12571 49513 12657 49569
rect 12713 49513 12799 49569
rect 12855 49513 12941 49569
rect 12997 49513 13083 49569
rect 13139 49513 13225 49569
rect 13281 49513 13367 49569
rect 13423 49513 13509 49569
rect 13565 49513 13651 49569
rect 13707 49513 13793 49569
rect 13849 49513 13935 49569
rect 13991 49513 14077 49569
rect 14133 49513 14219 49569
rect 14275 49513 14361 49569
rect 14417 49513 14503 49569
rect 14559 49513 14645 49569
rect 14701 49513 14787 49569
rect 14843 49513 15000 49569
rect 0 49427 15000 49513
rect 0 49371 161 49427
rect 217 49371 303 49427
rect 359 49371 445 49427
rect 501 49371 587 49427
rect 643 49371 729 49427
rect 785 49371 871 49427
rect 927 49371 1013 49427
rect 1069 49371 1155 49427
rect 1211 49371 1297 49427
rect 1353 49371 1439 49427
rect 1495 49371 1581 49427
rect 1637 49371 1723 49427
rect 1779 49371 1865 49427
rect 1921 49371 2007 49427
rect 2063 49371 2149 49427
rect 2205 49371 2291 49427
rect 2347 49371 2433 49427
rect 2489 49371 2575 49427
rect 2631 49371 2717 49427
rect 2773 49371 2859 49427
rect 2915 49371 3001 49427
rect 3057 49371 3143 49427
rect 3199 49371 3285 49427
rect 3341 49371 3427 49427
rect 3483 49371 3569 49427
rect 3625 49371 3711 49427
rect 3767 49371 3853 49427
rect 3909 49371 3995 49427
rect 4051 49371 4137 49427
rect 4193 49371 4279 49427
rect 4335 49371 4421 49427
rect 4477 49371 4563 49427
rect 4619 49371 4705 49427
rect 4761 49371 4847 49427
rect 4903 49371 4989 49427
rect 5045 49371 5131 49427
rect 5187 49371 5273 49427
rect 5329 49371 5415 49427
rect 5471 49371 5557 49427
rect 5613 49371 5699 49427
rect 5755 49371 5841 49427
rect 5897 49371 5983 49427
rect 6039 49371 6125 49427
rect 6181 49371 6267 49427
rect 6323 49371 6409 49427
rect 6465 49371 6551 49427
rect 6607 49371 6693 49427
rect 6749 49371 6835 49427
rect 6891 49371 6977 49427
rect 7033 49371 7119 49427
rect 7175 49371 7261 49427
rect 7317 49371 7403 49427
rect 7459 49371 7545 49427
rect 7601 49371 7687 49427
rect 7743 49371 7829 49427
rect 7885 49371 7971 49427
rect 8027 49371 8113 49427
rect 8169 49371 8255 49427
rect 8311 49371 8397 49427
rect 8453 49371 8539 49427
rect 8595 49371 8681 49427
rect 8737 49371 8823 49427
rect 8879 49371 8965 49427
rect 9021 49371 9107 49427
rect 9163 49371 9249 49427
rect 9305 49371 9391 49427
rect 9447 49371 9533 49427
rect 9589 49371 9675 49427
rect 9731 49371 9817 49427
rect 9873 49371 9959 49427
rect 10015 49371 10101 49427
rect 10157 49371 10243 49427
rect 10299 49371 10385 49427
rect 10441 49371 10527 49427
rect 10583 49371 10669 49427
rect 10725 49371 10811 49427
rect 10867 49371 10953 49427
rect 11009 49371 11095 49427
rect 11151 49371 11237 49427
rect 11293 49371 11379 49427
rect 11435 49371 11521 49427
rect 11577 49371 11663 49427
rect 11719 49371 11805 49427
rect 11861 49371 11947 49427
rect 12003 49371 12089 49427
rect 12145 49371 12231 49427
rect 12287 49371 12373 49427
rect 12429 49371 12515 49427
rect 12571 49371 12657 49427
rect 12713 49371 12799 49427
rect 12855 49371 12941 49427
rect 12997 49371 13083 49427
rect 13139 49371 13225 49427
rect 13281 49371 13367 49427
rect 13423 49371 13509 49427
rect 13565 49371 13651 49427
rect 13707 49371 13793 49427
rect 13849 49371 13935 49427
rect 13991 49371 14077 49427
rect 14133 49371 14219 49427
rect 14275 49371 14361 49427
rect 14417 49371 14503 49427
rect 14559 49371 14645 49427
rect 14701 49371 14787 49427
rect 14843 49371 15000 49427
rect 0 49285 15000 49371
rect 0 49229 161 49285
rect 217 49229 303 49285
rect 359 49229 445 49285
rect 501 49229 587 49285
rect 643 49229 729 49285
rect 785 49229 871 49285
rect 927 49229 1013 49285
rect 1069 49229 1155 49285
rect 1211 49229 1297 49285
rect 1353 49229 1439 49285
rect 1495 49229 1581 49285
rect 1637 49229 1723 49285
rect 1779 49229 1865 49285
rect 1921 49229 2007 49285
rect 2063 49229 2149 49285
rect 2205 49229 2291 49285
rect 2347 49229 2433 49285
rect 2489 49229 2575 49285
rect 2631 49229 2717 49285
rect 2773 49229 2859 49285
rect 2915 49229 3001 49285
rect 3057 49229 3143 49285
rect 3199 49229 3285 49285
rect 3341 49229 3427 49285
rect 3483 49229 3569 49285
rect 3625 49229 3711 49285
rect 3767 49229 3853 49285
rect 3909 49229 3995 49285
rect 4051 49229 4137 49285
rect 4193 49229 4279 49285
rect 4335 49229 4421 49285
rect 4477 49229 4563 49285
rect 4619 49229 4705 49285
rect 4761 49229 4847 49285
rect 4903 49229 4989 49285
rect 5045 49229 5131 49285
rect 5187 49229 5273 49285
rect 5329 49229 5415 49285
rect 5471 49229 5557 49285
rect 5613 49229 5699 49285
rect 5755 49229 5841 49285
rect 5897 49229 5983 49285
rect 6039 49229 6125 49285
rect 6181 49229 6267 49285
rect 6323 49229 6409 49285
rect 6465 49229 6551 49285
rect 6607 49229 6693 49285
rect 6749 49229 6835 49285
rect 6891 49229 6977 49285
rect 7033 49229 7119 49285
rect 7175 49229 7261 49285
rect 7317 49229 7403 49285
rect 7459 49229 7545 49285
rect 7601 49229 7687 49285
rect 7743 49229 7829 49285
rect 7885 49229 7971 49285
rect 8027 49229 8113 49285
rect 8169 49229 8255 49285
rect 8311 49229 8397 49285
rect 8453 49229 8539 49285
rect 8595 49229 8681 49285
rect 8737 49229 8823 49285
rect 8879 49229 8965 49285
rect 9021 49229 9107 49285
rect 9163 49229 9249 49285
rect 9305 49229 9391 49285
rect 9447 49229 9533 49285
rect 9589 49229 9675 49285
rect 9731 49229 9817 49285
rect 9873 49229 9959 49285
rect 10015 49229 10101 49285
rect 10157 49229 10243 49285
rect 10299 49229 10385 49285
rect 10441 49229 10527 49285
rect 10583 49229 10669 49285
rect 10725 49229 10811 49285
rect 10867 49229 10953 49285
rect 11009 49229 11095 49285
rect 11151 49229 11237 49285
rect 11293 49229 11379 49285
rect 11435 49229 11521 49285
rect 11577 49229 11663 49285
rect 11719 49229 11805 49285
rect 11861 49229 11947 49285
rect 12003 49229 12089 49285
rect 12145 49229 12231 49285
rect 12287 49229 12373 49285
rect 12429 49229 12515 49285
rect 12571 49229 12657 49285
rect 12713 49229 12799 49285
rect 12855 49229 12941 49285
rect 12997 49229 13083 49285
rect 13139 49229 13225 49285
rect 13281 49229 13367 49285
rect 13423 49229 13509 49285
rect 13565 49229 13651 49285
rect 13707 49229 13793 49285
rect 13849 49229 13935 49285
rect 13991 49229 14077 49285
rect 14133 49229 14219 49285
rect 14275 49229 14361 49285
rect 14417 49229 14503 49285
rect 14559 49229 14645 49285
rect 14701 49229 14787 49285
rect 14843 49229 15000 49285
rect 0 49200 15000 49229
rect 0 48941 15000 49000
rect 0 48885 161 48941
rect 217 48885 303 48941
rect 359 48885 445 48941
rect 501 48885 587 48941
rect 643 48885 729 48941
rect 785 48885 871 48941
rect 927 48885 1013 48941
rect 1069 48885 1155 48941
rect 1211 48885 1297 48941
rect 1353 48885 1439 48941
rect 1495 48885 1581 48941
rect 1637 48885 1723 48941
rect 1779 48885 1865 48941
rect 1921 48885 2007 48941
rect 2063 48885 2149 48941
rect 2205 48885 2291 48941
rect 2347 48885 2433 48941
rect 2489 48885 2575 48941
rect 2631 48885 2717 48941
rect 2773 48885 2859 48941
rect 2915 48885 3001 48941
rect 3057 48885 3143 48941
rect 3199 48885 3285 48941
rect 3341 48885 3427 48941
rect 3483 48885 3569 48941
rect 3625 48885 3711 48941
rect 3767 48885 3853 48941
rect 3909 48885 3995 48941
rect 4051 48885 4137 48941
rect 4193 48885 4279 48941
rect 4335 48885 4421 48941
rect 4477 48885 4563 48941
rect 4619 48885 4705 48941
rect 4761 48885 4847 48941
rect 4903 48885 4989 48941
rect 5045 48885 5131 48941
rect 5187 48885 5273 48941
rect 5329 48885 5415 48941
rect 5471 48885 5557 48941
rect 5613 48885 5699 48941
rect 5755 48885 5841 48941
rect 5897 48885 5983 48941
rect 6039 48885 6125 48941
rect 6181 48885 6267 48941
rect 6323 48885 6409 48941
rect 6465 48885 6551 48941
rect 6607 48885 6693 48941
rect 6749 48885 6835 48941
rect 6891 48885 6977 48941
rect 7033 48885 7119 48941
rect 7175 48885 7261 48941
rect 7317 48885 7403 48941
rect 7459 48885 7545 48941
rect 7601 48885 7687 48941
rect 7743 48885 7829 48941
rect 7885 48885 7971 48941
rect 8027 48885 8113 48941
rect 8169 48885 8255 48941
rect 8311 48885 8397 48941
rect 8453 48885 8539 48941
rect 8595 48885 8681 48941
rect 8737 48885 8823 48941
rect 8879 48885 8965 48941
rect 9021 48885 9107 48941
rect 9163 48885 9249 48941
rect 9305 48885 9391 48941
rect 9447 48885 9533 48941
rect 9589 48885 9675 48941
rect 9731 48885 9817 48941
rect 9873 48885 9959 48941
rect 10015 48885 10101 48941
rect 10157 48885 10243 48941
rect 10299 48885 10385 48941
rect 10441 48885 10527 48941
rect 10583 48885 10669 48941
rect 10725 48885 10811 48941
rect 10867 48885 10953 48941
rect 11009 48885 11095 48941
rect 11151 48885 11237 48941
rect 11293 48885 11379 48941
rect 11435 48885 11521 48941
rect 11577 48885 11663 48941
rect 11719 48885 11805 48941
rect 11861 48885 11947 48941
rect 12003 48885 12089 48941
rect 12145 48885 12231 48941
rect 12287 48885 12373 48941
rect 12429 48885 12515 48941
rect 12571 48885 12657 48941
rect 12713 48885 12799 48941
rect 12855 48885 12941 48941
rect 12997 48885 13083 48941
rect 13139 48885 13225 48941
rect 13281 48885 13367 48941
rect 13423 48885 13509 48941
rect 13565 48885 13651 48941
rect 13707 48885 13793 48941
rect 13849 48885 13935 48941
rect 13991 48885 14077 48941
rect 14133 48885 14219 48941
rect 14275 48885 14361 48941
rect 14417 48885 14503 48941
rect 14559 48885 14645 48941
rect 14701 48885 14787 48941
rect 14843 48885 15000 48941
rect 0 48799 15000 48885
rect 0 48743 161 48799
rect 217 48743 303 48799
rect 359 48743 445 48799
rect 501 48743 587 48799
rect 643 48743 729 48799
rect 785 48743 871 48799
rect 927 48743 1013 48799
rect 1069 48743 1155 48799
rect 1211 48743 1297 48799
rect 1353 48743 1439 48799
rect 1495 48743 1581 48799
rect 1637 48743 1723 48799
rect 1779 48743 1865 48799
rect 1921 48743 2007 48799
rect 2063 48743 2149 48799
rect 2205 48743 2291 48799
rect 2347 48743 2433 48799
rect 2489 48743 2575 48799
rect 2631 48743 2717 48799
rect 2773 48743 2859 48799
rect 2915 48743 3001 48799
rect 3057 48743 3143 48799
rect 3199 48743 3285 48799
rect 3341 48743 3427 48799
rect 3483 48743 3569 48799
rect 3625 48743 3711 48799
rect 3767 48743 3853 48799
rect 3909 48743 3995 48799
rect 4051 48743 4137 48799
rect 4193 48743 4279 48799
rect 4335 48743 4421 48799
rect 4477 48743 4563 48799
rect 4619 48743 4705 48799
rect 4761 48743 4847 48799
rect 4903 48743 4989 48799
rect 5045 48743 5131 48799
rect 5187 48743 5273 48799
rect 5329 48743 5415 48799
rect 5471 48743 5557 48799
rect 5613 48743 5699 48799
rect 5755 48743 5841 48799
rect 5897 48743 5983 48799
rect 6039 48743 6125 48799
rect 6181 48743 6267 48799
rect 6323 48743 6409 48799
rect 6465 48743 6551 48799
rect 6607 48743 6693 48799
rect 6749 48743 6835 48799
rect 6891 48743 6977 48799
rect 7033 48743 7119 48799
rect 7175 48743 7261 48799
rect 7317 48743 7403 48799
rect 7459 48743 7545 48799
rect 7601 48743 7687 48799
rect 7743 48743 7829 48799
rect 7885 48743 7971 48799
rect 8027 48743 8113 48799
rect 8169 48743 8255 48799
rect 8311 48743 8397 48799
rect 8453 48743 8539 48799
rect 8595 48743 8681 48799
rect 8737 48743 8823 48799
rect 8879 48743 8965 48799
rect 9021 48743 9107 48799
rect 9163 48743 9249 48799
rect 9305 48743 9391 48799
rect 9447 48743 9533 48799
rect 9589 48743 9675 48799
rect 9731 48743 9817 48799
rect 9873 48743 9959 48799
rect 10015 48743 10101 48799
rect 10157 48743 10243 48799
rect 10299 48743 10385 48799
rect 10441 48743 10527 48799
rect 10583 48743 10669 48799
rect 10725 48743 10811 48799
rect 10867 48743 10953 48799
rect 11009 48743 11095 48799
rect 11151 48743 11237 48799
rect 11293 48743 11379 48799
rect 11435 48743 11521 48799
rect 11577 48743 11663 48799
rect 11719 48743 11805 48799
rect 11861 48743 11947 48799
rect 12003 48743 12089 48799
rect 12145 48743 12231 48799
rect 12287 48743 12373 48799
rect 12429 48743 12515 48799
rect 12571 48743 12657 48799
rect 12713 48743 12799 48799
rect 12855 48743 12941 48799
rect 12997 48743 13083 48799
rect 13139 48743 13225 48799
rect 13281 48743 13367 48799
rect 13423 48743 13509 48799
rect 13565 48743 13651 48799
rect 13707 48743 13793 48799
rect 13849 48743 13935 48799
rect 13991 48743 14077 48799
rect 14133 48743 14219 48799
rect 14275 48743 14361 48799
rect 14417 48743 14503 48799
rect 14559 48743 14645 48799
rect 14701 48743 14787 48799
rect 14843 48743 15000 48799
rect 0 48657 15000 48743
rect 0 48601 161 48657
rect 217 48601 303 48657
rect 359 48601 445 48657
rect 501 48601 587 48657
rect 643 48601 729 48657
rect 785 48601 871 48657
rect 927 48601 1013 48657
rect 1069 48601 1155 48657
rect 1211 48601 1297 48657
rect 1353 48601 1439 48657
rect 1495 48601 1581 48657
rect 1637 48601 1723 48657
rect 1779 48601 1865 48657
rect 1921 48601 2007 48657
rect 2063 48601 2149 48657
rect 2205 48601 2291 48657
rect 2347 48601 2433 48657
rect 2489 48601 2575 48657
rect 2631 48601 2717 48657
rect 2773 48601 2859 48657
rect 2915 48601 3001 48657
rect 3057 48601 3143 48657
rect 3199 48601 3285 48657
rect 3341 48601 3427 48657
rect 3483 48601 3569 48657
rect 3625 48601 3711 48657
rect 3767 48601 3853 48657
rect 3909 48601 3995 48657
rect 4051 48601 4137 48657
rect 4193 48601 4279 48657
rect 4335 48601 4421 48657
rect 4477 48601 4563 48657
rect 4619 48601 4705 48657
rect 4761 48601 4847 48657
rect 4903 48601 4989 48657
rect 5045 48601 5131 48657
rect 5187 48601 5273 48657
rect 5329 48601 5415 48657
rect 5471 48601 5557 48657
rect 5613 48601 5699 48657
rect 5755 48601 5841 48657
rect 5897 48601 5983 48657
rect 6039 48601 6125 48657
rect 6181 48601 6267 48657
rect 6323 48601 6409 48657
rect 6465 48601 6551 48657
rect 6607 48601 6693 48657
rect 6749 48601 6835 48657
rect 6891 48601 6977 48657
rect 7033 48601 7119 48657
rect 7175 48601 7261 48657
rect 7317 48601 7403 48657
rect 7459 48601 7545 48657
rect 7601 48601 7687 48657
rect 7743 48601 7829 48657
rect 7885 48601 7971 48657
rect 8027 48601 8113 48657
rect 8169 48601 8255 48657
rect 8311 48601 8397 48657
rect 8453 48601 8539 48657
rect 8595 48601 8681 48657
rect 8737 48601 8823 48657
rect 8879 48601 8965 48657
rect 9021 48601 9107 48657
rect 9163 48601 9249 48657
rect 9305 48601 9391 48657
rect 9447 48601 9533 48657
rect 9589 48601 9675 48657
rect 9731 48601 9817 48657
rect 9873 48601 9959 48657
rect 10015 48601 10101 48657
rect 10157 48601 10243 48657
rect 10299 48601 10385 48657
rect 10441 48601 10527 48657
rect 10583 48601 10669 48657
rect 10725 48601 10811 48657
rect 10867 48601 10953 48657
rect 11009 48601 11095 48657
rect 11151 48601 11237 48657
rect 11293 48601 11379 48657
rect 11435 48601 11521 48657
rect 11577 48601 11663 48657
rect 11719 48601 11805 48657
rect 11861 48601 11947 48657
rect 12003 48601 12089 48657
rect 12145 48601 12231 48657
rect 12287 48601 12373 48657
rect 12429 48601 12515 48657
rect 12571 48601 12657 48657
rect 12713 48601 12799 48657
rect 12855 48601 12941 48657
rect 12997 48601 13083 48657
rect 13139 48601 13225 48657
rect 13281 48601 13367 48657
rect 13423 48601 13509 48657
rect 13565 48601 13651 48657
rect 13707 48601 13793 48657
rect 13849 48601 13935 48657
rect 13991 48601 14077 48657
rect 14133 48601 14219 48657
rect 14275 48601 14361 48657
rect 14417 48601 14503 48657
rect 14559 48601 14645 48657
rect 14701 48601 14787 48657
rect 14843 48601 15000 48657
rect 0 48515 15000 48601
rect 0 48459 161 48515
rect 217 48459 303 48515
rect 359 48459 445 48515
rect 501 48459 587 48515
rect 643 48459 729 48515
rect 785 48459 871 48515
rect 927 48459 1013 48515
rect 1069 48459 1155 48515
rect 1211 48459 1297 48515
rect 1353 48459 1439 48515
rect 1495 48459 1581 48515
rect 1637 48459 1723 48515
rect 1779 48459 1865 48515
rect 1921 48459 2007 48515
rect 2063 48459 2149 48515
rect 2205 48459 2291 48515
rect 2347 48459 2433 48515
rect 2489 48459 2575 48515
rect 2631 48459 2717 48515
rect 2773 48459 2859 48515
rect 2915 48459 3001 48515
rect 3057 48459 3143 48515
rect 3199 48459 3285 48515
rect 3341 48459 3427 48515
rect 3483 48459 3569 48515
rect 3625 48459 3711 48515
rect 3767 48459 3853 48515
rect 3909 48459 3995 48515
rect 4051 48459 4137 48515
rect 4193 48459 4279 48515
rect 4335 48459 4421 48515
rect 4477 48459 4563 48515
rect 4619 48459 4705 48515
rect 4761 48459 4847 48515
rect 4903 48459 4989 48515
rect 5045 48459 5131 48515
rect 5187 48459 5273 48515
rect 5329 48459 5415 48515
rect 5471 48459 5557 48515
rect 5613 48459 5699 48515
rect 5755 48459 5841 48515
rect 5897 48459 5983 48515
rect 6039 48459 6125 48515
rect 6181 48459 6267 48515
rect 6323 48459 6409 48515
rect 6465 48459 6551 48515
rect 6607 48459 6693 48515
rect 6749 48459 6835 48515
rect 6891 48459 6977 48515
rect 7033 48459 7119 48515
rect 7175 48459 7261 48515
rect 7317 48459 7403 48515
rect 7459 48459 7545 48515
rect 7601 48459 7687 48515
rect 7743 48459 7829 48515
rect 7885 48459 7971 48515
rect 8027 48459 8113 48515
rect 8169 48459 8255 48515
rect 8311 48459 8397 48515
rect 8453 48459 8539 48515
rect 8595 48459 8681 48515
rect 8737 48459 8823 48515
rect 8879 48459 8965 48515
rect 9021 48459 9107 48515
rect 9163 48459 9249 48515
rect 9305 48459 9391 48515
rect 9447 48459 9533 48515
rect 9589 48459 9675 48515
rect 9731 48459 9817 48515
rect 9873 48459 9959 48515
rect 10015 48459 10101 48515
rect 10157 48459 10243 48515
rect 10299 48459 10385 48515
rect 10441 48459 10527 48515
rect 10583 48459 10669 48515
rect 10725 48459 10811 48515
rect 10867 48459 10953 48515
rect 11009 48459 11095 48515
rect 11151 48459 11237 48515
rect 11293 48459 11379 48515
rect 11435 48459 11521 48515
rect 11577 48459 11663 48515
rect 11719 48459 11805 48515
rect 11861 48459 11947 48515
rect 12003 48459 12089 48515
rect 12145 48459 12231 48515
rect 12287 48459 12373 48515
rect 12429 48459 12515 48515
rect 12571 48459 12657 48515
rect 12713 48459 12799 48515
rect 12855 48459 12941 48515
rect 12997 48459 13083 48515
rect 13139 48459 13225 48515
rect 13281 48459 13367 48515
rect 13423 48459 13509 48515
rect 13565 48459 13651 48515
rect 13707 48459 13793 48515
rect 13849 48459 13935 48515
rect 13991 48459 14077 48515
rect 14133 48459 14219 48515
rect 14275 48459 14361 48515
rect 14417 48459 14503 48515
rect 14559 48459 14645 48515
rect 14701 48459 14787 48515
rect 14843 48459 15000 48515
rect 0 48373 15000 48459
rect 0 48317 161 48373
rect 217 48317 303 48373
rect 359 48317 445 48373
rect 501 48317 587 48373
rect 643 48317 729 48373
rect 785 48317 871 48373
rect 927 48317 1013 48373
rect 1069 48317 1155 48373
rect 1211 48317 1297 48373
rect 1353 48317 1439 48373
rect 1495 48317 1581 48373
rect 1637 48317 1723 48373
rect 1779 48317 1865 48373
rect 1921 48317 2007 48373
rect 2063 48317 2149 48373
rect 2205 48317 2291 48373
rect 2347 48317 2433 48373
rect 2489 48317 2575 48373
rect 2631 48317 2717 48373
rect 2773 48317 2859 48373
rect 2915 48317 3001 48373
rect 3057 48317 3143 48373
rect 3199 48317 3285 48373
rect 3341 48317 3427 48373
rect 3483 48317 3569 48373
rect 3625 48317 3711 48373
rect 3767 48317 3853 48373
rect 3909 48317 3995 48373
rect 4051 48317 4137 48373
rect 4193 48317 4279 48373
rect 4335 48317 4421 48373
rect 4477 48317 4563 48373
rect 4619 48317 4705 48373
rect 4761 48317 4847 48373
rect 4903 48317 4989 48373
rect 5045 48317 5131 48373
rect 5187 48317 5273 48373
rect 5329 48317 5415 48373
rect 5471 48317 5557 48373
rect 5613 48317 5699 48373
rect 5755 48317 5841 48373
rect 5897 48317 5983 48373
rect 6039 48317 6125 48373
rect 6181 48317 6267 48373
rect 6323 48317 6409 48373
rect 6465 48317 6551 48373
rect 6607 48317 6693 48373
rect 6749 48317 6835 48373
rect 6891 48317 6977 48373
rect 7033 48317 7119 48373
rect 7175 48317 7261 48373
rect 7317 48317 7403 48373
rect 7459 48317 7545 48373
rect 7601 48317 7687 48373
rect 7743 48317 7829 48373
rect 7885 48317 7971 48373
rect 8027 48317 8113 48373
rect 8169 48317 8255 48373
rect 8311 48317 8397 48373
rect 8453 48317 8539 48373
rect 8595 48317 8681 48373
rect 8737 48317 8823 48373
rect 8879 48317 8965 48373
rect 9021 48317 9107 48373
rect 9163 48317 9249 48373
rect 9305 48317 9391 48373
rect 9447 48317 9533 48373
rect 9589 48317 9675 48373
rect 9731 48317 9817 48373
rect 9873 48317 9959 48373
rect 10015 48317 10101 48373
rect 10157 48317 10243 48373
rect 10299 48317 10385 48373
rect 10441 48317 10527 48373
rect 10583 48317 10669 48373
rect 10725 48317 10811 48373
rect 10867 48317 10953 48373
rect 11009 48317 11095 48373
rect 11151 48317 11237 48373
rect 11293 48317 11379 48373
rect 11435 48317 11521 48373
rect 11577 48317 11663 48373
rect 11719 48317 11805 48373
rect 11861 48317 11947 48373
rect 12003 48317 12089 48373
rect 12145 48317 12231 48373
rect 12287 48317 12373 48373
rect 12429 48317 12515 48373
rect 12571 48317 12657 48373
rect 12713 48317 12799 48373
rect 12855 48317 12941 48373
rect 12997 48317 13083 48373
rect 13139 48317 13225 48373
rect 13281 48317 13367 48373
rect 13423 48317 13509 48373
rect 13565 48317 13651 48373
rect 13707 48317 13793 48373
rect 13849 48317 13935 48373
rect 13991 48317 14077 48373
rect 14133 48317 14219 48373
rect 14275 48317 14361 48373
rect 14417 48317 14503 48373
rect 14559 48317 14645 48373
rect 14701 48317 14787 48373
rect 14843 48317 15000 48373
rect 0 48231 15000 48317
rect 0 48175 161 48231
rect 217 48175 303 48231
rect 359 48175 445 48231
rect 501 48175 587 48231
rect 643 48175 729 48231
rect 785 48175 871 48231
rect 927 48175 1013 48231
rect 1069 48175 1155 48231
rect 1211 48175 1297 48231
rect 1353 48175 1439 48231
rect 1495 48175 1581 48231
rect 1637 48175 1723 48231
rect 1779 48175 1865 48231
rect 1921 48175 2007 48231
rect 2063 48175 2149 48231
rect 2205 48175 2291 48231
rect 2347 48175 2433 48231
rect 2489 48175 2575 48231
rect 2631 48175 2717 48231
rect 2773 48175 2859 48231
rect 2915 48175 3001 48231
rect 3057 48175 3143 48231
rect 3199 48175 3285 48231
rect 3341 48175 3427 48231
rect 3483 48175 3569 48231
rect 3625 48175 3711 48231
rect 3767 48175 3853 48231
rect 3909 48175 3995 48231
rect 4051 48175 4137 48231
rect 4193 48175 4279 48231
rect 4335 48175 4421 48231
rect 4477 48175 4563 48231
rect 4619 48175 4705 48231
rect 4761 48175 4847 48231
rect 4903 48175 4989 48231
rect 5045 48175 5131 48231
rect 5187 48175 5273 48231
rect 5329 48175 5415 48231
rect 5471 48175 5557 48231
rect 5613 48175 5699 48231
rect 5755 48175 5841 48231
rect 5897 48175 5983 48231
rect 6039 48175 6125 48231
rect 6181 48175 6267 48231
rect 6323 48175 6409 48231
rect 6465 48175 6551 48231
rect 6607 48175 6693 48231
rect 6749 48175 6835 48231
rect 6891 48175 6977 48231
rect 7033 48175 7119 48231
rect 7175 48175 7261 48231
rect 7317 48175 7403 48231
rect 7459 48175 7545 48231
rect 7601 48175 7687 48231
rect 7743 48175 7829 48231
rect 7885 48175 7971 48231
rect 8027 48175 8113 48231
rect 8169 48175 8255 48231
rect 8311 48175 8397 48231
rect 8453 48175 8539 48231
rect 8595 48175 8681 48231
rect 8737 48175 8823 48231
rect 8879 48175 8965 48231
rect 9021 48175 9107 48231
rect 9163 48175 9249 48231
rect 9305 48175 9391 48231
rect 9447 48175 9533 48231
rect 9589 48175 9675 48231
rect 9731 48175 9817 48231
rect 9873 48175 9959 48231
rect 10015 48175 10101 48231
rect 10157 48175 10243 48231
rect 10299 48175 10385 48231
rect 10441 48175 10527 48231
rect 10583 48175 10669 48231
rect 10725 48175 10811 48231
rect 10867 48175 10953 48231
rect 11009 48175 11095 48231
rect 11151 48175 11237 48231
rect 11293 48175 11379 48231
rect 11435 48175 11521 48231
rect 11577 48175 11663 48231
rect 11719 48175 11805 48231
rect 11861 48175 11947 48231
rect 12003 48175 12089 48231
rect 12145 48175 12231 48231
rect 12287 48175 12373 48231
rect 12429 48175 12515 48231
rect 12571 48175 12657 48231
rect 12713 48175 12799 48231
rect 12855 48175 12941 48231
rect 12997 48175 13083 48231
rect 13139 48175 13225 48231
rect 13281 48175 13367 48231
rect 13423 48175 13509 48231
rect 13565 48175 13651 48231
rect 13707 48175 13793 48231
rect 13849 48175 13935 48231
rect 13991 48175 14077 48231
rect 14133 48175 14219 48231
rect 14275 48175 14361 48231
rect 14417 48175 14503 48231
rect 14559 48175 14645 48231
rect 14701 48175 14787 48231
rect 14843 48175 15000 48231
rect 0 48089 15000 48175
rect 0 48033 161 48089
rect 217 48033 303 48089
rect 359 48033 445 48089
rect 501 48033 587 48089
rect 643 48033 729 48089
rect 785 48033 871 48089
rect 927 48033 1013 48089
rect 1069 48033 1155 48089
rect 1211 48033 1297 48089
rect 1353 48033 1439 48089
rect 1495 48033 1581 48089
rect 1637 48033 1723 48089
rect 1779 48033 1865 48089
rect 1921 48033 2007 48089
rect 2063 48033 2149 48089
rect 2205 48033 2291 48089
rect 2347 48033 2433 48089
rect 2489 48033 2575 48089
rect 2631 48033 2717 48089
rect 2773 48033 2859 48089
rect 2915 48033 3001 48089
rect 3057 48033 3143 48089
rect 3199 48033 3285 48089
rect 3341 48033 3427 48089
rect 3483 48033 3569 48089
rect 3625 48033 3711 48089
rect 3767 48033 3853 48089
rect 3909 48033 3995 48089
rect 4051 48033 4137 48089
rect 4193 48033 4279 48089
rect 4335 48033 4421 48089
rect 4477 48033 4563 48089
rect 4619 48033 4705 48089
rect 4761 48033 4847 48089
rect 4903 48033 4989 48089
rect 5045 48033 5131 48089
rect 5187 48033 5273 48089
rect 5329 48033 5415 48089
rect 5471 48033 5557 48089
rect 5613 48033 5699 48089
rect 5755 48033 5841 48089
rect 5897 48033 5983 48089
rect 6039 48033 6125 48089
rect 6181 48033 6267 48089
rect 6323 48033 6409 48089
rect 6465 48033 6551 48089
rect 6607 48033 6693 48089
rect 6749 48033 6835 48089
rect 6891 48033 6977 48089
rect 7033 48033 7119 48089
rect 7175 48033 7261 48089
rect 7317 48033 7403 48089
rect 7459 48033 7545 48089
rect 7601 48033 7687 48089
rect 7743 48033 7829 48089
rect 7885 48033 7971 48089
rect 8027 48033 8113 48089
rect 8169 48033 8255 48089
rect 8311 48033 8397 48089
rect 8453 48033 8539 48089
rect 8595 48033 8681 48089
rect 8737 48033 8823 48089
rect 8879 48033 8965 48089
rect 9021 48033 9107 48089
rect 9163 48033 9249 48089
rect 9305 48033 9391 48089
rect 9447 48033 9533 48089
rect 9589 48033 9675 48089
rect 9731 48033 9817 48089
rect 9873 48033 9959 48089
rect 10015 48033 10101 48089
rect 10157 48033 10243 48089
rect 10299 48033 10385 48089
rect 10441 48033 10527 48089
rect 10583 48033 10669 48089
rect 10725 48033 10811 48089
rect 10867 48033 10953 48089
rect 11009 48033 11095 48089
rect 11151 48033 11237 48089
rect 11293 48033 11379 48089
rect 11435 48033 11521 48089
rect 11577 48033 11663 48089
rect 11719 48033 11805 48089
rect 11861 48033 11947 48089
rect 12003 48033 12089 48089
rect 12145 48033 12231 48089
rect 12287 48033 12373 48089
rect 12429 48033 12515 48089
rect 12571 48033 12657 48089
rect 12713 48033 12799 48089
rect 12855 48033 12941 48089
rect 12997 48033 13083 48089
rect 13139 48033 13225 48089
rect 13281 48033 13367 48089
rect 13423 48033 13509 48089
rect 13565 48033 13651 48089
rect 13707 48033 13793 48089
rect 13849 48033 13935 48089
rect 13991 48033 14077 48089
rect 14133 48033 14219 48089
rect 14275 48033 14361 48089
rect 14417 48033 14503 48089
rect 14559 48033 14645 48089
rect 14701 48033 14787 48089
rect 14843 48033 15000 48089
rect 0 47947 15000 48033
rect 0 47891 161 47947
rect 217 47891 303 47947
rect 359 47891 445 47947
rect 501 47891 587 47947
rect 643 47891 729 47947
rect 785 47891 871 47947
rect 927 47891 1013 47947
rect 1069 47891 1155 47947
rect 1211 47891 1297 47947
rect 1353 47891 1439 47947
rect 1495 47891 1581 47947
rect 1637 47891 1723 47947
rect 1779 47891 1865 47947
rect 1921 47891 2007 47947
rect 2063 47891 2149 47947
rect 2205 47891 2291 47947
rect 2347 47891 2433 47947
rect 2489 47891 2575 47947
rect 2631 47891 2717 47947
rect 2773 47891 2859 47947
rect 2915 47891 3001 47947
rect 3057 47891 3143 47947
rect 3199 47891 3285 47947
rect 3341 47891 3427 47947
rect 3483 47891 3569 47947
rect 3625 47891 3711 47947
rect 3767 47891 3853 47947
rect 3909 47891 3995 47947
rect 4051 47891 4137 47947
rect 4193 47891 4279 47947
rect 4335 47891 4421 47947
rect 4477 47891 4563 47947
rect 4619 47891 4705 47947
rect 4761 47891 4847 47947
rect 4903 47891 4989 47947
rect 5045 47891 5131 47947
rect 5187 47891 5273 47947
rect 5329 47891 5415 47947
rect 5471 47891 5557 47947
rect 5613 47891 5699 47947
rect 5755 47891 5841 47947
rect 5897 47891 5983 47947
rect 6039 47891 6125 47947
rect 6181 47891 6267 47947
rect 6323 47891 6409 47947
rect 6465 47891 6551 47947
rect 6607 47891 6693 47947
rect 6749 47891 6835 47947
rect 6891 47891 6977 47947
rect 7033 47891 7119 47947
rect 7175 47891 7261 47947
rect 7317 47891 7403 47947
rect 7459 47891 7545 47947
rect 7601 47891 7687 47947
rect 7743 47891 7829 47947
rect 7885 47891 7971 47947
rect 8027 47891 8113 47947
rect 8169 47891 8255 47947
rect 8311 47891 8397 47947
rect 8453 47891 8539 47947
rect 8595 47891 8681 47947
rect 8737 47891 8823 47947
rect 8879 47891 8965 47947
rect 9021 47891 9107 47947
rect 9163 47891 9249 47947
rect 9305 47891 9391 47947
rect 9447 47891 9533 47947
rect 9589 47891 9675 47947
rect 9731 47891 9817 47947
rect 9873 47891 9959 47947
rect 10015 47891 10101 47947
rect 10157 47891 10243 47947
rect 10299 47891 10385 47947
rect 10441 47891 10527 47947
rect 10583 47891 10669 47947
rect 10725 47891 10811 47947
rect 10867 47891 10953 47947
rect 11009 47891 11095 47947
rect 11151 47891 11237 47947
rect 11293 47891 11379 47947
rect 11435 47891 11521 47947
rect 11577 47891 11663 47947
rect 11719 47891 11805 47947
rect 11861 47891 11947 47947
rect 12003 47891 12089 47947
rect 12145 47891 12231 47947
rect 12287 47891 12373 47947
rect 12429 47891 12515 47947
rect 12571 47891 12657 47947
rect 12713 47891 12799 47947
rect 12855 47891 12941 47947
rect 12997 47891 13083 47947
rect 13139 47891 13225 47947
rect 13281 47891 13367 47947
rect 13423 47891 13509 47947
rect 13565 47891 13651 47947
rect 13707 47891 13793 47947
rect 13849 47891 13935 47947
rect 13991 47891 14077 47947
rect 14133 47891 14219 47947
rect 14275 47891 14361 47947
rect 14417 47891 14503 47947
rect 14559 47891 14645 47947
rect 14701 47891 14787 47947
rect 14843 47891 15000 47947
rect 0 47805 15000 47891
rect 0 47749 161 47805
rect 217 47749 303 47805
rect 359 47749 445 47805
rect 501 47749 587 47805
rect 643 47749 729 47805
rect 785 47749 871 47805
rect 927 47749 1013 47805
rect 1069 47749 1155 47805
rect 1211 47749 1297 47805
rect 1353 47749 1439 47805
rect 1495 47749 1581 47805
rect 1637 47749 1723 47805
rect 1779 47749 1865 47805
rect 1921 47749 2007 47805
rect 2063 47749 2149 47805
rect 2205 47749 2291 47805
rect 2347 47749 2433 47805
rect 2489 47749 2575 47805
rect 2631 47749 2717 47805
rect 2773 47749 2859 47805
rect 2915 47749 3001 47805
rect 3057 47749 3143 47805
rect 3199 47749 3285 47805
rect 3341 47749 3427 47805
rect 3483 47749 3569 47805
rect 3625 47749 3711 47805
rect 3767 47749 3853 47805
rect 3909 47749 3995 47805
rect 4051 47749 4137 47805
rect 4193 47749 4279 47805
rect 4335 47749 4421 47805
rect 4477 47749 4563 47805
rect 4619 47749 4705 47805
rect 4761 47749 4847 47805
rect 4903 47749 4989 47805
rect 5045 47749 5131 47805
rect 5187 47749 5273 47805
rect 5329 47749 5415 47805
rect 5471 47749 5557 47805
rect 5613 47749 5699 47805
rect 5755 47749 5841 47805
rect 5897 47749 5983 47805
rect 6039 47749 6125 47805
rect 6181 47749 6267 47805
rect 6323 47749 6409 47805
rect 6465 47749 6551 47805
rect 6607 47749 6693 47805
rect 6749 47749 6835 47805
rect 6891 47749 6977 47805
rect 7033 47749 7119 47805
rect 7175 47749 7261 47805
rect 7317 47749 7403 47805
rect 7459 47749 7545 47805
rect 7601 47749 7687 47805
rect 7743 47749 7829 47805
rect 7885 47749 7971 47805
rect 8027 47749 8113 47805
rect 8169 47749 8255 47805
rect 8311 47749 8397 47805
rect 8453 47749 8539 47805
rect 8595 47749 8681 47805
rect 8737 47749 8823 47805
rect 8879 47749 8965 47805
rect 9021 47749 9107 47805
rect 9163 47749 9249 47805
rect 9305 47749 9391 47805
rect 9447 47749 9533 47805
rect 9589 47749 9675 47805
rect 9731 47749 9817 47805
rect 9873 47749 9959 47805
rect 10015 47749 10101 47805
rect 10157 47749 10243 47805
rect 10299 47749 10385 47805
rect 10441 47749 10527 47805
rect 10583 47749 10669 47805
rect 10725 47749 10811 47805
rect 10867 47749 10953 47805
rect 11009 47749 11095 47805
rect 11151 47749 11237 47805
rect 11293 47749 11379 47805
rect 11435 47749 11521 47805
rect 11577 47749 11663 47805
rect 11719 47749 11805 47805
rect 11861 47749 11947 47805
rect 12003 47749 12089 47805
rect 12145 47749 12231 47805
rect 12287 47749 12373 47805
rect 12429 47749 12515 47805
rect 12571 47749 12657 47805
rect 12713 47749 12799 47805
rect 12855 47749 12941 47805
rect 12997 47749 13083 47805
rect 13139 47749 13225 47805
rect 13281 47749 13367 47805
rect 13423 47749 13509 47805
rect 13565 47749 13651 47805
rect 13707 47749 13793 47805
rect 13849 47749 13935 47805
rect 13991 47749 14077 47805
rect 14133 47749 14219 47805
rect 14275 47749 14361 47805
rect 14417 47749 14503 47805
rect 14559 47749 14645 47805
rect 14701 47749 14787 47805
rect 14843 47749 15000 47805
rect 0 47663 15000 47749
rect 0 47607 161 47663
rect 217 47607 303 47663
rect 359 47607 445 47663
rect 501 47607 587 47663
rect 643 47607 729 47663
rect 785 47607 871 47663
rect 927 47607 1013 47663
rect 1069 47607 1155 47663
rect 1211 47607 1297 47663
rect 1353 47607 1439 47663
rect 1495 47607 1581 47663
rect 1637 47607 1723 47663
rect 1779 47607 1865 47663
rect 1921 47607 2007 47663
rect 2063 47607 2149 47663
rect 2205 47607 2291 47663
rect 2347 47607 2433 47663
rect 2489 47607 2575 47663
rect 2631 47607 2717 47663
rect 2773 47607 2859 47663
rect 2915 47607 3001 47663
rect 3057 47607 3143 47663
rect 3199 47607 3285 47663
rect 3341 47607 3427 47663
rect 3483 47607 3569 47663
rect 3625 47607 3711 47663
rect 3767 47607 3853 47663
rect 3909 47607 3995 47663
rect 4051 47607 4137 47663
rect 4193 47607 4279 47663
rect 4335 47607 4421 47663
rect 4477 47607 4563 47663
rect 4619 47607 4705 47663
rect 4761 47607 4847 47663
rect 4903 47607 4989 47663
rect 5045 47607 5131 47663
rect 5187 47607 5273 47663
rect 5329 47607 5415 47663
rect 5471 47607 5557 47663
rect 5613 47607 5699 47663
rect 5755 47607 5841 47663
rect 5897 47607 5983 47663
rect 6039 47607 6125 47663
rect 6181 47607 6267 47663
rect 6323 47607 6409 47663
rect 6465 47607 6551 47663
rect 6607 47607 6693 47663
rect 6749 47607 6835 47663
rect 6891 47607 6977 47663
rect 7033 47607 7119 47663
rect 7175 47607 7261 47663
rect 7317 47607 7403 47663
rect 7459 47607 7545 47663
rect 7601 47607 7687 47663
rect 7743 47607 7829 47663
rect 7885 47607 7971 47663
rect 8027 47607 8113 47663
rect 8169 47607 8255 47663
rect 8311 47607 8397 47663
rect 8453 47607 8539 47663
rect 8595 47607 8681 47663
rect 8737 47607 8823 47663
rect 8879 47607 8965 47663
rect 9021 47607 9107 47663
rect 9163 47607 9249 47663
rect 9305 47607 9391 47663
rect 9447 47607 9533 47663
rect 9589 47607 9675 47663
rect 9731 47607 9817 47663
rect 9873 47607 9959 47663
rect 10015 47607 10101 47663
rect 10157 47607 10243 47663
rect 10299 47607 10385 47663
rect 10441 47607 10527 47663
rect 10583 47607 10669 47663
rect 10725 47607 10811 47663
rect 10867 47607 10953 47663
rect 11009 47607 11095 47663
rect 11151 47607 11237 47663
rect 11293 47607 11379 47663
rect 11435 47607 11521 47663
rect 11577 47607 11663 47663
rect 11719 47607 11805 47663
rect 11861 47607 11947 47663
rect 12003 47607 12089 47663
rect 12145 47607 12231 47663
rect 12287 47607 12373 47663
rect 12429 47607 12515 47663
rect 12571 47607 12657 47663
rect 12713 47607 12799 47663
rect 12855 47607 12941 47663
rect 12997 47607 13083 47663
rect 13139 47607 13225 47663
rect 13281 47607 13367 47663
rect 13423 47607 13509 47663
rect 13565 47607 13651 47663
rect 13707 47607 13793 47663
rect 13849 47607 13935 47663
rect 13991 47607 14077 47663
rect 14133 47607 14219 47663
rect 14275 47607 14361 47663
rect 14417 47607 14503 47663
rect 14559 47607 14645 47663
rect 14701 47607 14787 47663
rect 14843 47607 15000 47663
rect 0 47521 15000 47607
rect 0 47465 161 47521
rect 217 47465 303 47521
rect 359 47465 445 47521
rect 501 47465 587 47521
rect 643 47465 729 47521
rect 785 47465 871 47521
rect 927 47465 1013 47521
rect 1069 47465 1155 47521
rect 1211 47465 1297 47521
rect 1353 47465 1439 47521
rect 1495 47465 1581 47521
rect 1637 47465 1723 47521
rect 1779 47465 1865 47521
rect 1921 47465 2007 47521
rect 2063 47465 2149 47521
rect 2205 47465 2291 47521
rect 2347 47465 2433 47521
rect 2489 47465 2575 47521
rect 2631 47465 2717 47521
rect 2773 47465 2859 47521
rect 2915 47465 3001 47521
rect 3057 47465 3143 47521
rect 3199 47465 3285 47521
rect 3341 47465 3427 47521
rect 3483 47465 3569 47521
rect 3625 47465 3711 47521
rect 3767 47465 3853 47521
rect 3909 47465 3995 47521
rect 4051 47465 4137 47521
rect 4193 47465 4279 47521
rect 4335 47465 4421 47521
rect 4477 47465 4563 47521
rect 4619 47465 4705 47521
rect 4761 47465 4847 47521
rect 4903 47465 4989 47521
rect 5045 47465 5131 47521
rect 5187 47465 5273 47521
rect 5329 47465 5415 47521
rect 5471 47465 5557 47521
rect 5613 47465 5699 47521
rect 5755 47465 5841 47521
rect 5897 47465 5983 47521
rect 6039 47465 6125 47521
rect 6181 47465 6267 47521
rect 6323 47465 6409 47521
rect 6465 47465 6551 47521
rect 6607 47465 6693 47521
rect 6749 47465 6835 47521
rect 6891 47465 6977 47521
rect 7033 47465 7119 47521
rect 7175 47465 7261 47521
rect 7317 47465 7403 47521
rect 7459 47465 7545 47521
rect 7601 47465 7687 47521
rect 7743 47465 7829 47521
rect 7885 47465 7971 47521
rect 8027 47465 8113 47521
rect 8169 47465 8255 47521
rect 8311 47465 8397 47521
rect 8453 47465 8539 47521
rect 8595 47465 8681 47521
rect 8737 47465 8823 47521
rect 8879 47465 8965 47521
rect 9021 47465 9107 47521
rect 9163 47465 9249 47521
rect 9305 47465 9391 47521
rect 9447 47465 9533 47521
rect 9589 47465 9675 47521
rect 9731 47465 9817 47521
rect 9873 47465 9959 47521
rect 10015 47465 10101 47521
rect 10157 47465 10243 47521
rect 10299 47465 10385 47521
rect 10441 47465 10527 47521
rect 10583 47465 10669 47521
rect 10725 47465 10811 47521
rect 10867 47465 10953 47521
rect 11009 47465 11095 47521
rect 11151 47465 11237 47521
rect 11293 47465 11379 47521
rect 11435 47465 11521 47521
rect 11577 47465 11663 47521
rect 11719 47465 11805 47521
rect 11861 47465 11947 47521
rect 12003 47465 12089 47521
rect 12145 47465 12231 47521
rect 12287 47465 12373 47521
rect 12429 47465 12515 47521
rect 12571 47465 12657 47521
rect 12713 47465 12799 47521
rect 12855 47465 12941 47521
rect 12997 47465 13083 47521
rect 13139 47465 13225 47521
rect 13281 47465 13367 47521
rect 13423 47465 13509 47521
rect 13565 47465 13651 47521
rect 13707 47465 13793 47521
rect 13849 47465 13935 47521
rect 13991 47465 14077 47521
rect 14133 47465 14219 47521
rect 14275 47465 14361 47521
rect 14417 47465 14503 47521
rect 14559 47465 14645 47521
rect 14701 47465 14787 47521
rect 14843 47465 15000 47521
rect 0 47379 15000 47465
rect 0 47323 161 47379
rect 217 47323 303 47379
rect 359 47323 445 47379
rect 501 47323 587 47379
rect 643 47323 729 47379
rect 785 47323 871 47379
rect 927 47323 1013 47379
rect 1069 47323 1155 47379
rect 1211 47323 1297 47379
rect 1353 47323 1439 47379
rect 1495 47323 1581 47379
rect 1637 47323 1723 47379
rect 1779 47323 1865 47379
rect 1921 47323 2007 47379
rect 2063 47323 2149 47379
rect 2205 47323 2291 47379
rect 2347 47323 2433 47379
rect 2489 47323 2575 47379
rect 2631 47323 2717 47379
rect 2773 47323 2859 47379
rect 2915 47323 3001 47379
rect 3057 47323 3143 47379
rect 3199 47323 3285 47379
rect 3341 47323 3427 47379
rect 3483 47323 3569 47379
rect 3625 47323 3711 47379
rect 3767 47323 3853 47379
rect 3909 47323 3995 47379
rect 4051 47323 4137 47379
rect 4193 47323 4279 47379
rect 4335 47323 4421 47379
rect 4477 47323 4563 47379
rect 4619 47323 4705 47379
rect 4761 47323 4847 47379
rect 4903 47323 4989 47379
rect 5045 47323 5131 47379
rect 5187 47323 5273 47379
rect 5329 47323 5415 47379
rect 5471 47323 5557 47379
rect 5613 47323 5699 47379
rect 5755 47323 5841 47379
rect 5897 47323 5983 47379
rect 6039 47323 6125 47379
rect 6181 47323 6267 47379
rect 6323 47323 6409 47379
rect 6465 47323 6551 47379
rect 6607 47323 6693 47379
rect 6749 47323 6835 47379
rect 6891 47323 6977 47379
rect 7033 47323 7119 47379
rect 7175 47323 7261 47379
rect 7317 47323 7403 47379
rect 7459 47323 7545 47379
rect 7601 47323 7687 47379
rect 7743 47323 7829 47379
rect 7885 47323 7971 47379
rect 8027 47323 8113 47379
rect 8169 47323 8255 47379
rect 8311 47323 8397 47379
rect 8453 47323 8539 47379
rect 8595 47323 8681 47379
rect 8737 47323 8823 47379
rect 8879 47323 8965 47379
rect 9021 47323 9107 47379
rect 9163 47323 9249 47379
rect 9305 47323 9391 47379
rect 9447 47323 9533 47379
rect 9589 47323 9675 47379
rect 9731 47323 9817 47379
rect 9873 47323 9959 47379
rect 10015 47323 10101 47379
rect 10157 47323 10243 47379
rect 10299 47323 10385 47379
rect 10441 47323 10527 47379
rect 10583 47323 10669 47379
rect 10725 47323 10811 47379
rect 10867 47323 10953 47379
rect 11009 47323 11095 47379
rect 11151 47323 11237 47379
rect 11293 47323 11379 47379
rect 11435 47323 11521 47379
rect 11577 47323 11663 47379
rect 11719 47323 11805 47379
rect 11861 47323 11947 47379
rect 12003 47323 12089 47379
rect 12145 47323 12231 47379
rect 12287 47323 12373 47379
rect 12429 47323 12515 47379
rect 12571 47323 12657 47379
rect 12713 47323 12799 47379
rect 12855 47323 12941 47379
rect 12997 47323 13083 47379
rect 13139 47323 13225 47379
rect 13281 47323 13367 47379
rect 13423 47323 13509 47379
rect 13565 47323 13651 47379
rect 13707 47323 13793 47379
rect 13849 47323 13935 47379
rect 13991 47323 14077 47379
rect 14133 47323 14219 47379
rect 14275 47323 14361 47379
rect 14417 47323 14503 47379
rect 14559 47323 14645 47379
rect 14701 47323 14787 47379
rect 14843 47323 15000 47379
rect 0 47237 15000 47323
rect 0 47181 161 47237
rect 217 47181 303 47237
rect 359 47181 445 47237
rect 501 47181 587 47237
rect 643 47181 729 47237
rect 785 47181 871 47237
rect 927 47181 1013 47237
rect 1069 47181 1155 47237
rect 1211 47181 1297 47237
rect 1353 47181 1439 47237
rect 1495 47181 1581 47237
rect 1637 47181 1723 47237
rect 1779 47181 1865 47237
rect 1921 47181 2007 47237
rect 2063 47181 2149 47237
rect 2205 47181 2291 47237
rect 2347 47181 2433 47237
rect 2489 47181 2575 47237
rect 2631 47181 2717 47237
rect 2773 47181 2859 47237
rect 2915 47181 3001 47237
rect 3057 47181 3143 47237
rect 3199 47181 3285 47237
rect 3341 47181 3427 47237
rect 3483 47181 3569 47237
rect 3625 47181 3711 47237
rect 3767 47181 3853 47237
rect 3909 47181 3995 47237
rect 4051 47181 4137 47237
rect 4193 47181 4279 47237
rect 4335 47181 4421 47237
rect 4477 47181 4563 47237
rect 4619 47181 4705 47237
rect 4761 47181 4847 47237
rect 4903 47181 4989 47237
rect 5045 47181 5131 47237
rect 5187 47181 5273 47237
rect 5329 47181 5415 47237
rect 5471 47181 5557 47237
rect 5613 47181 5699 47237
rect 5755 47181 5841 47237
rect 5897 47181 5983 47237
rect 6039 47181 6125 47237
rect 6181 47181 6267 47237
rect 6323 47181 6409 47237
rect 6465 47181 6551 47237
rect 6607 47181 6693 47237
rect 6749 47181 6835 47237
rect 6891 47181 6977 47237
rect 7033 47181 7119 47237
rect 7175 47181 7261 47237
rect 7317 47181 7403 47237
rect 7459 47181 7545 47237
rect 7601 47181 7687 47237
rect 7743 47181 7829 47237
rect 7885 47181 7971 47237
rect 8027 47181 8113 47237
rect 8169 47181 8255 47237
rect 8311 47181 8397 47237
rect 8453 47181 8539 47237
rect 8595 47181 8681 47237
rect 8737 47181 8823 47237
rect 8879 47181 8965 47237
rect 9021 47181 9107 47237
rect 9163 47181 9249 47237
rect 9305 47181 9391 47237
rect 9447 47181 9533 47237
rect 9589 47181 9675 47237
rect 9731 47181 9817 47237
rect 9873 47181 9959 47237
rect 10015 47181 10101 47237
rect 10157 47181 10243 47237
rect 10299 47181 10385 47237
rect 10441 47181 10527 47237
rect 10583 47181 10669 47237
rect 10725 47181 10811 47237
rect 10867 47181 10953 47237
rect 11009 47181 11095 47237
rect 11151 47181 11237 47237
rect 11293 47181 11379 47237
rect 11435 47181 11521 47237
rect 11577 47181 11663 47237
rect 11719 47181 11805 47237
rect 11861 47181 11947 47237
rect 12003 47181 12089 47237
rect 12145 47181 12231 47237
rect 12287 47181 12373 47237
rect 12429 47181 12515 47237
rect 12571 47181 12657 47237
rect 12713 47181 12799 47237
rect 12855 47181 12941 47237
rect 12997 47181 13083 47237
rect 13139 47181 13225 47237
rect 13281 47181 13367 47237
rect 13423 47181 13509 47237
rect 13565 47181 13651 47237
rect 13707 47181 13793 47237
rect 13849 47181 13935 47237
rect 13991 47181 14077 47237
rect 14133 47181 14219 47237
rect 14275 47181 14361 47237
rect 14417 47181 14503 47237
rect 14559 47181 14645 47237
rect 14701 47181 14787 47237
rect 14843 47181 15000 47237
rect 0 47095 15000 47181
rect 0 47039 161 47095
rect 217 47039 303 47095
rect 359 47039 445 47095
rect 501 47039 587 47095
rect 643 47039 729 47095
rect 785 47039 871 47095
rect 927 47039 1013 47095
rect 1069 47039 1155 47095
rect 1211 47039 1297 47095
rect 1353 47039 1439 47095
rect 1495 47039 1581 47095
rect 1637 47039 1723 47095
rect 1779 47039 1865 47095
rect 1921 47039 2007 47095
rect 2063 47039 2149 47095
rect 2205 47039 2291 47095
rect 2347 47039 2433 47095
rect 2489 47039 2575 47095
rect 2631 47039 2717 47095
rect 2773 47039 2859 47095
rect 2915 47039 3001 47095
rect 3057 47039 3143 47095
rect 3199 47039 3285 47095
rect 3341 47039 3427 47095
rect 3483 47039 3569 47095
rect 3625 47039 3711 47095
rect 3767 47039 3853 47095
rect 3909 47039 3995 47095
rect 4051 47039 4137 47095
rect 4193 47039 4279 47095
rect 4335 47039 4421 47095
rect 4477 47039 4563 47095
rect 4619 47039 4705 47095
rect 4761 47039 4847 47095
rect 4903 47039 4989 47095
rect 5045 47039 5131 47095
rect 5187 47039 5273 47095
rect 5329 47039 5415 47095
rect 5471 47039 5557 47095
rect 5613 47039 5699 47095
rect 5755 47039 5841 47095
rect 5897 47039 5983 47095
rect 6039 47039 6125 47095
rect 6181 47039 6267 47095
rect 6323 47039 6409 47095
rect 6465 47039 6551 47095
rect 6607 47039 6693 47095
rect 6749 47039 6835 47095
rect 6891 47039 6977 47095
rect 7033 47039 7119 47095
rect 7175 47039 7261 47095
rect 7317 47039 7403 47095
rect 7459 47039 7545 47095
rect 7601 47039 7687 47095
rect 7743 47039 7829 47095
rect 7885 47039 7971 47095
rect 8027 47039 8113 47095
rect 8169 47039 8255 47095
rect 8311 47039 8397 47095
rect 8453 47039 8539 47095
rect 8595 47039 8681 47095
rect 8737 47039 8823 47095
rect 8879 47039 8965 47095
rect 9021 47039 9107 47095
rect 9163 47039 9249 47095
rect 9305 47039 9391 47095
rect 9447 47039 9533 47095
rect 9589 47039 9675 47095
rect 9731 47039 9817 47095
rect 9873 47039 9959 47095
rect 10015 47039 10101 47095
rect 10157 47039 10243 47095
rect 10299 47039 10385 47095
rect 10441 47039 10527 47095
rect 10583 47039 10669 47095
rect 10725 47039 10811 47095
rect 10867 47039 10953 47095
rect 11009 47039 11095 47095
rect 11151 47039 11237 47095
rect 11293 47039 11379 47095
rect 11435 47039 11521 47095
rect 11577 47039 11663 47095
rect 11719 47039 11805 47095
rect 11861 47039 11947 47095
rect 12003 47039 12089 47095
rect 12145 47039 12231 47095
rect 12287 47039 12373 47095
rect 12429 47039 12515 47095
rect 12571 47039 12657 47095
rect 12713 47039 12799 47095
rect 12855 47039 12941 47095
rect 12997 47039 13083 47095
rect 13139 47039 13225 47095
rect 13281 47039 13367 47095
rect 13423 47039 13509 47095
rect 13565 47039 13651 47095
rect 13707 47039 13793 47095
rect 13849 47039 13935 47095
rect 13991 47039 14077 47095
rect 14133 47039 14219 47095
rect 14275 47039 14361 47095
rect 14417 47039 14503 47095
rect 14559 47039 14645 47095
rect 14701 47039 14787 47095
rect 14843 47039 15000 47095
rect 0 46953 15000 47039
rect 0 46897 161 46953
rect 217 46897 303 46953
rect 359 46897 445 46953
rect 501 46897 587 46953
rect 643 46897 729 46953
rect 785 46897 871 46953
rect 927 46897 1013 46953
rect 1069 46897 1155 46953
rect 1211 46897 1297 46953
rect 1353 46897 1439 46953
rect 1495 46897 1581 46953
rect 1637 46897 1723 46953
rect 1779 46897 1865 46953
rect 1921 46897 2007 46953
rect 2063 46897 2149 46953
rect 2205 46897 2291 46953
rect 2347 46897 2433 46953
rect 2489 46897 2575 46953
rect 2631 46897 2717 46953
rect 2773 46897 2859 46953
rect 2915 46897 3001 46953
rect 3057 46897 3143 46953
rect 3199 46897 3285 46953
rect 3341 46897 3427 46953
rect 3483 46897 3569 46953
rect 3625 46897 3711 46953
rect 3767 46897 3853 46953
rect 3909 46897 3995 46953
rect 4051 46897 4137 46953
rect 4193 46897 4279 46953
rect 4335 46897 4421 46953
rect 4477 46897 4563 46953
rect 4619 46897 4705 46953
rect 4761 46897 4847 46953
rect 4903 46897 4989 46953
rect 5045 46897 5131 46953
rect 5187 46897 5273 46953
rect 5329 46897 5415 46953
rect 5471 46897 5557 46953
rect 5613 46897 5699 46953
rect 5755 46897 5841 46953
rect 5897 46897 5983 46953
rect 6039 46897 6125 46953
rect 6181 46897 6267 46953
rect 6323 46897 6409 46953
rect 6465 46897 6551 46953
rect 6607 46897 6693 46953
rect 6749 46897 6835 46953
rect 6891 46897 6977 46953
rect 7033 46897 7119 46953
rect 7175 46897 7261 46953
rect 7317 46897 7403 46953
rect 7459 46897 7545 46953
rect 7601 46897 7687 46953
rect 7743 46897 7829 46953
rect 7885 46897 7971 46953
rect 8027 46897 8113 46953
rect 8169 46897 8255 46953
rect 8311 46897 8397 46953
rect 8453 46897 8539 46953
rect 8595 46897 8681 46953
rect 8737 46897 8823 46953
rect 8879 46897 8965 46953
rect 9021 46897 9107 46953
rect 9163 46897 9249 46953
rect 9305 46897 9391 46953
rect 9447 46897 9533 46953
rect 9589 46897 9675 46953
rect 9731 46897 9817 46953
rect 9873 46897 9959 46953
rect 10015 46897 10101 46953
rect 10157 46897 10243 46953
rect 10299 46897 10385 46953
rect 10441 46897 10527 46953
rect 10583 46897 10669 46953
rect 10725 46897 10811 46953
rect 10867 46897 10953 46953
rect 11009 46897 11095 46953
rect 11151 46897 11237 46953
rect 11293 46897 11379 46953
rect 11435 46897 11521 46953
rect 11577 46897 11663 46953
rect 11719 46897 11805 46953
rect 11861 46897 11947 46953
rect 12003 46897 12089 46953
rect 12145 46897 12231 46953
rect 12287 46897 12373 46953
rect 12429 46897 12515 46953
rect 12571 46897 12657 46953
rect 12713 46897 12799 46953
rect 12855 46897 12941 46953
rect 12997 46897 13083 46953
rect 13139 46897 13225 46953
rect 13281 46897 13367 46953
rect 13423 46897 13509 46953
rect 13565 46897 13651 46953
rect 13707 46897 13793 46953
rect 13849 46897 13935 46953
rect 13991 46897 14077 46953
rect 14133 46897 14219 46953
rect 14275 46897 14361 46953
rect 14417 46897 14503 46953
rect 14559 46897 14645 46953
rect 14701 46897 14787 46953
rect 14843 46897 15000 46953
rect 0 46811 15000 46897
rect 0 46755 161 46811
rect 217 46755 303 46811
rect 359 46755 445 46811
rect 501 46755 587 46811
rect 643 46755 729 46811
rect 785 46755 871 46811
rect 927 46755 1013 46811
rect 1069 46755 1155 46811
rect 1211 46755 1297 46811
rect 1353 46755 1439 46811
rect 1495 46755 1581 46811
rect 1637 46755 1723 46811
rect 1779 46755 1865 46811
rect 1921 46755 2007 46811
rect 2063 46755 2149 46811
rect 2205 46755 2291 46811
rect 2347 46755 2433 46811
rect 2489 46755 2575 46811
rect 2631 46755 2717 46811
rect 2773 46755 2859 46811
rect 2915 46755 3001 46811
rect 3057 46755 3143 46811
rect 3199 46755 3285 46811
rect 3341 46755 3427 46811
rect 3483 46755 3569 46811
rect 3625 46755 3711 46811
rect 3767 46755 3853 46811
rect 3909 46755 3995 46811
rect 4051 46755 4137 46811
rect 4193 46755 4279 46811
rect 4335 46755 4421 46811
rect 4477 46755 4563 46811
rect 4619 46755 4705 46811
rect 4761 46755 4847 46811
rect 4903 46755 4989 46811
rect 5045 46755 5131 46811
rect 5187 46755 5273 46811
rect 5329 46755 5415 46811
rect 5471 46755 5557 46811
rect 5613 46755 5699 46811
rect 5755 46755 5841 46811
rect 5897 46755 5983 46811
rect 6039 46755 6125 46811
rect 6181 46755 6267 46811
rect 6323 46755 6409 46811
rect 6465 46755 6551 46811
rect 6607 46755 6693 46811
rect 6749 46755 6835 46811
rect 6891 46755 6977 46811
rect 7033 46755 7119 46811
rect 7175 46755 7261 46811
rect 7317 46755 7403 46811
rect 7459 46755 7545 46811
rect 7601 46755 7687 46811
rect 7743 46755 7829 46811
rect 7885 46755 7971 46811
rect 8027 46755 8113 46811
rect 8169 46755 8255 46811
rect 8311 46755 8397 46811
rect 8453 46755 8539 46811
rect 8595 46755 8681 46811
rect 8737 46755 8823 46811
rect 8879 46755 8965 46811
rect 9021 46755 9107 46811
rect 9163 46755 9249 46811
rect 9305 46755 9391 46811
rect 9447 46755 9533 46811
rect 9589 46755 9675 46811
rect 9731 46755 9817 46811
rect 9873 46755 9959 46811
rect 10015 46755 10101 46811
rect 10157 46755 10243 46811
rect 10299 46755 10385 46811
rect 10441 46755 10527 46811
rect 10583 46755 10669 46811
rect 10725 46755 10811 46811
rect 10867 46755 10953 46811
rect 11009 46755 11095 46811
rect 11151 46755 11237 46811
rect 11293 46755 11379 46811
rect 11435 46755 11521 46811
rect 11577 46755 11663 46811
rect 11719 46755 11805 46811
rect 11861 46755 11947 46811
rect 12003 46755 12089 46811
rect 12145 46755 12231 46811
rect 12287 46755 12373 46811
rect 12429 46755 12515 46811
rect 12571 46755 12657 46811
rect 12713 46755 12799 46811
rect 12855 46755 12941 46811
rect 12997 46755 13083 46811
rect 13139 46755 13225 46811
rect 13281 46755 13367 46811
rect 13423 46755 13509 46811
rect 13565 46755 13651 46811
rect 13707 46755 13793 46811
rect 13849 46755 13935 46811
rect 13991 46755 14077 46811
rect 14133 46755 14219 46811
rect 14275 46755 14361 46811
rect 14417 46755 14503 46811
rect 14559 46755 14645 46811
rect 14701 46755 14787 46811
rect 14843 46755 15000 46811
rect 0 46669 15000 46755
rect 0 46613 161 46669
rect 217 46613 303 46669
rect 359 46613 445 46669
rect 501 46613 587 46669
rect 643 46613 729 46669
rect 785 46613 871 46669
rect 927 46613 1013 46669
rect 1069 46613 1155 46669
rect 1211 46613 1297 46669
rect 1353 46613 1439 46669
rect 1495 46613 1581 46669
rect 1637 46613 1723 46669
rect 1779 46613 1865 46669
rect 1921 46613 2007 46669
rect 2063 46613 2149 46669
rect 2205 46613 2291 46669
rect 2347 46613 2433 46669
rect 2489 46613 2575 46669
rect 2631 46613 2717 46669
rect 2773 46613 2859 46669
rect 2915 46613 3001 46669
rect 3057 46613 3143 46669
rect 3199 46613 3285 46669
rect 3341 46613 3427 46669
rect 3483 46613 3569 46669
rect 3625 46613 3711 46669
rect 3767 46613 3853 46669
rect 3909 46613 3995 46669
rect 4051 46613 4137 46669
rect 4193 46613 4279 46669
rect 4335 46613 4421 46669
rect 4477 46613 4563 46669
rect 4619 46613 4705 46669
rect 4761 46613 4847 46669
rect 4903 46613 4989 46669
rect 5045 46613 5131 46669
rect 5187 46613 5273 46669
rect 5329 46613 5415 46669
rect 5471 46613 5557 46669
rect 5613 46613 5699 46669
rect 5755 46613 5841 46669
rect 5897 46613 5983 46669
rect 6039 46613 6125 46669
rect 6181 46613 6267 46669
rect 6323 46613 6409 46669
rect 6465 46613 6551 46669
rect 6607 46613 6693 46669
rect 6749 46613 6835 46669
rect 6891 46613 6977 46669
rect 7033 46613 7119 46669
rect 7175 46613 7261 46669
rect 7317 46613 7403 46669
rect 7459 46613 7545 46669
rect 7601 46613 7687 46669
rect 7743 46613 7829 46669
rect 7885 46613 7971 46669
rect 8027 46613 8113 46669
rect 8169 46613 8255 46669
rect 8311 46613 8397 46669
rect 8453 46613 8539 46669
rect 8595 46613 8681 46669
rect 8737 46613 8823 46669
rect 8879 46613 8965 46669
rect 9021 46613 9107 46669
rect 9163 46613 9249 46669
rect 9305 46613 9391 46669
rect 9447 46613 9533 46669
rect 9589 46613 9675 46669
rect 9731 46613 9817 46669
rect 9873 46613 9959 46669
rect 10015 46613 10101 46669
rect 10157 46613 10243 46669
rect 10299 46613 10385 46669
rect 10441 46613 10527 46669
rect 10583 46613 10669 46669
rect 10725 46613 10811 46669
rect 10867 46613 10953 46669
rect 11009 46613 11095 46669
rect 11151 46613 11237 46669
rect 11293 46613 11379 46669
rect 11435 46613 11521 46669
rect 11577 46613 11663 46669
rect 11719 46613 11805 46669
rect 11861 46613 11947 46669
rect 12003 46613 12089 46669
rect 12145 46613 12231 46669
rect 12287 46613 12373 46669
rect 12429 46613 12515 46669
rect 12571 46613 12657 46669
rect 12713 46613 12799 46669
rect 12855 46613 12941 46669
rect 12997 46613 13083 46669
rect 13139 46613 13225 46669
rect 13281 46613 13367 46669
rect 13423 46613 13509 46669
rect 13565 46613 13651 46669
rect 13707 46613 13793 46669
rect 13849 46613 13935 46669
rect 13991 46613 14077 46669
rect 14133 46613 14219 46669
rect 14275 46613 14361 46669
rect 14417 46613 14503 46669
rect 14559 46613 14645 46669
rect 14701 46613 14787 46669
rect 14843 46613 15000 46669
rect 0 46527 15000 46613
rect 0 46471 161 46527
rect 217 46471 303 46527
rect 359 46471 445 46527
rect 501 46471 587 46527
rect 643 46471 729 46527
rect 785 46471 871 46527
rect 927 46471 1013 46527
rect 1069 46471 1155 46527
rect 1211 46471 1297 46527
rect 1353 46471 1439 46527
rect 1495 46471 1581 46527
rect 1637 46471 1723 46527
rect 1779 46471 1865 46527
rect 1921 46471 2007 46527
rect 2063 46471 2149 46527
rect 2205 46471 2291 46527
rect 2347 46471 2433 46527
rect 2489 46471 2575 46527
rect 2631 46471 2717 46527
rect 2773 46471 2859 46527
rect 2915 46471 3001 46527
rect 3057 46471 3143 46527
rect 3199 46471 3285 46527
rect 3341 46471 3427 46527
rect 3483 46471 3569 46527
rect 3625 46471 3711 46527
rect 3767 46471 3853 46527
rect 3909 46471 3995 46527
rect 4051 46471 4137 46527
rect 4193 46471 4279 46527
rect 4335 46471 4421 46527
rect 4477 46471 4563 46527
rect 4619 46471 4705 46527
rect 4761 46471 4847 46527
rect 4903 46471 4989 46527
rect 5045 46471 5131 46527
rect 5187 46471 5273 46527
rect 5329 46471 5415 46527
rect 5471 46471 5557 46527
rect 5613 46471 5699 46527
rect 5755 46471 5841 46527
rect 5897 46471 5983 46527
rect 6039 46471 6125 46527
rect 6181 46471 6267 46527
rect 6323 46471 6409 46527
rect 6465 46471 6551 46527
rect 6607 46471 6693 46527
rect 6749 46471 6835 46527
rect 6891 46471 6977 46527
rect 7033 46471 7119 46527
rect 7175 46471 7261 46527
rect 7317 46471 7403 46527
rect 7459 46471 7545 46527
rect 7601 46471 7687 46527
rect 7743 46471 7829 46527
rect 7885 46471 7971 46527
rect 8027 46471 8113 46527
rect 8169 46471 8255 46527
rect 8311 46471 8397 46527
rect 8453 46471 8539 46527
rect 8595 46471 8681 46527
rect 8737 46471 8823 46527
rect 8879 46471 8965 46527
rect 9021 46471 9107 46527
rect 9163 46471 9249 46527
rect 9305 46471 9391 46527
rect 9447 46471 9533 46527
rect 9589 46471 9675 46527
rect 9731 46471 9817 46527
rect 9873 46471 9959 46527
rect 10015 46471 10101 46527
rect 10157 46471 10243 46527
rect 10299 46471 10385 46527
rect 10441 46471 10527 46527
rect 10583 46471 10669 46527
rect 10725 46471 10811 46527
rect 10867 46471 10953 46527
rect 11009 46471 11095 46527
rect 11151 46471 11237 46527
rect 11293 46471 11379 46527
rect 11435 46471 11521 46527
rect 11577 46471 11663 46527
rect 11719 46471 11805 46527
rect 11861 46471 11947 46527
rect 12003 46471 12089 46527
rect 12145 46471 12231 46527
rect 12287 46471 12373 46527
rect 12429 46471 12515 46527
rect 12571 46471 12657 46527
rect 12713 46471 12799 46527
rect 12855 46471 12941 46527
rect 12997 46471 13083 46527
rect 13139 46471 13225 46527
rect 13281 46471 13367 46527
rect 13423 46471 13509 46527
rect 13565 46471 13651 46527
rect 13707 46471 13793 46527
rect 13849 46471 13935 46527
rect 13991 46471 14077 46527
rect 14133 46471 14219 46527
rect 14275 46471 14361 46527
rect 14417 46471 14503 46527
rect 14559 46471 14645 46527
rect 14701 46471 14787 46527
rect 14843 46471 15000 46527
rect 0 46385 15000 46471
rect 0 46329 161 46385
rect 217 46329 303 46385
rect 359 46329 445 46385
rect 501 46329 587 46385
rect 643 46329 729 46385
rect 785 46329 871 46385
rect 927 46329 1013 46385
rect 1069 46329 1155 46385
rect 1211 46329 1297 46385
rect 1353 46329 1439 46385
rect 1495 46329 1581 46385
rect 1637 46329 1723 46385
rect 1779 46329 1865 46385
rect 1921 46329 2007 46385
rect 2063 46329 2149 46385
rect 2205 46329 2291 46385
rect 2347 46329 2433 46385
rect 2489 46329 2575 46385
rect 2631 46329 2717 46385
rect 2773 46329 2859 46385
rect 2915 46329 3001 46385
rect 3057 46329 3143 46385
rect 3199 46329 3285 46385
rect 3341 46329 3427 46385
rect 3483 46329 3569 46385
rect 3625 46329 3711 46385
rect 3767 46329 3853 46385
rect 3909 46329 3995 46385
rect 4051 46329 4137 46385
rect 4193 46329 4279 46385
rect 4335 46329 4421 46385
rect 4477 46329 4563 46385
rect 4619 46329 4705 46385
rect 4761 46329 4847 46385
rect 4903 46329 4989 46385
rect 5045 46329 5131 46385
rect 5187 46329 5273 46385
rect 5329 46329 5415 46385
rect 5471 46329 5557 46385
rect 5613 46329 5699 46385
rect 5755 46329 5841 46385
rect 5897 46329 5983 46385
rect 6039 46329 6125 46385
rect 6181 46329 6267 46385
rect 6323 46329 6409 46385
rect 6465 46329 6551 46385
rect 6607 46329 6693 46385
rect 6749 46329 6835 46385
rect 6891 46329 6977 46385
rect 7033 46329 7119 46385
rect 7175 46329 7261 46385
rect 7317 46329 7403 46385
rect 7459 46329 7545 46385
rect 7601 46329 7687 46385
rect 7743 46329 7829 46385
rect 7885 46329 7971 46385
rect 8027 46329 8113 46385
rect 8169 46329 8255 46385
rect 8311 46329 8397 46385
rect 8453 46329 8539 46385
rect 8595 46329 8681 46385
rect 8737 46329 8823 46385
rect 8879 46329 8965 46385
rect 9021 46329 9107 46385
rect 9163 46329 9249 46385
rect 9305 46329 9391 46385
rect 9447 46329 9533 46385
rect 9589 46329 9675 46385
rect 9731 46329 9817 46385
rect 9873 46329 9959 46385
rect 10015 46329 10101 46385
rect 10157 46329 10243 46385
rect 10299 46329 10385 46385
rect 10441 46329 10527 46385
rect 10583 46329 10669 46385
rect 10725 46329 10811 46385
rect 10867 46329 10953 46385
rect 11009 46329 11095 46385
rect 11151 46329 11237 46385
rect 11293 46329 11379 46385
rect 11435 46329 11521 46385
rect 11577 46329 11663 46385
rect 11719 46329 11805 46385
rect 11861 46329 11947 46385
rect 12003 46329 12089 46385
rect 12145 46329 12231 46385
rect 12287 46329 12373 46385
rect 12429 46329 12515 46385
rect 12571 46329 12657 46385
rect 12713 46329 12799 46385
rect 12855 46329 12941 46385
rect 12997 46329 13083 46385
rect 13139 46329 13225 46385
rect 13281 46329 13367 46385
rect 13423 46329 13509 46385
rect 13565 46329 13651 46385
rect 13707 46329 13793 46385
rect 13849 46329 13935 46385
rect 13991 46329 14077 46385
rect 14133 46329 14219 46385
rect 14275 46329 14361 46385
rect 14417 46329 14503 46385
rect 14559 46329 14645 46385
rect 14701 46329 14787 46385
rect 14843 46329 15000 46385
rect 0 46243 15000 46329
rect 0 46187 161 46243
rect 217 46187 303 46243
rect 359 46187 445 46243
rect 501 46187 587 46243
rect 643 46187 729 46243
rect 785 46187 871 46243
rect 927 46187 1013 46243
rect 1069 46187 1155 46243
rect 1211 46187 1297 46243
rect 1353 46187 1439 46243
rect 1495 46187 1581 46243
rect 1637 46187 1723 46243
rect 1779 46187 1865 46243
rect 1921 46187 2007 46243
rect 2063 46187 2149 46243
rect 2205 46187 2291 46243
rect 2347 46187 2433 46243
rect 2489 46187 2575 46243
rect 2631 46187 2717 46243
rect 2773 46187 2859 46243
rect 2915 46187 3001 46243
rect 3057 46187 3143 46243
rect 3199 46187 3285 46243
rect 3341 46187 3427 46243
rect 3483 46187 3569 46243
rect 3625 46187 3711 46243
rect 3767 46187 3853 46243
rect 3909 46187 3995 46243
rect 4051 46187 4137 46243
rect 4193 46187 4279 46243
rect 4335 46187 4421 46243
rect 4477 46187 4563 46243
rect 4619 46187 4705 46243
rect 4761 46187 4847 46243
rect 4903 46187 4989 46243
rect 5045 46187 5131 46243
rect 5187 46187 5273 46243
rect 5329 46187 5415 46243
rect 5471 46187 5557 46243
rect 5613 46187 5699 46243
rect 5755 46187 5841 46243
rect 5897 46187 5983 46243
rect 6039 46187 6125 46243
rect 6181 46187 6267 46243
rect 6323 46187 6409 46243
rect 6465 46187 6551 46243
rect 6607 46187 6693 46243
rect 6749 46187 6835 46243
rect 6891 46187 6977 46243
rect 7033 46187 7119 46243
rect 7175 46187 7261 46243
rect 7317 46187 7403 46243
rect 7459 46187 7545 46243
rect 7601 46187 7687 46243
rect 7743 46187 7829 46243
rect 7885 46187 7971 46243
rect 8027 46187 8113 46243
rect 8169 46187 8255 46243
rect 8311 46187 8397 46243
rect 8453 46187 8539 46243
rect 8595 46187 8681 46243
rect 8737 46187 8823 46243
rect 8879 46187 8965 46243
rect 9021 46187 9107 46243
rect 9163 46187 9249 46243
rect 9305 46187 9391 46243
rect 9447 46187 9533 46243
rect 9589 46187 9675 46243
rect 9731 46187 9817 46243
rect 9873 46187 9959 46243
rect 10015 46187 10101 46243
rect 10157 46187 10243 46243
rect 10299 46187 10385 46243
rect 10441 46187 10527 46243
rect 10583 46187 10669 46243
rect 10725 46187 10811 46243
rect 10867 46187 10953 46243
rect 11009 46187 11095 46243
rect 11151 46187 11237 46243
rect 11293 46187 11379 46243
rect 11435 46187 11521 46243
rect 11577 46187 11663 46243
rect 11719 46187 11805 46243
rect 11861 46187 11947 46243
rect 12003 46187 12089 46243
rect 12145 46187 12231 46243
rect 12287 46187 12373 46243
rect 12429 46187 12515 46243
rect 12571 46187 12657 46243
rect 12713 46187 12799 46243
rect 12855 46187 12941 46243
rect 12997 46187 13083 46243
rect 13139 46187 13225 46243
rect 13281 46187 13367 46243
rect 13423 46187 13509 46243
rect 13565 46187 13651 46243
rect 13707 46187 13793 46243
rect 13849 46187 13935 46243
rect 13991 46187 14077 46243
rect 14133 46187 14219 46243
rect 14275 46187 14361 46243
rect 14417 46187 14503 46243
rect 14559 46187 14645 46243
rect 14701 46187 14787 46243
rect 14843 46187 15000 46243
rect 0 46101 15000 46187
rect 0 46045 161 46101
rect 217 46045 303 46101
rect 359 46045 445 46101
rect 501 46045 587 46101
rect 643 46045 729 46101
rect 785 46045 871 46101
rect 927 46045 1013 46101
rect 1069 46045 1155 46101
rect 1211 46045 1297 46101
rect 1353 46045 1439 46101
rect 1495 46045 1581 46101
rect 1637 46045 1723 46101
rect 1779 46045 1865 46101
rect 1921 46045 2007 46101
rect 2063 46045 2149 46101
rect 2205 46045 2291 46101
rect 2347 46045 2433 46101
rect 2489 46045 2575 46101
rect 2631 46045 2717 46101
rect 2773 46045 2859 46101
rect 2915 46045 3001 46101
rect 3057 46045 3143 46101
rect 3199 46045 3285 46101
rect 3341 46045 3427 46101
rect 3483 46045 3569 46101
rect 3625 46045 3711 46101
rect 3767 46045 3853 46101
rect 3909 46045 3995 46101
rect 4051 46045 4137 46101
rect 4193 46045 4279 46101
rect 4335 46045 4421 46101
rect 4477 46045 4563 46101
rect 4619 46045 4705 46101
rect 4761 46045 4847 46101
rect 4903 46045 4989 46101
rect 5045 46045 5131 46101
rect 5187 46045 5273 46101
rect 5329 46045 5415 46101
rect 5471 46045 5557 46101
rect 5613 46045 5699 46101
rect 5755 46045 5841 46101
rect 5897 46045 5983 46101
rect 6039 46045 6125 46101
rect 6181 46045 6267 46101
rect 6323 46045 6409 46101
rect 6465 46045 6551 46101
rect 6607 46045 6693 46101
rect 6749 46045 6835 46101
rect 6891 46045 6977 46101
rect 7033 46045 7119 46101
rect 7175 46045 7261 46101
rect 7317 46045 7403 46101
rect 7459 46045 7545 46101
rect 7601 46045 7687 46101
rect 7743 46045 7829 46101
rect 7885 46045 7971 46101
rect 8027 46045 8113 46101
rect 8169 46045 8255 46101
rect 8311 46045 8397 46101
rect 8453 46045 8539 46101
rect 8595 46045 8681 46101
rect 8737 46045 8823 46101
rect 8879 46045 8965 46101
rect 9021 46045 9107 46101
rect 9163 46045 9249 46101
rect 9305 46045 9391 46101
rect 9447 46045 9533 46101
rect 9589 46045 9675 46101
rect 9731 46045 9817 46101
rect 9873 46045 9959 46101
rect 10015 46045 10101 46101
rect 10157 46045 10243 46101
rect 10299 46045 10385 46101
rect 10441 46045 10527 46101
rect 10583 46045 10669 46101
rect 10725 46045 10811 46101
rect 10867 46045 10953 46101
rect 11009 46045 11095 46101
rect 11151 46045 11237 46101
rect 11293 46045 11379 46101
rect 11435 46045 11521 46101
rect 11577 46045 11663 46101
rect 11719 46045 11805 46101
rect 11861 46045 11947 46101
rect 12003 46045 12089 46101
rect 12145 46045 12231 46101
rect 12287 46045 12373 46101
rect 12429 46045 12515 46101
rect 12571 46045 12657 46101
rect 12713 46045 12799 46101
rect 12855 46045 12941 46101
rect 12997 46045 13083 46101
rect 13139 46045 13225 46101
rect 13281 46045 13367 46101
rect 13423 46045 13509 46101
rect 13565 46045 13651 46101
rect 13707 46045 13793 46101
rect 13849 46045 13935 46101
rect 13991 46045 14077 46101
rect 14133 46045 14219 46101
rect 14275 46045 14361 46101
rect 14417 46045 14503 46101
rect 14559 46045 14645 46101
rect 14701 46045 14787 46101
rect 14843 46045 15000 46101
rect 0 46000 15000 46045
rect 0 45741 15000 45800
rect 0 45685 161 45741
rect 217 45685 303 45741
rect 359 45685 445 45741
rect 501 45685 587 45741
rect 643 45685 729 45741
rect 785 45685 871 45741
rect 927 45685 1013 45741
rect 1069 45685 1155 45741
rect 1211 45685 1297 45741
rect 1353 45685 1439 45741
rect 1495 45685 1581 45741
rect 1637 45685 1723 45741
rect 1779 45685 1865 45741
rect 1921 45685 2007 45741
rect 2063 45685 2149 45741
rect 2205 45685 2291 45741
rect 2347 45685 2433 45741
rect 2489 45685 2575 45741
rect 2631 45685 2717 45741
rect 2773 45685 2859 45741
rect 2915 45685 3001 45741
rect 3057 45685 3143 45741
rect 3199 45685 3285 45741
rect 3341 45685 3427 45741
rect 3483 45685 3569 45741
rect 3625 45685 3711 45741
rect 3767 45685 3853 45741
rect 3909 45685 3995 45741
rect 4051 45685 4137 45741
rect 4193 45685 4279 45741
rect 4335 45685 4421 45741
rect 4477 45685 4563 45741
rect 4619 45685 4705 45741
rect 4761 45685 4847 45741
rect 4903 45685 4989 45741
rect 5045 45685 5131 45741
rect 5187 45685 5273 45741
rect 5329 45685 5415 45741
rect 5471 45685 5557 45741
rect 5613 45685 5699 45741
rect 5755 45685 5841 45741
rect 5897 45685 5983 45741
rect 6039 45685 6125 45741
rect 6181 45685 6267 45741
rect 6323 45685 6409 45741
rect 6465 45685 6551 45741
rect 6607 45685 6693 45741
rect 6749 45685 6835 45741
rect 6891 45685 6977 45741
rect 7033 45685 7119 45741
rect 7175 45685 7261 45741
rect 7317 45685 7403 45741
rect 7459 45685 7545 45741
rect 7601 45685 7687 45741
rect 7743 45685 7829 45741
rect 7885 45685 7971 45741
rect 8027 45685 8113 45741
rect 8169 45685 8255 45741
rect 8311 45685 8397 45741
rect 8453 45685 8539 45741
rect 8595 45685 8681 45741
rect 8737 45685 8823 45741
rect 8879 45685 8965 45741
rect 9021 45685 9107 45741
rect 9163 45685 9249 45741
rect 9305 45685 9391 45741
rect 9447 45685 9533 45741
rect 9589 45685 9675 45741
rect 9731 45685 9817 45741
rect 9873 45685 9959 45741
rect 10015 45685 10101 45741
rect 10157 45685 10243 45741
rect 10299 45685 10385 45741
rect 10441 45685 10527 45741
rect 10583 45685 10669 45741
rect 10725 45685 10811 45741
rect 10867 45685 10953 45741
rect 11009 45685 11095 45741
rect 11151 45685 11237 45741
rect 11293 45685 11379 45741
rect 11435 45685 11521 45741
rect 11577 45685 11663 45741
rect 11719 45685 11805 45741
rect 11861 45685 11947 45741
rect 12003 45685 12089 45741
rect 12145 45685 12231 45741
rect 12287 45685 12373 45741
rect 12429 45685 12515 45741
rect 12571 45685 12657 45741
rect 12713 45685 12799 45741
rect 12855 45685 12941 45741
rect 12997 45685 13083 45741
rect 13139 45685 13225 45741
rect 13281 45685 13367 45741
rect 13423 45685 13509 45741
rect 13565 45685 13651 45741
rect 13707 45685 13793 45741
rect 13849 45685 13935 45741
rect 13991 45685 14077 45741
rect 14133 45685 14219 45741
rect 14275 45685 14361 45741
rect 14417 45685 14503 45741
rect 14559 45685 14645 45741
rect 14701 45685 14787 45741
rect 14843 45685 15000 45741
rect 0 45599 15000 45685
rect 0 45543 161 45599
rect 217 45543 303 45599
rect 359 45543 445 45599
rect 501 45543 587 45599
rect 643 45543 729 45599
rect 785 45543 871 45599
rect 927 45543 1013 45599
rect 1069 45543 1155 45599
rect 1211 45543 1297 45599
rect 1353 45543 1439 45599
rect 1495 45543 1581 45599
rect 1637 45543 1723 45599
rect 1779 45543 1865 45599
rect 1921 45543 2007 45599
rect 2063 45543 2149 45599
rect 2205 45543 2291 45599
rect 2347 45543 2433 45599
rect 2489 45543 2575 45599
rect 2631 45543 2717 45599
rect 2773 45543 2859 45599
rect 2915 45543 3001 45599
rect 3057 45543 3143 45599
rect 3199 45543 3285 45599
rect 3341 45543 3427 45599
rect 3483 45543 3569 45599
rect 3625 45543 3711 45599
rect 3767 45543 3853 45599
rect 3909 45543 3995 45599
rect 4051 45543 4137 45599
rect 4193 45543 4279 45599
rect 4335 45543 4421 45599
rect 4477 45543 4563 45599
rect 4619 45543 4705 45599
rect 4761 45543 4847 45599
rect 4903 45543 4989 45599
rect 5045 45543 5131 45599
rect 5187 45543 5273 45599
rect 5329 45543 5415 45599
rect 5471 45543 5557 45599
rect 5613 45543 5699 45599
rect 5755 45543 5841 45599
rect 5897 45543 5983 45599
rect 6039 45543 6125 45599
rect 6181 45543 6267 45599
rect 6323 45543 6409 45599
rect 6465 45543 6551 45599
rect 6607 45543 6693 45599
rect 6749 45543 6835 45599
rect 6891 45543 6977 45599
rect 7033 45543 7119 45599
rect 7175 45543 7261 45599
rect 7317 45543 7403 45599
rect 7459 45543 7545 45599
rect 7601 45543 7687 45599
rect 7743 45543 7829 45599
rect 7885 45543 7971 45599
rect 8027 45543 8113 45599
rect 8169 45543 8255 45599
rect 8311 45543 8397 45599
rect 8453 45543 8539 45599
rect 8595 45543 8681 45599
rect 8737 45543 8823 45599
rect 8879 45543 8965 45599
rect 9021 45543 9107 45599
rect 9163 45543 9249 45599
rect 9305 45543 9391 45599
rect 9447 45543 9533 45599
rect 9589 45543 9675 45599
rect 9731 45543 9817 45599
rect 9873 45543 9959 45599
rect 10015 45543 10101 45599
rect 10157 45543 10243 45599
rect 10299 45543 10385 45599
rect 10441 45543 10527 45599
rect 10583 45543 10669 45599
rect 10725 45543 10811 45599
rect 10867 45543 10953 45599
rect 11009 45543 11095 45599
rect 11151 45543 11237 45599
rect 11293 45543 11379 45599
rect 11435 45543 11521 45599
rect 11577 45543 11663 45599
rect 11719 45543 11805 45599
rect 11861 45543 11947 45599
rect 12003 45543 12089 45599
rect 12145 45543 12231 45599
rect 12287 45543 12373 45599
rect 12429 45543 12515 45599
rect 12571 45543 12657 45599
rect 12713 45543 12799 45599
rect 12855 45543 12941 45599
rect 12997 45543 13083 45599
rect 13139 45543 13225 45599
rect 13281 45543 13367 45599
rect 13423 45543 13509 45599
rect 13565 45543 13651 45599
rect 13707 45543 13793 45599
rect 13849 45543 13935 45599
rect 13991 45543 14077 45599
rect 14133 45543 14219 45599
rect 14275 45543 14361 45599
rect 14417 45543 14503 45599
rect 14559 45543 14645 45599
rect 14701 45543 14787 45599
rect 14843 45543 15000 45599
rect 0 45457 15000 45543
rect 0 45401 161 45457
rect 217 45401 303 45457
rect 359 45401 445 45457
rect 501 45401 587 45457
rect 643 45401 729 45457
rect 785 45401 871 45457
rect 927 45401 1013 45457
rect 1069 45401 1155 45457
rect 1211 45401 1297 45457
rect 1353 45401 1439 45457
rect 1495 45401 1581 45457
rect 1637 45401 1723 45457
rect 1779 45401 1865 45457
rect 1921 45401 2007 45457
rect 2063 45401 2149 45457
rect 2205 45401 2291 45457
rect 2347 45401 2433 45457
rect 2489 45401 2575 45457
rect 2631 45401 2717 45457
rect 2773 45401 2859 45457
rect 2915 45401 3001 45457
rect 3057 45401 3143 45457
rect 3199 45401 3285 45457
rect 3341 45401 3427 45457
rect 3483 45401 3569 45457
rect 3625 45401 3711 45457
rect 3767 45401 3853 45457
rect 3909 45401 3995 45457
rect 4051 45401 4137 45457
rect 4193 45401 4279 45457
rect 4335 45401 4421 45457
rect 4477 45401 4563 45457
rect 4619 45401 4705 45457
rect 4761 45401 4847 45457
rect 4903 45401 4989 45457
rect 5045 45401 5131 45457
rect 5187 45401 5273 45457
rect 5329 45401 5415 45457
rect 5471 45401 5557 45457
rect 5613 45401 5699 45457
rect 5755 45401 5841 45457
rect 5897 45401 5983 45457
rect 6039 45401 6125 45457
rect 6181 45401 6267 45457
rect 6323 45401 6409 45457
rect 6465 45401 6551 45457
rect 6607 45401 6693 45457
rect 6749 45401 6835 45457
rect 6891 45401 6977 45457
rect 7033 45401 7119 45457
rect 7175 45401 7261 45457
rect 7317 45401 7403 45457
rect 7459 45401 7545 45457
rect 7601 45401 7687 45457
rect 7743 45401 7829 45457
rect 7885 45401 7971 45457
rect 8027 45401 8113 45457
rect 8169 45401 8255 45457
rect 8311 45401 8397 45457
rect 8453 45401 8539 45457
rect 8595 45401 8681 45457
rect 8737 45401 8823 45457
rect 8879 45401 8965 45457
rect 9021 45401 9107 45457
rect 9163 45401 9249 45457
rect 9305 45401 9391 45457
rect 9447 45401 9533 45457
rect 9589 45401 9675 45457
rect 9731 45401 9817 45457
rect 9873 45401 9959 45457
rect 10015 45401 10101 45457
rect 10157 45401 10243 45457
rect 10299 45401 10385 45457
rect 10441 45401 10527 45457
rect 10583 45401 10669 45457
rect 10725 45401 10811 45457
rect 10867 45401 10953 45457
rect 11009 45401 11095 45457
rect 11151 45401 11237 45457
rect 11293 45401 11379 45457
rect 11435 45401 11521 45457
rect 11577 45401 11663 45457
rect 11719 45401 11805 45457
rect 11861 45401 11947 45457
rect 12003 45401 12089 45457
rect 12145 45401 12231 45457
rect 12287 45401 12373 45457
rect 12429 45401 12515 45457
rect 12571 45401 12657 45457
rect 12713 45401 12799 45457
rect 12855 45401 12941 45457
rect 12997 45401 13083 45457
rect 13139 45401 13225 45457
rect 13281 45401 13367 45457
rect 13423 45401 13509 45457
rect 13565 45401 13651 45457
rect 13707 45401 13793 45457
rect 13849 45401 13935 45457
rect 13991 45401 14077 45457
rect 14133 45401 14219 45457
rect 14275 45401 14361 45457
rect 14417 45401 14503 45457
rect 14559 45401 14645 45457
rect 14701 45401 14787 45457
rect 14843 45401 15000 45457
rect 0 45315 15000 45401
rect 0 45259 161 45315
rect 217 45259 303 45315
rect 359 45259 445 45315
rect 501 45259 587 45315
rect 643 45259 729 45315
rect 785 45259 871 45315
rect 927 45259 1013 45315
rect 1069 45259 1155 45315
rect 1211 45259 1297 45315
rect 1353 45259 1439 45315
rect 1495 45259 1581 45315
rect 1637 45259 1723 45315
rect 1779 45259 1865 45315
rect 1921 45259 2007 45315
rect 2063 45259 2149 45315
rect 2205 45259 2291 45315
rect 2347 45259 2433 45315
rect 2489 45259 2575 45315
rect 2631 45259 2717 45315
rect 2773 45259 2859 45315
rect 2915 45259 3001 45315
rect 3057 45259 3143 45315
rect 3199 45259 3285 45315
rect 3341 45259 3427 45315
rect 3483 45259 3569 45315
rect 3625 45259 3711 45315
rect 3767 45259 3853 45315
rect 3909 45259 3995 45315
rect 4051 45259 4137 45315
rect 4193 45259 4279 45315
rect 4335 45259 4421 45315
rect 4477 45259 4563 45315
rect 4619 45259 4705 45315
rect 4761 45259 4847 45315
rect 4903 45259 4989 45315
rect 5045 45259 5131 45315
rect 5187 45259 5273 45315
rect 5329 45259 5415 45315
rect 5471 45259 5557 45315
rect 5613 45259 5699 45315
rect 5755 45259 5841 45315
rect 5897 45259 5983 45315
rect 6039 45259 6125 45315
rect 6181 45259 6267 45315
rect 6323 45259 6409 45315
rect 6465 45259 6551 45315
rect 6607 45259 6693 45315
rect 6749 45259 6835 45315
rect 6891 45259 6977 45315
rect 7033 45259 7119 45315
rect 7175 45259 7261 45315
rect 7317 45259 7403 45315
rect 7459 45259 7545 45315
rect 7601 45259 7687 45315
rect 7743 45259 7829 45315
rect 7885 45259 7971 45315
rect 8027 45259 8113 45315
rect 8169 45259 8255 45315
rect 8311 45259 8397 45315
rect 8453 45259 8539 45315
rect 8595 45259 8681 45315
rect 8737 45259 8823 45315
rect 8879 45259 8965 45315
rect 9021 45259 9107 45315
rect 9163 45259 9249 45315
rect 9305 45259 9391 45315
rect 9447 45259 9533 45315
rect 9589 45259 9675 45315
rect 9731 45259 9817 45315
rect 9873 45259 9959 45315
rect 10015 45259 10101 45315
rect 10157 45259 10243 45315
rect 10299 45259 10385 45315
rect 10441 45259 10527 45315
rect 10583 45259 10669 45315
rect 10725 45259 10811 45315
rect 10867 45259 10953 45315
rect 11009 45259 11095 45315
rect 11151 45259 11237 45315
rect 11293 45259 11379 45315
rect 11435 45259 11521 45315
rect 11577 45259 11663 45315
rect 11719 45259 11805 45315
rect 11861 45259 11947 45315
rect 12003 45259 12089 45315
rect 12145 45259 12231 45315
rect 12287 45259 12373 45315
rect 12429 45259 12515 45315
rect 12571 45259 12657 45315
rect 12713 45259 12799 45315
rect 12855 45259 12941 45315
rect 12997 45259 13083 45315
rect 13139 45259 13225 45315
rect 13281 45259 13367 45315
rect 13423 45259 13509 45315
rect 13565 45259 13651 45315
rect 13707 45259 13793 45315
rect 13849 45259 13935 45315
rect 13991 45259 14077 45315
rect 14133 45259 14219 45315
rect 14275 45259 14361 45315
rect 14417 45259 14503 45315
rect 14559 45259 14645 45315
rect 14701 45259 14787 45315
rect 14843 45259 15000 45315
rect 0 45173 15000 45259
rect 0 45117 161 45173
rect 217 45117 303 45173
rect 359 45117 445 45173
rect 501 45117 587 45173
rect 643 45117 729 45173
rect 785 45117 871 45173
rect 927 45117 1013 45173
rect 1069 45117 1155 45173
rect 1211 45117 1297 45173
rect 1353 45117 1439 45173
rect 1495 45117 1581 45173
rect 1637 45117 1723 45173
rect 1779 45117 1865 45173
rect 1921 45117 2007 45173
rect 2063 45117 2149 45173
rect 2205 45117 2291 45173
rect 2347 45117 2433 45173
rect 2489 45117 2575 45173
rect 2631 45117 2717 45173
rect 2773 45117 2859 45173
rect 2915 45117 3001 45173
rect 3057 45117 3143 45173
rect 3199 45117 3285 45173
rect 3341 45117 3427 45173
rect 3483 45117 3569 45173
rect 3625 45117 3711 45173
rect 3767 45117 3853 45173
rect 3909 45117 3995 45173
rect 4051 45117 4137 45173
rect 4193 45117 4279 45173
rect 4335 45117 4421 45173
rect 4477 45117 4563 45173
rect 4619 45117 4705 45173
rect 4761 45117 4847 45173
rect 4903 45117 4989 45173
rect 5045 45117 5131 45173
rect 5187 45117 5273 45173
rect 5329 45117 5415 45173
rect 5471 45117 5557 45173
rect 5613 45117 5699 45173
rect 5755 45117 5841 45173
rect 5897 45117 5983 45173
rect 6039 45117 6125 45173
rect 6181 45117 6267 45173
rect 6323 45117 6409 45173
rect 6465 45117 6551 45173
rect 6607 45117 6693 45173
rect 6749 45117 6835 45173
rect 6891 45117 6977 45173
rect 7033 45117 7119 45173
rect 7175 45117 7261 45173
rect 7317 45117 7403 45173
rect 7459 45117 7545 45173
rect 7601 45117 7687 45173
rect 7743 45117 7829 45173
rect 7885 45117 7971 45173
rect 8027 45117 8113 45173
rect 8169 45117 8255 45173
rect 8311 45117 8397 45173
rect 8453 45117 8539 45173
rect 8595 45117 8681 45173
rect 8737 45117 8823 45173
rect 8879 45117 8965 45173
rect 9021 45117 9107 45173
rect 9163 45117 9249 45173
rect 9305 45117 9391 45173
rect 9447 45117 9533 45173
rect 9589 45117 9675 45173
rect 9731 45117 9817 45173
rect 9873 45117 9959 45173
rect 10015 45117 10101 45173
rect 10157 45117 10243 45173
rect 10299 45117 10385 45173
rect 10441 45117 10527 45173
rect 10583 45117 10669 45173
rect 10725 45117 10811 45173
rect 10867 45117 10953 45173
rect 11009 45117 11095 45173
rect 11151 45117 11237 45173
rect 11293 45117 11379 45173
rect 11435 45117 11521 45173
rect 11577 45117 11663 45173
rect 11719 45117 11805 45173
rect 11861 45117 11947 45173
rect 12003 45117 12089 45173
rect 12145 45117 12231 45173
rect 12287 45117 12373 45173
rect 12429 45117 12515 45173
rect 12571 45117 12657 45173
rect 12713 45117 12799 45173
rect 12855 45117 12941 45173
rect 12997 45117 13083 45173
rect 13139 45117 13225 45173
rect 13281 45117 13367 45173
rect 13423 45117 13509 45173
rect 13565 45117 13651 45173
rect 13707 45117 13793 45173
rect 13849 45117 13935 45173
rect 13991 45117 14077 45173
rect 14133 45117 14219 45173
rect 14275 45117 14361 45173
rect 14417 45117 14503 45173
rect 14559 45117 14645 45173
rect 14701 45117 14787 45173
rect 14843 45117 15000 45173
rect 0 45031 15000 45117
rect 0 44975 161 45031
rect 217 44975 303 45031
rect 359 44975 445 45031
rect 501 44975 587 45031
rect 643 44975 729 45031
rect 785 44975 871 45031
rect 927 44975 1013 45031
rect 1069 44975 1155 45031
rect 1211 44975 1297 45031
rect 1353 44975 1439 45031
rect 1495 44975 1581 45031
rect 1637 44975 1723 45031
rect 1779 44975 1865 45031
rect 1921 44975 2007 45031
rect 2063 44975 2149 45031
rect 2205 44975 2291 45031
rect 2347 44975 2433 45031
rect 2489 44975 2575 45031
rect 2631 44975 2717 45031
rect 2773 44975 2859 45031
rect 2915 44975 3001 45031
rect 3057 44975 3143 45031
rect 3199 44975 3285 45031
rect 3341 44975 3427 45031
rect 3483 44975 3569 45031
rect 3625 44975 3711 45031
rect 3767 44975 3853 45031
rect 3909 44975 3995 45031
rect 4051 44975 4137 45031
rect 4193 44975 4279 45031
rect 4335 44975 4421 45031
rect 4477 44975 4563 45031
rect 4619 44975 4705 45031
rect 4761 44975 4847 45031
rect 4903 44975 4989 45031
rect 5045 44975 5131 45031
rect 5187 44975 5273 45031
rect 5329 44975 5415 45031
rect 5471 44975 5557 45031
rect 5613 44975 5699 45031
rect 5755 44975 5841 45031
rect 5897 44975 5983 45031
rect 6039 44975 6125 45031
rect 6181 44975 6267 45031
rect 6323 44975 6409 45031
rect 6465 44975 6551 45031
rect 6607 44975 6693 45031
rect 6749 44975 6835 45031
rect 6891 44975 6977 45031
rect 7033 44975 7119 45031
rect 7175 44975 7261 45031
rect 7317 44975 7403 45031
rect 7459 44975 7545 45031
rect 7601 44975 7687 45031
rect 7743 44975 7829 45031
rect 7885 44975 7971 45031
rect 8027 44975 8113 45031
rect 8169 44975 8255 45031
rect 8311 44975 8397 45031
rect 8453 44975 8539 45031
rect 8595 44975 8681 45031
rect 8737 44975 8823 45031
rect 8879 44975 8965 45031
rect 9021 44975 9107 45031
rect 9163 44975 9249 45031
rect 9305 44975 9391 45031
rect 9447 44975 9533 45031
rect 9589 44975 9675 45031
rect 9731 44975 9817 45031
rect 9873 44975 9959 45031
rect 10015 44975 10101 45031
rect 10157 44975 10243 45031
rect 10299 44975 10385 45031
rect 10441 44975 10527 45031
rect 10583 44975 10669 45031
rect 10725 44975 10811 45031
rect 10867 44975 10953 45031
rect 11009 44975 11095 45031
rect 11151 44975 11237 45031
rect 11293 44975 11379 45031
rect 11435 44975 11521 45031
rect 11577 44975 11663 45031
rect 11719 44975 11805 45031
rect 11861 44975 11947 45031
rect 12003 44975 12089 45031
rect 12145 44975 12231 45031
rect 12287 44975 12373 45031
rect 12429 44975 12515 45031
rect 12571 44975 12657 45031
rect 12713 44975 12799 45031
rect 12855 44975 12941 45031
rect 12997 44975 13083 45031
rect 13139 44975 13225 45031
rect 13281 44975 13367 45031
rect 13423 44975 13509 45031
rect 13565 44975 13651 45031
rect 13707 44975 13793 45031
rect 13849 44975 13935 45031
rect 13991 44975 14077 45031
rect 14133 44975 14219 45031
rect 14275 44975 14361 45031
rect 14417 44975 14503 45031
rect 14559 44975 14645 45031
rect 14701 44975 14787 45031
rect 14843 44975 15000 45031
rect 0 44889 15000 44975
rect 0 44833 161 44889
rect 217 44833 303 44889
rect 359 44833 445 44889
rect 501 44833 587 44889
rect 643 44833 729 44889
rect 785 44833 871 44889
rect 927 44833 1013 44889
rect 1069 44833 1155 44889
rect 1211 44833 1297 44889
rect 1353 44833 1439 44889
rect 1495 44833 1581 44889
rect 1637 44833 1723 44889
rect 1779 44833 1865 44889
rect 1921 44833 2007 44889
rect 2063 44833 2149 44889
rect 2205 44833 2291 44889
rect 2347 44833 2433 44889
rect 2489 44833 2575 44889
rect 2631 44833 2717 44889
rect 2773 44833 2859 44889
rect 2915 44833 3001 44889
rect 3057 44833 3143 44889
rect 3199 44833 3285 44889
rect 3341 44833 3427 44889
rect 3483 44833 3569 44889
rect 3625 44833 3711 44889
rect 3767 44833 3853 44889
rect 3909 44833 3995 44889
rect 4051 44833 4137 44889
rect 4193 44833 4279 44889
rect 4335 44833 4421 44889
rect 4477 44833 4563 44889
rect 4619 44833 4705 44889
rect 4761 44833 4847 44889
rect 4903 44833 4989 44889
rect 5045 44833 5131 44889
rect 5187 44833 5273 44889
rect 5329 44833 5415 44889
rect 5471 44833 5557 44889
rect 5613 44833 5699 44889
rect 5755 44833 5841 44889
rect 5897 44833 5983 44889
rect 6039 44833 6125 44889
rect 6181 44833 6267 44889
rect 6323 44833 6409 44889
rect 6465 44833 6551 44889
rect 6607 44833 6693 44889
rect 6749 44833 6835 44889
rect 6891 44833 6977 44889
rect 7033 44833 7119 44889
rect 7175 44833 7261 44889
rect 7317 44833 7403 44889
rect 7459 44833 7545 44889
rect 7601 44833 7687 44889
rect 7743 44833 7829 44889
rect 7885 44833 7971 44889
rect 8027 44833 8113 44889
rect 8169 44833 8255 44889
rect 8311 44833 8397 44889
rect 8453 44833 8539 44889
rect 8595 44833 8681 44889
rect 8737 44833 8823 44889
rect 8879 44833 8965 44889
rect 9021 44833 9107 44889
rect 9163 44833 9249 44889
rect 9305 44833 9391 44889
rect 9447 44833 9533 44889
rect 9589 44833 9675 44889
rect 9731 44833 9817 44889
rect 9873 44833 9959 44889
rect 10015 44833 10101 44889
rect 10157 44833 10243 44889
rect 10299 44833 10385 44889
rect 10441 44833 10527 44889
rect 10583 44833 10669 44889
rect 10725 44833 10811 44889
rect 10867 44833 10953 44889
rect 11009 44833 11095 44889
rect 11151 44833 11237 44889
rect 11293 44833 11379 44889
rect 11435 44833 11521 44889
rect 11577 44833 11663 44889
rect 11719 44833 11805 44889
rect 11861 44833 11947 44889
rect 12003 44833 12089 44889
rect 12145 44833 12231 44889
rect 12287 44833 12373 44889
rect 12429 44833 12515 44889
rect 12571 44833 12657 44889
rect 12713 44833 12799 44889
rect 12855 44833 12941 44889
rect 12997 44833 13083 44889
rect 13139 44833 13225 44889
rect 13281 44833 13367 44889
rect 13423 44833 13509 44889
rect 13565 44833 13651 44889
rect 13707 44833 13793 44889
rect 13849 44833 13935 44889
rect 13991 44833 14077 44889
rect 14133 44833 14219 44889
rect 14275 44833 14361 44889
rect 14417 44833 14503 44889
rect 14559 44833 14645 44889
rect 14701 44833 14787 44889
rect 14843 44833 15000 44889
rect 0 44747 15000 44833
rect 0 44691 161 44747
rect 217 44691 303 44747
rect 359 44691 445 44747
rect 501 44691 587 44747
rect 643 44691 729 44747
rect 785 44691 871 44747
rect 927 44691 1013 44747
rect 1069 44691 1155 44747
rect 1211 44691 1297 44747
rect 1353 44691 1439 44747
rect 1495 44691 1581 44747
rect 1637 44691 1723 44747
rect 1779 44691 1865 44747
rect 1921 44691 2007 44747
rect 2063 44691 2149 44747
rect 2205 44691 2291 44747
rect 2347 44691 2433 44747
rect 2489 44691 2575 44747
rect 2631 44691 2717 44747
rect 2773 44691 2859 44747
rect 2915 44691 3001 44747
rect 3057 44691 3143 44747
rect 3199 44691 3285 44747
rect 3341 44691 3427 44747
rect 3483 44691 3569 44747
rect 3625 44691 3711 44747
rect 3767 44691 3853 44747
rect 3909 44691 3995 44747
rect 4051 44691 4137 44747
rect 4193 44691 4279 44747
rect 4335 44691 4421 44747
rect 4477 44691 4563 44747
rect 4619 44691 4705 44747
rect 4761 44691 4847 44747
rect 4903 44691 4989 44747
rect 5045 44691 5131 44747
rect 5187 44691 5273 44747
rect 5329 44691 5415 44747
rect 5471 44691 5557 44747
rect 5613 44691 5699 44747
rect 5755 44691 5841 44747
rect 5897 44691 5983 44747
rect 6039 44691 6125 44747
rect 6181 44691 6267 44747
rect 6323 44691 6409 44747
rect 6465 44691 6551 44747
rect 6607 44691 6693 44747
rect 6749 44691 6835 44747
rect 6891 44691 6977 44747
rect 7033 44691 7119 44747
rect 7175 44691 7261 44747
rect 7317 44691 7403 44747
rect 7459 44691 7545 44747
rect 7601 44691 7687 44747
rect 7743 44691 7829 44747
rect 7885 44691 7971 44747
rect 8027 44691 8113 44747
rect 8169 44691 8255 44747
rect 8311 44691 8397 44747
rect 8453 44691 8539 44747
rect 8595 44691 8681 44747
rect 8737 44691 8823 44747
rect 8879 44691 8965 44747
rect 9021 44691 9107 44747
rect 9163 44691 9249 44747
rect 9305 44691 9391 44747
rect 9447 44691 9533 44747
rect 9589 44691 9675 44747
rect 9731 44691 9817 44747
rect 9873 44691 9959 44747
rect 10015 44691 10101 44747
rect 10157 44691 10243 44747
rect 10299 44691 10385 44747
rect 10441 44691 10527 44747
rect 10583 44691 10669 44747
rect 10725 44691 10811 44747
rect 10867 44691 10953 44747
rect 11009 44691 11095 44747
rect 11151 44691 11237 44747
rect 11293 44691 11379 44747
rect 11435 44691 11521 44747
rect 11577 44691 11663 44747
rect 11719 44691 11805 44747
rect 11861 44691 11947 44747
rect 12003 44691 12089 44747
rect 12145 44691 12231 44747
rect 12287 44691 12373 44747
rect 12429 44691 12515 44747
rect 12571 44691 12657 44747
rect 12713 44691 12799 44747
rect 12855 44691 12941 44747
rect 12997 44691 13083 44747
rect 13139 44691 13225 44747
rect 13281 44691 13367 44747
rect 13423 44691 13509 44747
rect 13565 44691 13651 44747
rect 13707 44691 13793 44747
rect 13849 44691 13935 44747
rect 13991 44691 14077 44747
rect 14133 44691 14219 44747
rect 14275 44691 14361 44747
rect 14417 44691 14503 44747
rect 14559 44691 14645 44747
rect 14701 44691 14787 44747
rect 14843 44691 15000 44747
rect 0 44605 15000 44691
rect 0 44549 161 44605
rect 217 44549 303 44605
rect 359 44549 445 44605
rect 501 44549 587 44605
rect 643 44549 729 44605
rect 785 44549 871 44605
rect 927 44549 1013 44605
rect 1069 44549 1155 44605
rect 1211 44549 1297 44605
rect 1353 44549 1439 44605
rect 1495 44549 1581 44605
rect 1637 44549 1723 44605
rect 1779 44549 1865 44605
rect 1921 44549 2007 44605
rect 2063 44549 2149 44605
rect 2205 44549 2291 44605
rect 2347 44549 2433 44605
rect 2489 44549 2575 44605
rect 2631 44549 2717 44605
rect 2773 44549 2859 44605
rect 2915 44549 3001 44605
rect 3057 44549 3143 44605
rect 3199 44549 3285 44605
rect 3341 44549 3427 44605
rect 3483 44549 3569 44605
rect 3625 44549 3711 44605
rect 3767 44549 3853 44605
rect 3909 44549 3995 44605
rect 4051 44549 4137 44605
rect 4193 44549 4279 44605
rect 4335 44549 4421 44605
rect 4477 44549 4563 44605
rect 4619 44549 4705 44605
rect 4761 44549 4847 44605
rect 4903 44549 4989 44605
rect 5045 44549 5131 44605
rect 5187 44549 5273 44605
rect 5329 44549 5415 44605
rect 5471 44549 5557 44605
rect 5613 44549 5699 44605
rect 5755 44549 5841 44605
rect 5897 44549 5983 44605
rect 6039 44549 6125 44605
rect 6181 44549 6267 44605
rect 6323 44549 6409 44605
rect 6465 44549 6551 44605
rect 6607 44549 6693 44605
rect 6749 44549 6835 44605
rect 6891 44549 6977 44605
rect 7033 44549 7119 44605
rect 7175 44549 7261 44605
rect 7317 44549 7403 44605
rect 7459 44549 7545 44605
rect 7601 44549 7687 44605
rect 7743 44549 7829 44605
rect 7885 44549 7971 44605
rect 8027 44549 8113 44605
rect 8169 44549 8255 44605
rect 8311 44549 8397 44605
rect 8453 44549 8539 44605
rect 8595 44549 8681 44605
rect 8737 44549 8823 44605
rect 8879 44549 8965 44605
rect 9021 44549 9107 44605
rect 9163 44549 9249 44605
rect 9305 44549 9391 44605
rect 9447 44549 9533 44605
rect 9589 44549 9675 44605
rect 9731 44549 9817 44605
rect 9873 44549 9959 44605
rect 10015 44549 10101 44605
rect 10157 44549 10243 44605
rect 10299 44549 10385 44605
rect 10441 44549 10527 44605
rect 10583 44549 10669 44605
rect 10725 44549 10811 44605
rect 10867 44549 10953 44605
rect 11009 44549 11095 44605
rect 11151 44549 11237 44605
rect 11293 44549 11379 44605
rect 11435 44549 11521 44605
rect 11577 44549 11663 44605
rect 11719 44549 11805 44605
rect 11861 44549 11947 44605
rect 12003 44549 12089 44605
rect 12145 44549 12231 44605
rect 12287 44549 12373 44605
rect 12429 44549 12515 44605
rect 12571 44549 12657 44605
rect 12713 44549 12799 44605
rect 12855 44549 12941 44605
rect 12997 44549 13083 44605
rect 13139 44549 13225 44605
rect 13281 44549 13367 44605
rect 13423 44549 13509 44605
rect 13565 44549 13651 44605
rect 13707 44549 13793 44605
rect 13849 44549 13935 44605
rect 13991 44549 14077 44605
rect 14133 44549 14219 44605
rect 14275 44549 14361 44605
rect 14417 44549 14503 44605
rect 14559 44549 14645 44605
rect 14701 44549 14787 44605
rect 14843 44549 15000 44605
rect 0 44463 15000 44549
rect 0 44407 161 44463
rect 217 44407 303 44463
rect 359 44407 445 44463
rect 501 44407 587 44463
rect 643 44407 729 44463
rect 785 44407 871 44463
rect 927 44407 1013 44463
rect 1069 44407 1155 44463
rect 1211 44407 1297 44463
rect 1353 44407 1439 44463
rect 1495 44407 1581 44463
rect 1637 44407 1723 44463
rect 1779 44407 1865 44463
rect 1921 44407 2007 44463
rect 2063 44407 2149 44463
rect 2205 44407 2291 44463
rect 2347 44407 2433 44463
rect 2489 44407 2575 44463
rect 2631 44407 2717 44463
rect 2773 44407 2859 44463
rect 2915 44407 3001 44463
rect 3057 44407 3143 44463
rect 3199 44407 3285 44463
rect 3341 44407 3427 44463
rect 3483 44407 3569 44463
rect 3625 44407 3711 44463
rect 3767 44407 3853 44463
rect 3909 44407 3995 44463
rect 4051 44407 4137 44463
rect 4193 44407 4279 44463
rect 4335 44407 4421 44463
rect 4477 44407 4563 44463
rect 4619 44407 4705 44463
rect 4761 44407 4847 44463
rect 4903 44407 4989 44463
rect 5045 44407 5131 44463
rect 5187 44407 5273 44463
rect 5329 44407 5415 44463
rect 5471 44407 5557 44463
rect 5613 44407 5699 44463
rect 5755 44407 5841 44463
rect 5897 44407 5983 44463
rect 6039 44407 6125 44463
rect 6181 44407 6267 44463
rect 6323 44407 6409 44463
rect 6465 44407 6551 44463
rect 6607 44407 6693 44463
rect 6749 44407 6835 44463
rect 6891 44407 6977 44463
rect 7033 44407 7119 44463
rect 7175 44407 7261 44463
rect 7317 44407 7403 44463
rect 7459 44407 7545 44463
rect 7601 44407 7687 44463
rect 7743 44407 7829 44463
rect 7885 44407 7971 44463
rect 8027 44407 8113 44463
rect 8169 44407 8255 44463
rect 8311 44407 8397 44463
rect 8453 44407 8539 44463
rect 8595 44407 8681 44463
rect 8737 44407 8823 44463
rect 8879 44407 8965 44463
rect 9021 44407 9107 44463
rect 9163 44407 9249 44463
rect 9305 44407 9391 44463
rect 9447 44407 9533 44463
rect 9589 44407 9675 44463
rect 9731 44407 9817 44463
rect 9873 44407 9959 44463
rect 10015 44407 10101 44463
rect 10157 44407 10243 44463
rect 10299 44407 10385 44463
rect 10441 44407 10527 44463
rect 10583 44407 10669 44463
rect 10725 44407 10811 44463
rect 10867 44407 10953 44463
rect 11009 44407 11095 44463
rect 11151 44407 11237 44463
rect 11293 44407 11379 44463
rect 11435 44407 11521 44463
rect 11577 44407 11663 44463
rect 11719 44407 11805 44463
rect 11861 44407 11947 44463
rect 12003 44407 12089 44463
rect 12145 44407 12231 44463
rect 12287 44407 12373 44463
rect 12429 44407 12515 44463
rect 12571 44407 12657 44463
rect 12713 44407 12799 44463
rect 12855 44407 12941 44463
rect 12997 44407 13083 44463
rect 13139 44407 13225 44463
rect 13281 44407 13367 44463
rect 13423 44407 13509 44463
rect 13565 44407 13651 44463
rect 13707 44407 13793 44463
rect 13849 44407 13935 44463
rect 13991 44407 14077 44463
rect 14133 44407 14219 44463
rect 14275 44407 14361 44463
rect 14417 44407 14503 44463
rect 14559 44407 14645 44463
rect 14701 44407 14787 44463
rect 14843 44407 15000 44463
rect 0 44321 15000 44407
rect 0 44265 161 44321
rect 217 44265 303 44321
rect 359 44265 445 44321
rect 501 44265 587 44321
rect 643 44265 729 44321
rect 785 44265 871 44321
rect 927 44265 1013 44321
rect 1069 44265 1155 44321
rect 1211 44265 1297 44321
rect 1353 44265 1439 44321
rect 1495 44265 1581 44321
rect 1637 44265 1723 44321
rect 1779 44265 1865 44321
rect 1921 44265 2007 44321
rect 2063 44265 2149 44321
rect 2205 44265 2291 44321
rect 2347 44265 2433 44321
rect 2489 44265 2575 44321
rect 2631 44265 2717 44321
rect 2773 44265 2859 44321
rect 2915 44265 3001 44321
rect 3057 44265 3143 44321
rect 3199 44265 3285 44321
rect 3341 44265 3427 44321
rect 3483 44265 3569 44321
rect 3625 44265 3711 44321
rect 3767 44265 3853 44321
rect 3909 44265 3995 44321
rect 4051 44265 4137 44321
rect 4193 44265 4279 44321
rect 4335 44265 4421 44321
rect 4477 44265 4563 44321
rect 4619 44265 4705 44321
rect 4761 44265 4847 44321
rect 4903 44265 4989 44321
rect 5045 44265 5131 44321
rect 5187 44265 5273 44321
rect 5329 44265 5415 44321
rect 5471 44265 5557 44321
rect 5613 44265 5699 44321
rect 5755 44265 5841 44321
rect 5897 44265 5983 44321
rect 6039 44265 6125 44321
rect 6181 44265 6267 44321
rect 6323 44265 6409 44321
rect 6465 44265 6551 44321
rect 6607 44265 6693 44321
rect 6749 44265 6835 44321
rect 6891 44265 6977 44321
rect 7033 44265 7119 44321
rect 7175 44265 7261 44321
rect 7317 44265 7403 44321
rect 7459 44265 7545 44321
rect 7601 44265 7687 44321
rect 7743 44265 7829 44321
rect 7885 44265 7971 44321
rect 8027 44265 8113 44321
rect 8169 44265 8255 44321
rect 8311 44265 8397 44321
rect 8453 44265 8539 44321
rect 8595 44265 8681 44321
rect 8737 44265 8823 44321
rect 8879 44265 8965 44321
rect 9021 44265 9107 44321
rect 9163 44265 9249 44321
rect 9305 44265 9391 44321
rect 9447 44265 9533 44321
rect 9589 44265 9675 44321
rect 9731 44265 9817 44321
rect 9873 44265 9959 44321
rect 10015 44265 10101 44321
rect 10157 44265 10243 44321
rect 10299 44265 10385 44321
rect 10441 44265 10527 44321
rect 10583 44265 10669 44321
rect 10725 44265 10811 44321
rect 10867 44265 10953 44321
rect 11009 44265 11095 44321
rect 11151 44265 11237 44321
rect 11293 44265 11379 44321
rect 11435 44265 11521 44321
rect 11577 44265 11663 44321
rect 11719 44265 11805 44321
rect 11861 44265 11947 44321
rect 12003 44265 12089 44321
rect 12145 44265 12231 44321
rect 12287 44265 12373 44321
rect 12429 44265 12515 44321
rect 12571 44265 12657 44321
rect 12713 44265 12799 44321
rect 12855 44265 12941 44321
rect 12997 44265 13083 44321
rect 13139 44265 13225 44321
rect 13281 44265 13367 44321
rect 13423 44265 13509 44321
rect 13565 44265 13651 44321
rect 13707 44265 13793 44321
rect 13849 44265 13935 44321
rect 13991 44265 14077 44321
rect 14133 44265 14219 44321
rect 14275 44265 14361 44321
rect 14417 44265 14503 44321
rect 14559 44265 14645 44321
rect 14701 44265 14787 44321
rect 14843 44265 15000 44321
rect 0 44179 15000 44265
rect 0 44123 161 44179
rect 217 44123 303 44179
rect 359 44123 445 44179
rect 501 44123 587 44179
rect 643 44123 729 44179
rect 785 44123 871 44179
rect 927 44123 1013 44179
rect 1069 44123 1155 44179
rect 1211 44123 1297 44179
rect 1353 44123 1439 44179
rect 1495 44123 1581 44179
rect 1637 44123 1723 44179
rect 1779 44123 1865 44179
rect 1921 44123 2007 44179
rect 2063 44123 2149 44179
rect 2205 44123 2291 44179
rect 2347 44123 2433 44179
rect 2489 44123 2575 44179
rect 2631 44123 2717 44179
rect 2773 44123 2859 44179
rect 2915 44123 3001 44179
rect 3057 44123 3143 44179
rect 3199 44123 3285 44179
rect 3341 44123 3427 44179
rect 3483 44123 3569 44179
rect 3625 44123 3711 44179
rect 3767 44123 3853 44179
rect 3909 44123 3995 44179
rect 4051 44123 4137 44179
rect 4193 44123 4279 44179
rect 4335 44123 4421 44179
rect 4477 44123 4563 44179
rect 4619 44123 4705 44179
rect 4761 44123 4847 44179
rect 4903 44123 4989 44179
rect 5045 44123 5131 44179
rect 5187 44123 5273 44179
rect 5329 44123 5415 44179
rect 5471 44123 5557 44179
rect 5613 44123 5699 44179
rect 5755 44123 5841 44179
rect 5897 44123 5983 44179
rect 6039 44123 6125 44179
rect 6181 44123 6267 44179
rect 6323 44123 6409 44179
rect 6465 44123 6551 44179
rect 6607 44123 6693 44179
rect 6749 44123 6835 44179
rect 6891 44123 6977 44179
rect 7033 44123 7119 44179
rect 7175 44123 7261 44179
rect 7317 44123 7403 44179
rect 7459 44123 7545 44179
rect 7601 44123 7687 44179
rect 7743 44123 7829 44179
rect 7885 44123 7971 44179
rect 8027 44123 8113 44179
rect 8169 44123 8255 44179
rect 8311 44123 8397 44179
rect 8453 44123 8539 44179
rect 8595 44123 8681 44179
rect 8737 44123 8823 44179
rect 8879 44123 8965 44179
rect 9021 44123 9107 44179
rect 9163 44123 9249 44179
rect 9305 44123 9391 44179
rect 9447 44123 9533 44179
rect 9589 44123 9675 44179
rect 9731 44123 9817 44179
rect 9873 44123 9959 44179
rect 10015 44123 10101 44179
rect 10157 44123 10243 44179
rect 10299 44123 10385 44179
rect 10441 44123 10527 44179
rect 10583 44123 10669 44179
rect 10725 44123 10811 44179
rect 10867 44123 10953 44179
rect 11009 44123 11095 44179
rect 11151 44123 11237 44179
rect 11293 44123 11379 44179
rect 11435 44123 11521 44179
rect 11577 44123 11663 44179
rect 11719 44123 11805 44179
rect 11861 44123 11947 44179
rect 12003 44123 12089 44179
rect 12145 44123 12231 44179
rect 12287 44123 12373 44179
rect 12429 44123 12515 44179
rect 12571 44123 12657 44179
rect 12713 44123 12799 44179
rect 12855 44123 12941 44179
rect 12997 44123 13083 44179
rect 13139 44123 13225 44179
rect 13281 44123 13367 44179
rect 13423 44123 13509 44179
rect 13565 44123 13651 44179
rect 13707 44123 13793 44179
rect 13849 44123 13935 44179
rect 13991 44123 14077 44179
rect 14133 44123 14219 44179
rect 14275 44123 14361 44179
rect 14417 44123 14503 44179
rect 14559 44123 14645 44179
rect 14701 44123 14787 44179
rect 14843 44123 15000 44179
rect 0 44037 15000 44123
rect 0 43981 161 44037
rect 217 43981 303 44037
rect 359 43981 445 44037
rect 501 43981 587 44037
rect 643 43981 729 44037
rect 785 43981 871 44037
rect 927 43981 1013 44037
rect 1069 43981 1155 44037
rect 1211 43981 1297 44037
rect 1353 43981 1439 44037
rect 1495 43981 1581 44037
rect 1637 43981 1723 44037
rect 1779 43981 1865 44037
rect 1921 43981 2007 44037
rect 2063 43981 2149 44037
rect 2205 43981 2291 44037
rect 2347 43981 2433 44037
rect 2489 43981 2575 44037
rect 2631 43981 2717 44037
rect 2773 43981 2859 44037
rect 2915 43981 3001 44037
rect 3057 43981 3143 44037
rect 3199 43981 3285 44037
rect 3341 43981 3427 44037
rect 3483 43981 3569 44037
rect 3625 43981 3711 44037
rect 3767 43981 3853 44037
rect 3909 43981 3995 44037
rect 4051 43981 4137 44037
rect 4193 43981 4279 44037
rect 4335 43981 4421 44037
rect 4477 43981 4563 44037
rect 4619 43981 4705 44037
rect 4761 43981 4847 44037
rect 4903 43981 4989 44037
rect 5045 43981 5131 44037
rect 5187 43981 5273 44037
rect 5329 43981 5415 44037
rect 5471 43981 5557 44037
rect 5613 43981 5699 44037
rect 5755 43981 5841 44037
rect 5897 43981 5983 44037
rect 6039 43981 6125 44037
rect 6181 43981 6267 44037
rect 6323 43981 6409 44037
rect 6465 43981 6551 44037
rect 6607 43981 6693 44037
rect 6749 43981 6835 44037
rect 6891 43981 6977 44037
rect 7033 43981 7119 44037
rect 7175 43981 7261 44037
rect 7317 43981 7403 44037
rect 7459 43981 7545 44037
rect 7601 43981 7687 44037
rect 7743 43981 7829 44037
rect 7885 43981 7971 44037
rect 8027 43981 8113 44037
rect 8169 43981 8255 44037
rect 8311 43981 8397 44037
rect 8453 43981 8539 44037
rect 8595 43981 8681 44037
rect 8737 43981 8823 44037
rect 8879 43981 8965 44037
rect 9021 43981 9107 44037
rect 9163 43981 9249 44037
rect 9305 43981 9391 44037
rect 9447 43981 9533 44037
rect 9589 43981 9675 44037
rect 9731 43981 9817 44037
rect 9873 43981 9959 44037
rect 10015 43981 10101 44037
rect 10157 43981 10243 44037
rect 10299 43981 10385 44037
rect 10441 43981 10527 44037
rect 10583 43981 10669 44037
rect 10725 43981 10811 44037
rect 10867 43981 10953 44037
rect 11009 43981 11095 44037
rect 11151 43981 11237 44037
rect 11293 43981 11379 44037
rect 11435 43981 11521 44037
rect 11577 43981 11663 44037
rect 11719 43981 11805 44037
rect 11861 43981 11947 44037
rect 12003 43981 12089 44037
rect 12145 43981 12231 44037
rect 12287 43981 12373 44037
rect 12429 43981 12515 44037
rect 12571 43981 12657 44037
rect 12713 43981 12799 44037
rect 12855 43981 12941 44037
rect 12997 43981 13083 44037
rect 13139 43981 13225 44037
rect 13281 43981 13367 44037
rect 13423 43981 13509 44037
rect 13565 43981 13651 44037
rect 13707 43981 13793 44037
rect 13849 43981 13935 44037
rect 13991 43981 14077 44037
rect 14133 43981 14219 44037
rect 14275 43981 14361 44037
rect 14417 43981 14503 44037
rect 14559 43981 14645 44037
rect 14701 43981 14787 44037
rect 14843 43981 15000 44037
rect 0 43895 15000 43981
rect 0 43839 161 43895
rect 217 43839 303 43895
rect 359 43839 445 43895
rect 501 43839 587 43895
rect 643 43839 729 43895
rect 785 43839 871 43895
rect 927 43839 1013 43895
rect 1069 43839 1155 43895
rect 1211 43839 1297 43895
rect 1353 43839 1439 43895
rect 1495 43839 1581 43895
rect 1637 43839 1723 43895
rect 1779 43839 1865 43895
rect 1921 43839 2007 43895
rect 2063 43839 2149 43895
rect 2205 43839 2291 43895
rect 2347 43839 2433 43895
rect 2489 43839 2575 43895
rect 2631 43839 2717 43895
rect 2773 43839 2859 43895
rect 2915 43839 3001 43895
rect 3057 43839 3143 43895
rect 3199 43839 3285 43895
rect 3341 43839 3427 43895
rect 3483 43839 3569 43895
rect 3625 43839 3711 43895
rect 3767 43839 3853 43895
rect 3909 43839 3995 43895
rect 4051 43839 4137 43895
rect 4193 43839 4279 43895
rect 4335 43839 4421 43895
rect 4477 43839 4563 43895
rect 4619 43839 4705 43895
rect 4761 43839 4847 43895
rect 4903 43839 4989 43895
rect 5045 43839 5131 43895
rect 5187 43839 5273 43895
rect 5329 43839 5415 43895
rect 5471 43839 5557 43895
rect 5613 43839 5699 43895
rect 5755 43839 5841 43895
rect 5897 43839 5983 43895
rect 6039 43839 6125 43895
rect 6181 43839 6267 43895
rect 6323 43839 6409 43895
rect 6465 43839 6551 43895
rect 6607 43839 6693 43895
rect 6749 43839 6835 43895
rect 6891 43839 6977 43895
rect 7033 43839 7119 43895
rect 7175 43839 7261 43895
rect 7317 43839 7403 43895
rect 7459 43839 7545 43895
rect 7601 43839 7687 43895
rect 7743 43839 7829 43895
rect 7885 43839 7971 43895
rect 8027 43839 8113 43895
rect 8169 43839 8255 43895
rect 8311 43839 8397 43895
rect 8453 43839 8539 43895
rect 8595 43839 8681 43895
rect 8737 43839 8823 43895
rect 8879 43839 8965 43895
rect 9021 43839 9107 43895
rect 9163 43839 9249 43895
rect 9305 43839 9391 43895
rect 9447 43839 9533 43895
rect 9589 43839 9675 43895
rect 9731 43839 9817 43895
rect 9873 43839 9959 43895
rect 10015 43839 10101 43895
rect 10157 43839 10243 43895
rect 10299 43839 10385 43895
rect 10441 43839 10527 43895
rect 10583 43839 10669 43895
rect 10725 43839 10811 43895
rect 10867 43839 10953 43895
rect 11009 43839 11095 43895
rect 11151 43839 11237 43895
rect 11293 43839 11379 43895
rect 11435 43839 11521 43895
rect 11577 43839 11663 43895
rect 11719 43839 11805 43895
rect 11861 43839 11947 43895
rect 12003 43839 12089 43895
rect 12145 43839 12231 43895
rect 12287 43839 12373 43895
rect 12429 43839 12515 43895
rect 12571 43839 12657 43895
rect 12713 43839 12799 43895
rect 12855 43839 12941 43895
rect 12997 43839 13083 43895
rect 13139 43839 13225 43895
rect 13281 43839 13367 43895
rect 13423 43839 13509 43895
rect 13565 43839 13651 43895
rect 13707 43839 13793 43895
rect 13849 43839 13935 43895
rect 13991 43839 14077 43895
rect 14133 43839 14219 43895
rect 14275 43839 14361 43895
rect 14417 43839 14503 43895
rect 14559 43839 14645 43895
rect 14701 43839 14787 43895
rect 14843 43839 15000 43895
rect 0 43753 15000 43839
rect 0 43697 161 43753
rect 217 43697 303 43753
rect 359 43697 445 43753
rect 501 43697 587 43753
rect 643 43697 729 43753
rect 785 43697 871 43753
rect 927 43697 1013 43753
rect 1069 43697 1155 43753
rect 1211 43697 1297 43753
rect 1353 43697 1439 43753
rect 1495 43697 1581 43753
rect 1637 43697 1723 43753
rect 1779 43697 1865 43753
rect 1921 43697 2007 43753
rect 2063 43697 2149 43753
rect 2205 43697 2291 43753
rect 2347 43697 2433 43753
rect 2489 43697 2575 43753
rect 2631 43697 2717 43753
rect 2773 43697 2859 43753
rect 2915 43697 3001 43753
rect 3057 43697 3143 43753
rect 3199 43697 3285 43753
rect 3341 43697 3427 43753
rect 3483 43697 3569 43753
rect 3625 43697 3711 43753
rect 3767 43697 3853 43753
rect 3909 43697 3995 43753
rect 4051 43697 4137 43753
rect 4193 43697 4279 43753
rect 4335 43697 4421 43753
rect 4477 43697 4563 43753
rect 4619 43697 4705 43753
rect 4761 43697 4847 43753
rect 4903 43697 4989 43753
rect 5045 43697 5131 43753
rect 5187 43697 5273 43753
rect 5329 43697 5415 43753
rect 5471 43697 5557 43753
rect 5613 43697 5699 43753
rect 5755 43697 5841 43753
rect 5897 43697 5983 43753
rect 6039 43697 6125 43753
rect 6181 43697 6267 43753
rect 6323 43697 6409 43753
rect 6465 43697 6551 43753
rect 6607 43697 6693 43753
rect 6749 43697 6835 43753
rect 6891 43697 6977 43753
rect 7033 43697 7119 43753
rect 7175 43697 7261 43753
rect 7317 43697 7403 43753
rect 7459 43697 7545 43753
rect 7601 43697 7687 43753
rect 7743 43697 7829 43753
rect 7885 43697 7971 43753
rect 8027 43697 8113 43753
rect 8169 43697 8255 43753
rect 8311 43697 8397 43753
rect 8453 43697 8539 43753
rect 8595 43697 8681 43753
rect 8737 43697 8823 43753
rect 8879 43697 8965 43753
rect 9021 43697 9107 43753
rect 9163 43697 9249 43753
rect 9305 43697 9391 43753
rect 9447 43697 9533 43753
rect 9589 43697 9675 43753
rect 9731 43697 9817 43753
rect 9873 43697 9959 43753
rect 10015 43697 10101 43753
rect 10157 43697 10243 43753
rect 10299 43697 10385 43753
rect 10441 43697 10527 43753
rect 10583 43697 10669 43753
rect 10725 43697 10811 43753
rect 10867 43697 10953 43753
rect 11009 43697 11095 43753
rect 11151 43697 11237 43753
rect 11293 43697 11379 43753
rect 11435 43697 11521 43753
rect 11577 43697 11663 43753
rect 11719 43697 11805 43753
rect 11861 43697 11947 43753
rect 12003 43697 12089 43753
rect 12145 43697 12231 43753
rect 12287 43697 12373 43753
rect 12429 43697 12515 43753
rect 12571 43697 12657 43753
rect 12713 43697 12799 43753
rect 12855 43697 12941 43753
rect 12997 43697 13083 43753
rect 13139 43697 13225 43753
rect 13281 43697 13367 43753
rect 13423 43697 13509 43753
rect 13565 43697 13651 43753
rect 13707 43697 13793 43753
rect 13849 43697 13935 43753
rect 13991 43697 14077 43753
rect 14133 43697 14219 43753
rect 14275 43697 14361 43753
rect 14417 43697 14503 43753
rect 14559 43697 14645 43753
rect 14701 43697 14787 43753
rect 14843 43697 15000 43753
rect 0 43611 15000 43697
rect 0 43555 161 43611
rect 217 43555 303 43611
rect 359 43555 445 43611
rect 501 43555 587 43611
rect 643 43555 729 43611
rect 785 43555 871 43611
rect 927 43555 1013 43611
rect 1069 43555 1155 43611
rect 1211 43555 1297 43611
rect 1353 43555 1439 43611
rect 1495 43555 1581 43611
rect 1637 43555 1723 43611
rect 1779 43555 1865 43611
rect 1921 43555 2007 43611
rect 2063 43555 2149 43611
rect 2205 43555 2291 43611
rect 2347 43555 2433 43611
rect 2489 43555 2575 43611
rect 2631 43555 2717 43611
rect 2773 43555 2859 43611
rect 2915 43555 3001 43611
rect 3057 43555 3143 43611
rect 3199 43555 3285 43611
rect 3341 43555 3427 43611
rect 3483 43555 3569 43611
rect 3625 43555 3711 43611
rect 3767 43555 3853 43611
rect 3909 43555 3995 43611
rect 4051 43555 4137 43611
rect 4193 43555 4279 43611
rect 4335 43555 4421 43611
rect 4477 43555 4563 43611
rect 4619 43555 4705 43611
rect 4761 43555 4847 43611
rect 4903 43555 4989 43611
rect 5045 43555 5131 43611
rect 5187 43555 5273 43611
rect 5329 43555 5415 43611
rect 5471 43555 5557 43611
rect 5613 43555 5699 43611
rect 5755 43555 5841 43611
rect 5897 43555 5983 43611
rect 6039 43555 6125 43611
rect 6181 43555 6267 43611
rect 6323 43555 6409 43611
rect 6465 43555 6551 43611
rect 6607 43555 6693 43611
rect 6749 43555 6835 43611
rect 6891 43555 6977 43611
rect 7033 43555 7119 43611
rect 7175 43555 7261 43611
rect 7317 43555 7403 43611
rect 7459 43555 7545 43611
rect 7601 43555 7687 43611
rect 7743 43555 7829 43611
rect 7885 43555 7971 43611
rect 8027 43555 8113 43611
rect 8169 43555 8255 43611
rect 8311 43555 8397 43611
rect 8453 43555 8539 43611
rect 8595 43555 8681 43611
rect 8737 43555 8823 43611
rect 8879 43555 8965 43611
rect 9021 43555 9107 43611
rect 9163 43555 9249 43611
rect 9305 43555 9391 43611
rect 9447 43555 9533 43611
rect 9589 43555 9675 43611
rect 9731 43555 9817 43611
rect 9873 43555 9959 43611
rect 10015 43555 10101 43611
rect 10157 43555 10243 43611
rect 10299 43555 10385 43611
rect 10441 43555 10527 43611
rect 10583 43555 10669 43611
rect 10725 43555 10811 43611
rect 10867 43555 10953 43611
rect 11009 43555 11095 43611
rect 11151 43555 11237 43611
rect 11293 43555 11379 43611
rect 11435 43555 11521 43611
rect 11577 43555 11663 43611
rect 11719 43555 11805 43611
rect 11861 43555 11947 43611
rect 12003 43555 12089 43611
rect 12145 43555 12231 43611
rect 12287 43555 12373 43611
rect 12429 43555 12515 43611
rect 12571 43555 12657 43611
rect 12713 43555 12799 43611
rect 12855 43555 12941 43611
rect 12997 43555 13083 43611
rect 13139 43555 13225 43611
rect 13281 43555 13367 43611
rect 13423 43555 13509 43611
rect 13565 43555 13651 43611
rect 13707 43555 13793 43611
rect 13849 43555 13935 43611
rect 13991 43555 14077 43611
rect 14133 43555 14219 43611
rect 14275 43555 14361 43611
rect 14417 43555 14503 43611
rect 14559 43555 14645 43611
rect 14701 43555 14787 43611
rect 14843 43555 15000 43611
rect 0 43469 15000 43555
rect 0 43413 161 43469
rect 217 43413 303 43469
rect 359 43413 445 43469
rect 501 43413 587 43469
rect 643 43413 729 43469
rect 785 43413 871 43469
rect 927 43413 1013 43469
rect 1069 43413 1155 43469
rect 1211 43413 1297 43469
rect 1353 43413 1439 43469
rect 1495 43413 1581 43469
rect 1637 43413 1723 43469
rect 1779 43413 1865 43469
rect 1921 43413 2007 43469
rect 2063 43413 2149 43469
rect 2205 43413 2291 43469
rect 2347 43413 2433 43469
rect 2489 43413 2575 43469
rect 2631 43413 2717 43469
rect 2773 43413 2859 43469
rect 2915 43413 3001 43469
rect 3057 43413 3143 43469
rect 3199 43413 3285 43469
rect 3341 43413 3427 43469
rect 3483 43413 3569 43469
rect 3625 43413 3711 43469
rect 3767 43413 3853 43469
rect 3909 43413 3995 43469
rect 4051 43413 4137 43469
rect 4193 43413 4279 43469
rect 4335 43413 4421 43469
rect 4477 43413 4563 43469
rect 4619 43413 4705 43469
rect 4761 43413 4847 43469
rect 4903 43413 4989 43469
rect 5045 43413 5131 43469
rect 5187 43413 5273 43469
rect 5329 43413 5415 43469
rect 5471 43413 5557 43469
rect 5613 43413 5699 43469
rect 5755 43413 5841 43469
rect 5897 43413 5983 43469
rect 6039 43413 6125 43469
rect 6181 43413 6267 43469
rect 6323 43413 6409 43469
rect 6465 43413 6551 43469
rect 6607 43413 6693 43469
rect 6749 43413 6835 43469
rect 6891 43413 6977 43469
rect 7033 43413 7119 43469
rect 7175 43413 7261 43469
rect 7317 43413 7403 43469
rect 7459 43413 7545 43469
rect 7601 43413 7687 43469
rect 7743 43413 7829 43469
rect 7885 43413 7971 43469
rect 8027 43413 8113 43469
rect 8169 43413 8255 43469
rect 8311 43413 8397 43469
rect 8453 43413 8539 43469
rect 8595 43413 8681 43469
rect 8737 43413 8823 43469
rect 8879 43413 8965 43469
rect 9021 43413 9107 43469
rect 9163 43413 9249 43469
rect 9305 43413 9391 43469
rect 9447 43413 9533 43469
rect 9589 43413 9675 43469
rect 9731 43413 9817 43469
rect 9873 43413 9959 43469
rect 10015 43413 10101 43469
rect 10157 43413 10243 43469
rect 10299 43413 10385 43469
rect 10441 43413 10527 43469
rect 10583 43413 10669 43469
rect 10725 43413 10811 43469
rect 10867 43413 10953 43469
rect 11009 43413 11095 43469
rect 11151 43413 11237 43469
rect 11293 43413 11379 43469
rect 11435 43413 11521 43469
rect 11577 43413 11663 43469
rect 11719 43413 11805 43469
rect 11861 43413 11947 43469
rect 12003 43413 12089 43469
rect 12145 43413 12231 43469
rect 12287 43413 12373 43469
rect 12429 43413 12515 43469
rect 12571 43413 12657 43469
rect 12713 43413 12799 43469
rect 12855 43413 12941 43469
rect 12997 43413 13083 43469
rect 13139 43413 13225 43469
rect 13281 43413 13367 43469
rect 13423 43413 13509 43469
rect 13565 43413 13651 43469
rect 13707 43413 13793 43469
rect 13849 43413 13935 43469
rect 13991 43413 14077 43469
rect 14133 43413 14219 43469
rect 14275 43413 14361 43469
rect 14417 43413 14503 43469
rect 14559 43413 14645 43469
rect 14701 43413 14787 43469
rect 14843 43413 15000 43469
rect 0 43327 15000 43413
rect 0 43271 161 43327
rect 217 43271 303 43327
rect 359 43271 445 43327
rect 501 43271 587 43327
rect 643 43271 729 43327
rect 785 43271 871 43327
rect 927 43271 1013 43327
rect 1069 43271 1155 43327
rect 1211 43271 1297 43327
rect 1353 43271 1439 43327
rect 1495 43271 1581 43327
rect 1637 43271 1723 43327
rect 1779 43271 1865 43327
rect 1921 43271 2007 43327
rect 2063 43271 2149 43327
rect 2205 43271 2291 43327
rect 2347 43271 2433 43327
rect 2489 43271 2575 43327
rect 2631 43271 2717 43327
rect 2773 43271 2859 43327
rect 2915 43271 3001 43327
rect 3057 43271 3143 43327
rect 3199 43271 3285 43327
rect 3341 43271 3427 43327
rect 3483 43271 3569 43327
rect 3625 43271 3711 43327
rect 3767 43271 3853 43327
rect 3909 43271 3995 43327
rect 4051 43271 4137 43327
rect 4193 43271 4279 43327
rect 4335 43271 4421 43327
rect 4477 43271 4563 43327
rect 4619 43271 4705 43327
rect 4761 43271 4847 43327
rect 4903 43271 4989 43327
rect 5045 43271 5131 43327
rect 5187 43271 5273 43327
rect 5329 43271 5415 43327
rect 5471 43271 5557 43327
rect 5613 43271 5699 43327
rect 5755 43271 5841 43327
rect 5897 43271 5983 43327
rect 6039 43271 6125 43327
rect 6181 43271 6267 43327
rect 6323 43271 6409 43327
rect 6465 43271 6551 43327
rect 6607 43271 6693 43327
rect 6749 43271 6835 43327
rect 6891 43271 6977 43327
rect 7033 43271 7119 43327
rect 7175 43271 7261 43327
rect 7317 43271 7403 43327
rect 7459 43271 7545 43327
rect 7601 43271 7687 43327
rect 7743 43271 7829 43327
rect 7885 43271 7971 43327
rect 8027 43271 8113 43327
rect 8169 43271 8255 43327
rect 8311 43271 8397 43327
rect 8453 43271 8539 43327
rect 8595 43271 8681 43327
rect 8737 43271 8823 43327
rect 8879 43271 8965 43327
rect 9021 43271 9107 43327
rect 9163 43271 9249 43327
rect 9305 43271 9391 43327
rect 9447 43271 9533 43327
rect 9589 43271 9675 43327
rect 9731 43271 9817 43327
rect 9873 43271 9959 43327
rect 10015 43271 10101 43327
rect 10157 43271 10243 43327
rect 10299 43271 10385 43327
rect 10441 43271 10527 43327
rect 10583 43271 10669 43327
rect 10725 43271 10811 43327
rect 10867 43271 10953 43327
rect 11009 43271 11095 43327
rect 11151 43271 11237 43327
rect 11293 43271 11379 43327
rect 11435 43271 11521 43327
rect 11577 43271 11663 43327
rect 11719 43271 11805 43327
rect 11861 43271 11947 43327
rect 12003 43271 12089 43327
rect 12145 43271 12231 43327
rect 12287 43271 12373 43327
rect 12429 43271 12515 43327
rect 12571 43271 12657 43327
rect 12713 43271 12799 43327
rect 12855 43271 12941 43327
rect 12997 43271 13083 43327
rect 13139 43271 13225 43327
rect 13281 43271 13367 43327
rect 13423 43271 13509 43327
rect 13565 43271 13651 43327
rect 13707 43271 13793 43327
rect 13849 43271 13935 43327
rect 13991 43271 14077 43327
rect 14133 43271 14219 43327
rect 14275 43271 14361 43327
rect 14417 43271 14503 43327
rect 14559 43271 14645 43327
rect 14701 43271 14787 43327
rect 14843 43271 15000 43327
rect 0 43185 15000 43271
rect 0 43129 161 43185
rect 217 43129 303 43185
rect 359 43129 445 43185
rect 501 43129 587 43185
rect 643 43129 729 43185
rect 785 43129 871 43185
rect 927 43129 1013 43185
rect 1069 43129 1155 43185
rect 1211 43129 1297 43185
rect 1353 43129 1439 43185
rect 1495 43129 1581 43185
rect 1637 43129 1723 43185
rect 1779 43129 1865 43185
rect 1921 43129 2007 43185
rect 2063 43129 2149 43185
rect 2205 43129 2291 43185
rect 2347 43129 2433 43185
rect 2489 43129 2575 43185
rect 2631 43129 2717 43185
rect 2773 43129 2859 43185
rect 2915 43129 3001 43185
rect 3057 43129 3143 43185
rect 3199 43129 3285 43185
rect 3341 43129 3427 43185
rect 3483 43129 3569 43185
rect 3625 43129 3711 43185
rect 3767 43129 3853 43185
rect 3909 43129 3995 43185
rect 4051 43129 4137 43185
rect 4193 43129 4279 43185
rect 4335 43129 4421 43185
rect 4477 43129 4563 43185
rect 4619 43129 4705 43185
rect 4761 43129 4847 43185
rect 4903 43129 4989 43185
rect 5045 43129 5131 43185
rect 5187 43129 5273 43185
rect 5329 43129 5415 43185
rect 5471 43129 5557 43185
rect 5613 43129 5699 43185
rect 5755 43129 5841 43185
rect 5897 43129 5983 43185
rect 6039 43129 6125 43185
rect 6181 43129 6267 43185
rect 6323 43129 6409 43185
rect 6465 43129 6551 43185
rect 6607 43129 6693 43185
rect 6749 43129 6835 43185
rect 6891 43129 6977 43185
rect 7033 43129 7119 43185
rect 7175 43129 7261 43185
rect 7317 43129 7403 43185
rect 7459 43129 7545 43185
rect 7601 43129 7687 43185
rect 7743 43129 7829 43185
rect 7885 43129 7971 43185
rect 8027 43129 8113 43185
rect 8169 43129 8255 43185
rect 8311 43129 8397 43185
rect 8453 43129 8539 43185
rect 8595 43129 8681 43185
rect 8737 43129 8823 43185
rect 8879 43129 8965 43185
rect 9021 43129 9107 43185
rect 9163 43129 9249 43185
rect 9305 43129 9391 43185
rect 9447 43129 9533 43185
rect 9589 43129 9675 43185
rect 9731 43129 9817 43185
rect 9873 43129 9959 43185
rect 10015 43129 10101 43185
rect 10157 43129 10243 43185
rect 10299 43129 10385 43185
rect 10441 43129 10527 43185
rect 10583 43129 10669 43185
rect 10725 43129 10811 43185
rect 10867 43129 10953 43185
rect 11009 43129 11095 43185
rect 11151 43129 11237 43185
rect 11293 43129 11379 43185
rect 11435 43129 11521 43185
rect 11577 43129 11663 43185
rect 11719 43129 11805 43185
rect 11861 43129 11947 43185
rect 12003 43129 12089 43185
rect 12145 43129 12231 43185
rect 12287 43129 12373 43185
rect 12429 43129 12515 43185
rect 12571 43129 12657 43185
rect 12713 43129 12799 43185
rect 12855 43129 12941 43185
rect 12997 43129 13083 43185
rect 13139 43129 13225 43185
rect 13281 43129 13367 43185
rect 13423 43129 13509 43185
rect 13565 43129 13651 43185
rect 13707 43129 13793 43185
rect 13849 43129 13935 43185
rect 13991 43129 14077 43185
rect 14133 43129 14219 43185
rect 14275 43129 14361 43185
rect 14417 43129 14503 43185
rect 14559 43129 14645 43185
rect 14701 43129 14787 43185
rect 14843 43129 15000 43185
rect 0 43043 15000 43129
rect 0 42987 161 43043
rect 217 42987 303 43043
rect 359 42987 445 43043
rect 501 42987 587 43043
rect 643 42987 729 43043
rect 785 42987 871 43043
rect 927 42987 1013 43043
rect 1069 42987 1155 43043
rect 1211 42987 1297 43043
rect 1353 42987 1439 43043
rect 1495 42987 1581 43043
rect 1637 42987 1723 43043
rect 1779 42987 1865 43043
rect 1921 42987 2007 43043
rect 2063 42987 2149 43043
rect 2205 42987 2291 43043
rect 2347 42987 2433 43043
rect 2489 42987 2575 43043
rect 2631 42987 2717 43043
rect 2773 42987 2859 43043
rect 2915 42987 3001 43043
rect 3057 42987 3143 43043
rect 3199 42987 3285 43043
rect 3341 42987 3427 43043
rect 3483 42987 3569 43043
rect 3625 42987 3711 43043
rect 3767 42987 3853 43043
rect 3909 42987 3995 43043
rect 4051 42987 4137 43043
rect 4193 42987 4279 43043
rect 4335 42987 4421 43043
rect 4477 42987 4563 43043
rect 4619 42987 4705 43043
rect 4761 42987 4847 43043
rect 4903 42987 4989 43043
rect 5045 42987 5131 43043
rect 5187 42987 5273 43043
rect 5329 42987 5415 43043
rect 5471 42987 5557 43043
rect 5613 42987 5699 43043
rect 5755 42987 5841 43043
rect 5897 42987 5983 43043
rect 6039 42987 6125 43043
rect 6181 42987 6267 43043
rect 6323 42987 6409 43043
rect 6465 42987 6551 43043
rect 6607 42987 6693 43043
rect 6749 42987 6835 43043
rect 6891 42987 6977 43043
rect 7033 42987 7119 43043
rect 7175 42987 7261 43043
rect 7317 42987 7403 43043
rect 7459 42987 7545 43043
rect 7601 42987 7687 43043
rect 7743 42987 7829 43043
rect 7885 42987 7971 43043
rect 8027 42987 8113 43043
rect 8169 42987 8255 43043
rect 8311 42987 8397 43043
rect 8453 42987 8539 43043
rect 8595 42987 8681 43043
rect 8737 42987 8823 43043
rect 8879 42987 8965 43043
rect 9021 42987 9107 43043
rect 9163 42987 9249 43043
rect 9305 42987 9391 43043
rect 9447 42987 9533 43043
rect 9589 42987 9675 43043
rect 9731 42987 9817 43043
rect 9873 42987 9959 43043
rect 10015 42987 10101 43043
rect 10157 42987 10243 43043
rect 10299 42987 10385 43043
rect 10441 42987 10527 43043
rect 10583 42987 10669 43043
rect 10725 42987 10811 43043
rect 10867 42987 10953 43043
rect 11009 42987 11095 43043
rect 11151 42987 11237 43043
rect 11293 42987 11379 43043
rect 11435 42987 11521 43043
rect 11577 42987 11663 43043
rect 11719 42987 11805 43043
rect 11861 42987 11947 43043
rect 12003 42987 12089 43043
rect 12145 42987 12231 43043
rect 12287 42987 12373 43043
rect 12429 42987 12515 43043
rect 12571 42987 12657 43043
rect 12713 42987 12799 43043
rect 12855 42987 12941 43043
rect 12997 42987 13083 43043
rect 13139 42987 13225 43043
rect 13281 42987 13367 43043
rect 13423 42987 13509 43043
rect 13565 42987 13651 43043
rect 13707 42987 13793 43043
rect 13849 42987 13935 43043
rect 13991 42987 14077 43043
rect 14133 42987 14219 43043
rect 14275 42987 14361 43043
rect 14417 42987 14503 43043
rect 14559 42987 14645 43043
rect 14701 42987 14787 43043
rect 14843 42987 15000 43043
rect 0 42901 15000 42987
rect 0 42845 161 42901
rect 217 42845 303 42901
rect 359 42845 445 42901
rect 501 42845 587 42901
rect 643 42845 729 42901
rect 785 42845 871 42901
rect 927 42845 1013 42901
rect 1069 42845 1155 42901
rect 1211 42845 1297 42901
rect 1353 42845 1439 42901
rect 1495 42845 1581 42901
rect 1637 42845 1723 42901
rect 1779 42845 1865 42901
rect 1921 42845 2007 42901
rect 2063 42845 2149 42901
rect 2205 42845 2291 42901
rect 2347 42845 2433 42901
rect 2489 42845 2575 42901
rect 2631 42845 2717 42901
rect 2773 42845 2859 42901
rect 2915 42845 3001 42901
rect 3057 42845 3143 42901
rect 3199 42845 3285 42901
rect 3341 42845 3427 42901
rect 3483 42845 3569 42901
rect 3625 42845 3711 42901
rect 3767 42845 3853 42901
rect 3909 42845 3995 42901
rect 4051 42845 4137 42901
rect 4193 42845 4279 42901
rect 4335 42845 4421 42901
rect 4477 42845 4563 42901
rect 4619 42845 4705 42901
rect 4761 42845 4847 42901
rect 4903 42845 4989 42901
rect 5045 42845 5131 42901
rect 5187 42845 5273 42901
rect 5329 42845 5415 42901
rect 5471 42845 5557 42901
rect 5613 42845 5699 42901
rect 5755 42845 5841 42901
rect 5897 42845 5983 42901
rect 6039 42845 6125 42901
rect 6181 42845 6267 42901
rect 6323 42845 6409 42901
rect 6465 42845 6551 42901
rect 6607 42845 6693 42901
rect 6749 42845 6835 42901
rect 6891 42845 6977 42901
rect 7033 42845 7119 42901
rect 7175 42845 7261 42901
rect 7317 42845 7403 42901
rect 7459 42845 7545 42901
rect 7601 42845 7687 42901
rect 7743 42845 7829 42901
rect 7885 42845 7971 42901
rect 8027 42845 8113 42901
rect 8169 42845 8255 42901
rect 8311 42845 8397 42901
rect 8453 42845 8539 42901
rect 8595 42845 8681 42901
rect 8737 42845 8823 42901
rect 8879 42845 8965 42901
rect 9021 42845 9107 42901
rect 9163 42845 9249 42901
rect 9305 42845 9391 42901
rect 9447 42845 9533 42901
rect 9589 42845 9675 42901
rect 9731 42845 9817 42901
rect 9873 42845 9959 42901
rect 10015 42845 10101 42901
rect 10157 42845 10243 42901
rect 10299 42845 10385 42901
rect 10441 42845 10527 42901
rect 10583 42845 10669 42901
rect 10725 42845 10811 42901
rect 10867 42845 10953 42901
rect 11009 42845 11095 42901
rect 11151 42845 11237 42901
rect 11293 42845 11379 42901
rect 11435 42845 11521 42901
rect 11577 42845 11663 42901
rect 11719 42845 11805 42901
rect 11861 42845 11947 42901
rect 12003 42845 12089 42901
rect 12145 42845 12231 42901
rect 12287 42845 12373 42901
rect 12429 42845 12515 42901
rect 12571 42845 12657 42901
rect 12713 42845 12799 42901
rect 12855 42845 12941 42901
rect 12997 42845 13083 42901
rect 13139 42845 13225 42901
rect 13281 42845 13367 42901
rect 13423 42845 13509 42901
rect 13565 42845 13651 42901
rect 13707 42845 13793 42901
rect 13849 42845 13935 42901
rect 13991 42845 14077 42901
rect 14133 42845 14219 42901
rect 14275 42845 14361 42901
rect 14417 42845 14503 42901
rect 14559 42845 14645 42901
rect 14701 42845 14787 42901
rect 14843 42845 15000 42901
rect 0 42800 15000 42845
rect 937 42600 3937 42800
rect 4337 42600 7337 42800
rect 7737 42600 10737 42800
rect 11137 42600 14137 42800
rect 0 42563 15000 42600
rect 0 42507 161 42563
rect 217 42507 303 42563
rect 359 42507 445 42563
rect 501 42507 587 42563
rect 643 42507 729 42563
rect 785 42507 871 42563
rect 927 42507 1013 42563
rect 1069 42507 1155 42563
rect 1211 42507 1297 42563
rect 1353 42507 1439 42563
rect 1495 42507 1581 42563
rect 1637 42507 1723 42563
rect 1779 42507 1865 42563
rect 1921 42507 2007 42563
rect 2063 42507 2149 42563
rect 2205 42507 2291 42563
rect 2347 42507 2433 42563
rect 2489 42507 2575 42563
rect 2631 42507 2717 42563
rect 2773 42507 2859 42563
rect 2915 42507 3001 42563
rect 3057 42507 3143 42563
rect 3199 42507 3285 42563
rect 3341 42507 3427 42563
rect 3483 42507 3569 42563
rect 3625 42507 3711 42563
rect 3767 42507 3853 42563
rect 3909 42507 3995 42563
rect 4051 42507 4137 42563
rect 4193 42507 4279 42563
rect 4335 42507 4421 42563
rect 4477 42507 4563 42563
rect 4619 42507 4705 42563
rect 4761 42507 4847 42563
rect 4903 42507 4989 42563
rect 5045 42507 5131 42563
rect 5187 42507 5273 42563
rect 5329 42507 5415 42563
rect 5471 42507 5557 42563
rect 5613 42507 5699 42563
rect 5755 42507 5841 42563
rect 5897 42507 5983 42563
rect 6039 42507 6125 42563
rect 6181 42507 6267 42563
rect 6323 42507 6409 42563
rect 6465 42507 6551 42563
rect 6607 42507 6693 42563
rect 6749 42507 6835 42563
rect 6891 42507 6977 42563
rect 7033 42507 7119 42563
rect 7175 42507 7261 42563
rect 7317 42507 7403 42563
rect 7459 42507 7545 42563
rect 7601 42507 7687 42563
rect 7743 42507 7829 42563
rect 7885 42507 7971 42563
rect 8027 42507 8113 42563
rect 8169 42507 8255 42563
rect 8311 42507 8397 42563
rect 8453 42507 8539 42563
rect 8595 42507 8681 42563
rect 8737 42507 8823 42563
rect 8879 42507 8965 42563
rect 9021 42507 9107 42563
rect 9163 42507 9249 42563
rect 9305 42507 9391 42563
rect 9447 42507 9533 42563
rect 9589 42507 9675 42563
rect 9731 42507 9817 42563
rect 9873 42507 9959 42563
rect 10015 42507 10101 42563
rect 10157 42507 10243 42563
rect 10299 42507 10385 42563
rect 10441 42507 10527 42563
rect 10583 42507 10669 42563
rect 10725 42507 10811 42563
rect 10867 42507 10953 42563
rect 11009 42507 11095 42563
rect 11151 42507 11237 42563
rect 11293 42507 11379 42563
rect 11435 42507 11521 42563
rect 11577 42507 11663 42563
rect 11719 42507 11805 42563
rect 11861 42507 11947 42563
rect 12003 42507 12089 42563
rect 12145 42507 12231 42563
rect 12287 42507 12373 42563
rect 12429 42507 12515 42563
rect 12571 42507 12657 42563
rect 12713 42507 12799 42563
rect 12855 42507 12941 42563
rect 12997 42507 13083 42563
rect 13139 42507 13225 42563
rect 13281 42507 13367 42563
rect 13423 42507 13509 42563
rect 13565 42507 13651 42563
rect 13707 42507 13793 42563
rect 13849 42507 13935 42563
rect 13991 42507 14077 42563
rect 14133 42507 14219 42563
rect 14275 42507 14361 42563
rect 14417 42507 14503 42563
rect 14559 42507 14645 42563
rect 14701 42507 14787 42563
rect 14843 42507 15000 42563
rect 0 42421 15000 42507
rect 0 42365 161 42421
rect 217 42365 303 42421
rect 359 42365 445 42421
rect 501 42365 587 42421
rect 643 42365 729 42421
rect 785 42365 871 42421
rect 927 42365 1013 42421
rect 1069 42365 1155 42421
rect 1211 42365 1297 42421
rect 1353 42365 1439 42421
rect 1495 42365 1581 42421
rect 1637 42365 1723 42421
rect 1779 42365 1865 42421
rect 1921 42365 2007 42421
rect 2063 42365 2149 42421
rect 2205 42365 2291 42421
rect 2347 42365 2433 42421
rect 2489 42365 2575 42421
rect 2631 42365 2717 42421
rect 2773 42365 2859 42421
rect 2915 42365 3001 42421
rect 3057 42365 3143 42421
rect 3199 42365 3285 42421
rect 3341 42365 3427 42421
rect 3483 42365 3569 42421
rect 3625 42365 3711 42421
rect 3767 42365 3853 42421
rect 3909 42365 3995 42421
rect 4051 42365 4137 42421
rect 4193 42365 4279 42421
rect 4335 42365 4421 42421
rect 4477 42365 4563 42421
rect 4619 42365 4705 42421
rect 4761 42365 4847 42421
rect 4903 42365 4989 42421
rect 5045 42365 5131 42421
rect 5187 42365 5273 42421
rect 5329 42365 5415 42421
rect 5471 42365 5557 42421
rect 5613 42365 5699 42421
rect 5755 42365 5841 42421
rect 5897 42365 5983 42421
rect 6039 42365 6125 42421
rect 6181 42365 6267 42421
rect 6323 42365 6409 42421
rect 6465 42365 6551 42421
rect 6607 42365 6693 42421
rect 6749 42365 6835 42421
rect 6891 42365 6977 42421
rect 7033 42365 7119 42421
rect 7175 42365 7261 42421
rect 7317 42365 7403 42421
rect 7459 42365 7545 42421
rect 7601 42365 7687 42421
rect 7743 42365 7829 42421
rect 7885 42365 7971 42421
rect 8027 42365 8113 42421
rect 8169 42365 8255 42421
rect 8311 42365 8397 42421
rect 8453 42365 8539 42421
rect 8595 42365 8681 42421
rect 8737 42365 8823 42421
rect 8879 42365 8965 42421
rect 9021 42365 9107 42421
rect 9163 42365 9249 42421
rect 9305 42365 9391 42421
rect 9447 42365 9533 42421
rect 9589 42365 9675 42421
rect 9731 42365 9817 42421
rect 9873 42365 9959 42421
rect 10015 42365 10101 42421
rect 10157 42365 10243 42421
rect 10299 42365 10385 42421
rect 10441 42365 10527 42421
rect 10583 42365 10669 42421
rect 10725 42365 10811 42421
rect 10867 42365 10953 42421
rect 11009 42365 11095 42421
rect 11151 42365 11237 42421
rect 11293 42365 11379 42421
rect 11435 42365 11521 42421
rect 11577 42365 11663 42421
rect 11719 42365 11805 42421
rect 11861 42365 11947 42421
rect 12003 42365 12089 42421
rect 12145 42365 12231 42421
rect 12287 42365 12373 42421
rect 12429 42365 12515 42421
rect 12571 42365 12657 42421
rect 12713 42365 12799 42421
rect 12855 42365 12941 42421
rect 12997 42365 13083 42421
rect 13139 42365 13225 42421
rect 13281 42365 13367 42421
rect 13423 42365 13509 42421
rect 13565 42365 13651 42421
rect 13707 42365 13793 42421
rect 13849 42365 13935 42421
rect 13991 42365 14077 42421
rect 14133 42365 14219 42421
rect 14275 42365 14361 42421
rect 14417 42365 14503 42421
rect 14559 42365 14645 42421
rect 14701 42365 14787 42421
rect 14843 42365 15000 42421
rect 0 42279 15000 42365
rect 0 42223 161 42279
rect 217 42223 303 42279
rect 359 42223 445 42279
rect 501 42223 587 42279
rect 643 42223 729 42279
rect 785 42223 871 42279
rect 927 42223 1013 42279
rect 1069 42223 1155 42279
rect 1211 42223 1297 42279
rect 1353 42223 1439 42279
rect 1495 42223 1581 42279
rect 1637 42223 1723 42279
rect 1779 42223 1865 42279
rect 1921 42223 2007 42279
rect 2063 42223 2149 42279
rect 2205 42223 2291 42279
rect 2347 42223 2433 42279
rect 2489 42223 2575 42279
rect 2631 42223 2717 42279
rect 2773 42223 2859 42279
rect 2915 42223 3001 42279
rect 3057 42223 3143 42279
rect 3199 42223 3285 42279
rect 3341 42223 3427 42279
rect 3483 42223 3569 42279
rect 3625 42223 3711 42279
rect 3767 42223 3853 42279
rect 3909 42223 3995 42279
rect 4051 42223 4137 42279
rect 4193 42223 4279 42279
rect 4335 42223 4421 42279
rect 4477 42223 4563 42279
rect 4619 42223 4705 42279
rect 4761 42223 4847 42279
rect 4903 42223 4989 42279
rect 5045 42223 5131 42279
rect 5187 42223 5273 42279
rect 5329 42223 5415 42279
rect 5471 42223 5557 42279
rect 5613 42223 5699 42279
rect 5755 42223 5841 42279
rect 5897 42223 5983 42279
rect 6039 42223 6125 42279
rect 6181 42223 6267 42279
rect 6323 42223 6409 42279
rect 6465 42223 6551 42279
rect 6607 42223 6693 42279
rect 6749 42223 6835 42279
rect 6891 42223 6977 42279
rect 7033 42223 7119 42279
rect 7175 42223 7261 42279
rect 7317 42223 7403 42279
rect 7459 42223 7545 42279
rect 7601 42223 7687 42279
rect 7743 42223 7829 42279
rect 7885 42223 7971 42279
rect 8027 42223 8113 42279
rect 8169 42223 8255 42279
rect 8311 42223 8397 42279
rect 8453 42223 8539 42279
rect 8595 42223 8681 42279
rect 8737 42223 8823 42279
rect 8879 42223 8965 42279
rect 9021 42223 9107 42279
rect 9163 42223 9249 42279
rect 9305 42223 9391 42279
rect 9447 42223 9533 42279
rect 9589 42223 9675 42279
rect 9731 42223 9817 42279
rect 9873 42223 9959 42279
rect 10015 42223 10101 42279
rect 10157 42223 10243 42279
rect 10299 42223 10385 42279
rect 10441 42223 10527 42279
rect 10583 42223 10669 42279
rect 10725 42223 10811 42279
rect 10867 42223 10953 42279
rect 11009 42223 11095 42279
rect 11151 42223 11237 42279
rect 11293 42223 11379 42279
rect 11435 42223 11521 42279
rect 11577 42223 11663 42279
rect 11719 42223 11805 42279
rect 11861 42223 11947 42279
rect 12003 42223 12089 42279
rect 12145 42223 12231 42279
rect 12287 42223 12373 42279
rect 12429 42223 12515 42279
rect 12571 42223 12657 42279
rect 12713 42223 12799 42279
rect 12855 42223 12941 42279
rect 12997 42223 13083 42279
rect 13139 42223 13225 42279
rect 13281 42223 13367 42279
rect 13423 42223 13509 42279
rect 13565 42223 13651 42279
rect 13707 42223 13793 42279
rect 13849 42223 13935 42279
rect 13991 42223 14077 42279
rect 14133 42223 14219 42279
rect 14275 42223 14361 42279
rect 14417 42223 14503 42279
rect 14559 42223 14645 42279
rect 14701 42223 14787 42279
rect 14843 42223 15000 42279
rect 0 42137 15000 42223
rect 0 42081 161 42137
rect 217 42081 303 42137
rect 359 42081 445 42137
rect 501 42081 587 42137
rect 643 42081 729 42137
rect 785 42081 871 42137
rect 927 42081 1013 42137
rect 1069 42081 1155 42137
rect 1211 42081 1297 42137
rect 1353 42081 1439 42137
rect 1495 42081 1581 42137
rect 1637 42081 1723 42137
rect 1779 42081 1865 42137
rect 1921 42081 2007 42137
rect 2063 42081 2149 42137
rect 2205 42081 2291 42137
rect 2347 42081 2433 42137
rect 2489 42081 2575 42137
rect 2631 42081 2717 42137
rect 2773 42081 2859 42137
rect 2915 42081 3001 42137
rect 3057 42081 3143 42137
rect 3199 42081 3285 42137
rect 3341 42081 3427 42137
rect 3483 42081 3569 42137
rect 3625 42081 3711 42137
rect 3767 42081 3853 42137
rect 3909 42081 3995 42137
rect 4051 42081 4137 42137
rect 4193 42081 4279 42137
rect 4335 42081 4421 42137
rect 4477 42081 4563 42137
rect 4619 42081 4705 42137
rect 4761 42081 4847 42137
rect 4903 42081 4989 42137
rect 5045 42081 5131 42137
rect 5187 42081 5273 42137
rect 5329 42081 5415 42137
rect 5471 42081 5557 42137
rect 5613 42081 5699 42137
rect 5755 42081 5841 42137
rect 5897 42081 5983 42137
rect 6039 42081 6125 42137
rect 6181 42081 6267 42137
rect 6323 42081 6409 42137
rect 6465 42081 6551 42137
rect 6607 42081 6693 42137
rect 6749 42081 6835 42137
rect 6891 42081 6977 42137
rect 7033 42081 7119 42137
rect 7175 42081 7261 42137
rect 7317 42081 7403 42137
rect 7459 42081 7545 42137
rect 7601 42081 7687 42137
rect 7743 42081 7829 42137
rect 7885 42081 7971 42137
rect 8027 42081 8113 42137
rect 8169 42081 8255 42137
rect 8311 42081 8397 42137
rect 8453 42081 8539 42137
rect 8595 42081 8681 42137
rect 8737 42081 8823 42137
rect 8879 42081 8965 42137
rect 9021 42081 9107 42137
rect 9163 42081 9249 42137
rect 9305 42081 9391 42137
rect 9447 42081 9533 42137
rect 9589 42081 9675 42137
rect 9731 42081 9817 42137
rect 9873 42081 9959 42137
rect 10015 42081 10101 42137
rect 10157 42081 10243 42137
rect 10299 42081 10385 42137
rect 10441 42081 10527 42137
rect 10583 42081 10669 42137
rect 10725 42081 10811 42137
rect 10867 42081 10953 42137
rect 11009 42081 11095 42137
rect 11151 42081 11237 42137
rect 11293 42081 11379 42137
rect 11435 42081 11521 42137
rect 11577 42081 11663 42137
rect 11719 42081 11805 42137
rect 11861 42081 11947 42137
rect 12003 42081 12089 42137
rect 12145 42081 12231 42137
rect 12287 42081 12373 42137
rect 12429 42081 12515 42137
rect 12571 42081 12657 42137
rect 12713 42081 12799 42137
rect 12855 42081 12941 42137
rect 12997 42081 13083 42137
rect 13139 42081 13225 42137
rect 13281 42081 13367 42137
rect 13423 42081 13509 42137
rect 13565 42081 13651 42137
rect 13707 42081 13793 42137
rect 13849 42081 13935 42137
rect 13991 42081 14077 42137
rect 14133 42081 14219 42137
rect 14275 42081 14361 42137
rect 14417 42081 14503 42137
rect 14559 42081 14645 42137
rect 14701 42081 14787 42137
rect 14843 42081 15000 42137
rect 0 41995 15000 42081
rect 0 41939 161 41995
rect 217 41939 303 41995
rect 359 41939 445 41995
rect 501 41939 587 41995
rect 643 41939 729 41995
rect 785 41939 871 41995
rect 927 41939 1013 41995
rect 1069 41939 1155 41995
rect 1211 41939 1297 41995
rect 1353 41939 1439 41995
rect 1495 41939 1581 41995
rect 1637 41939 1723 41995
rect 1779 41939 1865 41995
rect 1921 41939 2007 41995
rect 2063 41939 2149 41995
rect 2205 41939 2291 41995
rect 2347 41939 2433 41995
rect 2489 41939 2575 41995
rect 2631 41939 2717 41995
rect 2773 41939 2859 41995
rect 2915 41939 3001 41995
rect 3057 41939 3143 41995
rect 3199 41939 3285 41995
rect 3341 41939 3427 41995
rect 3483 41939 3569 41995
rect 3625 41939 3711 41995
rect 3767 41939 3853 41995
rect 3909 41939 3995 41995
rect 4051 41939 4137 41995
rect 4193 41939 4279 41995
rect 4335 41939 4421 41995
rect 4477 41939 4563 41995
rect 4619 41939 4705 41995
rect 4761 41939 4847 41995
rect 4903 41939 4989 41995
rect 5045 41939 5131 41995
rect 5187 41939 5273 41995
rect 5329 41939 5415 41995
rect 5471 41939 5557 41995
rect 5613 41939 5699 41995
rect 5755 41939 5841 41995
rect 5897 41939 5983 41995
rect 6039 41939 6125 41995
rect 6181 41939 6267 41995
rect 6323 41939 6409 41995
rect 6465 41939 6551 41995
rect 6607 41939 6693 41995
rect 6749 41939 6835 41995
rect 6891 41939 6977 41995
rect 7033 41939 7119 41995
rect 7175 41939 7261 41995
rect 7317 41939 7403 41995
rect 7459 41939 7545 41995
rect 7601 41939 7687 41995
rect 7743 41939 7829 41995
rect 7885 41939 7971 41995
rect 8027 41939 8113 41995
rect 8169 41939 8255 41995
rect 8311 41939 8397 41995
rect 8453 41939 8539 41995
rect 8595 41939 8681 41995
rect 8737 41939 8823 41995
rect 8879 41939 8965 41995
rect 9021 41939 9107 41995
rect 9163 41939 9249 41995
rect 9305 41939 9391 41995
rect 9447 41939 9533 41995
rect 9589 41939 9675 41995
rect 9731 41939 9817 41995
rect 9873 41939 9959 41995
rect 10015 41939 10101 41995
rect 10157 41939 10243 41995
rect 10299 41939 10385 41995
rect 10441 41939 10527 41995
rect 10583 41939 10669 41995
rect 10725 41939 10811 41995
rect 10867 41939 10953 41995
rect 11009 41939 11095 41995
rect 11151 41939 11237 41995
rect 11293 41939 11379 41995
rect 11435 41939 11521 41995
rect 11577 41939 11663 41995
rect 11719 41939 11805 41995
rect 11861 41939 11947 41995
rect 12003 41939 12089 41995
rect 12145 41939 12231 41995
rect 12287 41939 12373 41995
rect 12429 41939 12515 41995
rect 12571 41939 12657 41995
rect 12713 41939 12799 41995
rect 12855 41939 12941 41995
rect 12997 41939 13083 41995
rect 13139 41939 13225 41995
rect 13281 41939 13367 41995
rect 13423 41939 13509 41995
rect 13565 41939 13651 41995
rect 13707 41939 13793 41995
rect 13849 41939 13935 41995
rect 13991 41939 14077 41995
rect 14133 41939 14219 41995
rect 14275 41939 14361 41995
rect 14417 41939 14503 41995
rect 14559 41939 14645 41995
rect 14701 41939 14787 41995
rect 14843 41939 15000 41995
rect 0 41853 15000 41939
rect 0 41797 161 41853
rect 217 41797 303 41853
rect 359 41797 445 41853
rect 501 41797 587 41853
rect 643 41797 729 41853
rect 785 41797 871 41853
rect 927 41797 1013 41853
rect 1069 41797 1155 41853
rect 1211 41797 1297 41853
rect 1353 41797 1439 41853
rect 1495 41797 1581 41853
rect 1637 41797 1723 41853
rect 1779 41797 1865 41853
rect 1921 41797 2007 41853
rect 2063 41797 2149 41853
rect 2205 41797 2291 41853
rect 2347 41797 2433 41853
rect 2489 41797 2575 41853
rect 2631 41797 2717 41853
rect 2773 41797 2859 41853
rect 2915 41797 3001 41853
rect 3057 41797 3143 41853
rect 3199 41797 3285 41853
rect 3341 41797 3427 41853
rect 3483 41797 3569 41853
rect 3625 41797 3711 41853
rect 3767 41797 3853 41853
rect 3909 41797 3995 41853
rect 4051 41797 4137 41853
rect 4193 41797 4279 41853
rect 4335 41797 4421 41853
rect 4477 41797 4563 41853
rect 4619 41797 4705 41853
rect 4761 41797 4847 41853
rect 4903 41797 4989 41853
rect 5045 41797 5131 41853
rect 5187 41797 5273 41853
rect 5329 41797 5415 41853
rect 5471 41797 5557 41853
rect 5613 41797 5699 41853
rect 5755 41797 5841 41853
rect 5897 41797 5983 41853
rect 6039 41797 6125 41853
rect 6181 41797 6267 41853
rect 6323 41797 6409 41853
rect 6465 41797 6551 41853
rect 6607 41797 6693 41853
rect 6749 41797 6835 41853
rect 6891 41797 6977 41853
rect 7033 41797 7119 41853
rect 7175 41797 7261 41853
rect 7317 41797 7403 41853
rect 7459 41797 7545 41853
rect 7601 41797 7687 41853
rect 7743 41797 7829 41853
rect 7885 41797 7971 41853
rect 8027 41797 8113 41853
rect 8169 41797 8255 41853
rect 8311 41797 8397 41853
rect 8453 41797 8539 41853
rect 8595 41797 8681 41853
rect 8737 41797 8823 41853
rect 8879 41797 8965 41853
rect 9021 41797 9107 41853
rect 9163 41797 9249 41853
rect 9305 41797 9391 41853
rect 9447 41797 9533 41853
rect 9589 41797 9675 41853
rect 9731 41797 9817 41853
rect 9873 41797 9959 41853
rect 10015 41797 10101 41853
rect 10157 41797 10243 41853
rect 10299 41797 10385 41853
rect 10441 41797 10527 41853
rect 10583 41797 10669 41853
rect 10725 41797 10811 41853
rect 10867 41797 10953 41853
rect 11009 41797 11095 41853
rect 11151 41797 11237 41853
rect 11293 41797 11379 41853
rect 11435 41797 11521 41853
rect 11577 41797 11663 41853
rect 11719 41797 11805 41853
rect 11861 41797 11947 41853
rect 12003 41797 12089 41853
rect 12145 41797 12231 41853
rect 12287 41797 12373 41853
rect 12429 41797 12515 41853
rect 12571 41797 12657 41853
rect 12713 41797 12799 41853
rect 12855 41797 12941 41853
rect 12997 41797 13083 41853
rect 13139 41797 13225 41853
rect 13281 41797 13367 41853
rect 13423 41797 13509 41853
rect 13565 41797 13651 41853
rect 13707 41797 13793 41853
rect 13849 41797 13935 41853
rect 13991 41797 14077 41853
rect 14133 41797 14219 41853
rect 14275 41797 14361 41853
rect 14417 41797 14503 41853
rect 14559 41797 14645 41853
rect 14701 41797 14787 41853
rect 14843 41797 15000 41853
rect 0 41711 15000 41797
rect 0 41655 161 41711
rect 217 41655 303 41711
rect 359 41655 445 41711
rect 501 41655 587 41711
rect 643 41655 729 41711
rect 785 41655 871 41711
rect 927 41655 1013 41711
rect 1069 41655 1155 41711
rect 1211 41655 1297 41711
rect 1353 41655 1439 41711
rect 1495 41655 1581 41711
rect 1637 41655 1723 41711
rect 1779 41655 1865 41711
rect 1921 41655 2007 41711
rect 2063 41655 2149 41711
rect 2205 41655 2291 41711
rect 2347 41655 2433 41711
rect 2489 41655 2575 41711
rect 2631 41655 2717 41711
rect 2773 41655 2859 41711
rect 2915 41655 3001 41711
rect 3057 41655 3143 41711
rect 3199 41655 3285 41711
rect 3341 41655 3427 41711
rect 3483 41655 3569 41711
rect 3625 41655 3711 41711
rect 3767 41655 3853 41711
rect 3909 41655 3995 41711
rect 4051 41655 4137 41711
rect 4193 41655 4279 41711
rect 4335 41655 4421 41711
rect 4477 41655 4563 41711
rect 4619 41655 4705 41711
rect 4761 41655 4847 41711
rect 4903 41655 4989 41711
rect 5045 41655 5131 41711
rect 5187 41655 5273 41711
rect 5329 41655 5415 41711
rect 5471 41655 5557 41711
rect 5613 41655 5699 41711
rect 5755 41655 5841 41711
rect 5897 41655 5983 41711
rect 6039 41655 6125 41711
rect 6181 41655 6267 41711
rect 6323 41655 6409 41711
rect 6465 41655 6551 41711
rect 6607 41655 6693 41711
rect 6749 41655 6835 41711
rect 6891 41655 6977 41711
rect 7033 41655 7119 41711
rect 7175 41655 7261 41711
rect 7317 41655 7403 41711
rect 7459 41655 7545 41711
rect 7601 41655 7687 41711
rect 7743 41655 7829 41711
rect 7885 41655 7971 41711
rect 8027 41655 8113 41711
rect 8169 41655 8255 41711
rect 8311 41655 8397 41711
rect 8453 41655 8539 41711
rect 8595 41655 8681 41711
rect 8737 41655 8823 41711
rect 8879 41655 8965 41711
rect 9021 41655 9107 41711
rect 9163 41655 9249 41711
rect 9305 41655 9391 41711
rect 9447 41655 9533 41711
rect 9589 41655 9675 41711
rect 9731 41655 9817 41711
rect 9873 41655 9959 41711
rect 10015 41655 10101 41711
rect 10157 41655 10243 41711
rect 10299 41655 10385 41711
rect 10441 41655 10527 41711
rect 10583 41655 10669 41711
rect 10725 41655 10811 41711
rect 10867 41655 10953 41711
rect 11009 41655 11095 41711
rect 11151 41655 11237 41711
rect 11293 41655 11379 41711
rect 11435 41655 11521 41711
rect 11577 41655 11663 41711
rect 11719 41655 11805 41711
rect 11861 41655 11947 41711
rect 12003 41655 12089 41711
rect 12145 41655 12231 41711
rect 12287 41655 12373 41711
rect 12429 41655 12515 41711
rect 12571 41655 12657 41711
rect 12713 41655 12799 41711
rect 12855 41655 12941 41711
rect 12997 41655 13083 41711
rect 13139 41655 13225 41711
rect 13281 41655 13367 41711
rect 13423 41655 13509 41711
rect 13565 41655 13651 41711
rect 13707 41655 13793 41711
rect 13849 41655 13935 41711
rect 13991 41655 14077 41711
rect 14133 41655 14219 41711
rect 14275 41655 14361 41711
rect 14417 41655 14503 41711
rect 14559 41655 14645 41711
rect 14701 41655 14787 41711
rect 14843 41655 15000 41711
rect 0 41569 15000 41655
rect 0 41513 161 41569
rect 217 41513 303 41569
rect 359 41513 445 41569
rect 501 41513 587 41569
rect 643 41513 729 41569
rect 785 41513 871 41569
rect 927 41513 1013 41569
rect 1069 41513 1155 41569
rect 1211 41513 1297 41569
rect 1353 41513 1439 41569
rect 1495 41513 1581 41569
rect 1637 41513 1723 41569
rect 1779 41513 1865 41569
rect 1921 41513 2007 41569
rect 2063 41513 2149 41569
rect 2205 41513 2291 41569
rect 2347 41513 2433 41569
rect 2489 41513 2575 41569
rect 2631 41513 2717 41569
rect 2773 41513 2859 41569
rect 2915 41513 3001 41569
rect 3057 41513 3143 41569
rect 3199 41513 3285 41569
rect 3341 41513 3427 41569
rect 3483 41513 3569 41569
rect 3625 41513 3711 41569
rect 3767 41513 3853 41569
rect 3909 41513 3995 41569
rect 4051 41513 4137 41569
rect 4193 41513 4279 41569
rect 4335 41513 4421 41569
rect 4477 41513 4563 41569
rect 4619 41513 4705 41569
rect 4761 41513 4847 41569
rect 4903 41513 4989 41569
rect 5045 41513 5131 41569
rect 5187 41513 5273 41569
rect 5329 41513 5415 41569
rect 5471 41513 5557 41569
rect 5613 41513 5699 41569
rect 5755 41513 5841 41569
rect 5897 41513 5983 41569
rect 6039 41513 6125 41569
rect 6181 41513 6267 41569
rect 6323 41513 6409 41569
rect 6465 41513 6551 41569
rect 6607 41513 6693 41569
rect 6749 41513 6835 41569
rect 6891 41513 6977 41569
rect 7033 41513 7119 41569
rect 7175 41513 7261 41569
rect 7317 41513 7403 41569
rect 7459 41513 7545 41569
rect 7601 41513 7687 41569
rect 7743 41513 7829 41569
rect 7885 41513 7971 41569
rect 8027 41513 8113 41569
rect 8169 41513 8255 41569
rect 8311 41513 8397 41569
rect 8453 41513 8539 41569
rect 8595 41513 8681 41569
rect 8737 41513 8823 41569
rect 8879 41513 8965 41569
rect 9021 41513 9107 41569
rect 9163 41513 9249 41569
rect 9305 41513 9391 41569
rect 9447 41513 9533 41569
rect 9589 41513 9675 41569
rect 9731 41513 9817 41569
rect 9873 41513 9959 41569
rect 10015 41513 10101 41569
rect 10157 41513 10243 41569
rect 10299 41513 10385 41569
rect 10441 41513 10527 41569
rect 10583 41513 10669 41569
rect 10725 41513 10811 41569
rect 10867 41513 10953 41569
rect 11009 41513 11095 41569
rect 11151 41513 11237 41569
rect 11293 41513 11379 41569
rect 11435 41513 11521 41569
rect 11577 41513 11663 41569
rect 11719 41513 11805 41569
rect 11861 41513 11947 41569
rect 12003 41513 12089 41569
rect 12145 41513 12231 41569
rect 12287 41513 12373 41569
rect 12429 41513 12515 41569
rect 12571 41513 12657 41569
rect 12713 41513 12799 41569
rect 12855 41513 12941 41569
rect 12997 41513 13083 41569
rect 13139 41513 13225 41569
rect 13281 41513 13367 41569
rect 13423 41513 13509 41569
rect 13565 41513 13651 41569
rect 13707 41513 13793 41569
rect 13849 41513 13935 41569
rect 13991 41513 14077 41569
rect 14133 41513 14219 41569
rect 14275 41513 14361 41569
rect 14417 41513 14503 41569
rect 14559 41513 14645 41569
rect 14701 41513 14787 41569
rect 14843 41513 15000 41569
rect 0 41427 15000 41513
rect 0 41371 161 41427
rect 217 41371 303 41427
rect 359 41371 445 41427
rect 501 41371 587 41427
rect 643 41371 729 41427
rect 785 41371 871 41427
rect 927 41371 1013 41427
rect 1069 41371 1155 41427
rect 1211 41371 1297 41427
rect 1353 41371 1439 41427
rect 1495 41371 1581 41427
rect 1637 41371 1723 41427
rect 1779 41371 1865 41427
rect 1921 41371 2007 41427
rect 2063 41371 2149 41427
rect 2205 41371 2291 41427
rect 2347 41371 2433 41427
rect 2489 41371 2575 41427
rect 2631 41371 2717 41427
rect 2773 41371 2859 41427
rect 2915 41371 3001 41427
rect 3057 41371 3143 41427
rect 3199 41371 3285 41427
rect 3341 41371 3427 41427
rect 3483 41371 3569 41427
rect 3625 41371 3711 41427
rect 3767 41371 3853 41427
rect 3909 41371 3995 41427
rect 4051 41371 4137 41427
rect 4193 41371 4279 41427
rect 4335 41371 4421 41427
rect 4477 41371 4563 41427
rect 4619 41371 4705 41427
rect 4761 41371 4847 41427
rect 4903 41371 4989 41427
rect 5045 41371 5131 41427
rect 5187 41371 5273 41427
rect 5329 41371 5415 41427
rect 5471 41371 5557 41427
rect 5613 41371 5699 41427
rect 5755 41371 5841 41427
rect 5897 41371 5983 41427
rect 6039 41371 6125 41427
rect 6181 41371 6267 41427
rect 6323 41371 6409 41427
rect 6465 41371 6551 41427
rect 6607 41371 6693 41427
rect 6749 41371 6835 41427
rect 6891 41371 6977 41427
rect 7033 41371 7119 41427
rect 7175 41371 7261 41427
rect 7317 41371 7403 41427
rect 7459 41371 7545 41427
rect 7601 41371 7687 41427
rect 7743 41371 7829 41427
rect 7885 41371 7971 41427
rect 8027 41371 8113 41427
rect 8169 41371 8255 41427
rect 8311 41371 8397 41427
rect 8453 41371 8539 41427
rect 8595 41371 8681 41427
rect 8737 41371 8823 41427
rect 8879 41371 8965 41427
rect 9021 41371 9107 41427
rect 9163 41371 9249 41427
rect 9305 41371 9391 41427
rect 9447 41371 9533 41427
rect 9589 41371 9675 41427
rect 9731 41371 9817 41427
rect 9873 41371 9959 41427
rect 10015 41371 10101 41427
rect 10157 41371 10243 41427
rect 10299 41371 10385 41427
rect 10441 41371 10527 41427
rect 10583 41371 10669 41427
rect 10725 41371 10811 41427
rect 10867 41371 10953 41427
rect 11009 41371 11095 41427
rect 11151 41371 11237 41427
rect 11293 41371 11379 41427
rect 11435 41371 11521 41427
rect 11577 41371 11663 41427
rect 11719 41371 11805 41427
rect 11861 41371 11947 41427
rect 12003 41371 12089 41427
rect 12145 41371 12231 41427
rect 12287 41371 12373 41427
rect 12429 41371 12515 41427
rect 12571 41371 12657 41427
rect 12713 41371 12799 41427
rect 12855 41371 12941 41427
rect 12997 41371 13083 41427
rect 13139 41371 13225 41427
rect 13281 41371 13367 41427
rect 13423 41371 13509 41427
rect 13565 41371 13651 41427
rect 13707 41371 13793 41427
rect 13849 41371 13935 41427
rect 13991 41371 14077 41427
rect 14133 41371 14219 41427
rect 14275 41371 14361 41427
rect 14417 41371 14503 41427
rect 14559 41371 14645 41427
rect 14701 41371 14787 41427
rect 14843 41371 15000 41427
rect 0 41285 15000 41371
rect 0 41229 161 41285
rect 217 41229 303 41285
rect 359 41229 445 41285
rect 501 41229 587 41285
rect 643 41229 729 41285
rect 785 41229 871 41285
rect 927 41229 1013 41285
rect 1069 41229 1155 41285
rect 1211 41229 1297 41285
rect 1353 41229 1439 41285
rect 1495 41229 1581 41285
rect 1637 41229 1723 41285
rect 1779 41229 1865 41285
rect 1921 41229 2007 41285
rect 2063 41229 2149 41285
rect 2205 41229 2291 41285
rect 2347 41229 2433 41285
rect 2489 41229 2575 41285
rect 2631 41229 2717 41285
rect 2773 41229 2859 41285
rect 2915 41229 3001 41285
rect 3057 41229 3143 41285
rect 3199 41229 3285 41285
rect 3341 41229 3427 41285
rect 3483 41229 3569 41285
rect 3625 41229 3711 41285
rect 3767 41229 3853 41285
rect 3909 41229 3995 41285
rect 4051 41229 4137 41285
rect 4193 41229 4279 41285
rect 4335 41229 4421 41285
rect 4477 41229 4563 41285
rect 4619 41229 4705 41285
rect 4761 41229 4847 41285
rect 4903 41229 4989 41285
rect 5045 41229 5131 41285
rect 5187 41229 5273 41285
rect 5329 41229 5415 41285
rect 5471 41229 5557 41285
rect 5613 41229 5699 41285
rect 5755 41229 5841 41285
rect 5897 41229 5983 41285
rect 6039 41229 6125 41285
rect 6181 41229 6267 41285
rect 6323 41229 6409 41285
rect 6465 41229 6551 41285
rect 6607 41229 6693 41285
rect 6749 41229 6835 41285
rect 6891 41229 6977 41285
rect 7033 41229 7119 41285
rect 7175 41229 7261 41285
rect 7317 41229 7403 41285
rect 7459 41229 7545 41285
rect 7601 41229 7687 41285
rect 7743 41229 7829 41285
rect 7885 41229 7971 41285
rect 8027 41229 8113 41285
rect 8169 41229 8255 41285
rect 8311 41229 8397 41285
rect 8453 41229 8539 41285
rect 8595 41229 8681 41285
rect 8737 41229 8823 41285
rect 8879 41229 8965 41285
rect 9021 41229 9107 41285
rect 9163 41229 9249 41285
rect 9305 41229 9391 41285
rect 9447 41229 9533 41285
rect 9589 41229 9675 41285
rect 9731 41229 9817 41285
rect 9873 41229 9959 41285
rect 10015 41229 10101 41285
rect 10157 41229 10243 41285
rect 10299 41229 10385 41285
rect 10441 41229 10527 41285
rect 10583 41229 10669 41285
rect 10725 41229 10811 41285
rect 10867 41229 10953 41285
rect 11009 41229 11095 41285
rect 11151 41229 11237 41285
rect 11293 41229 11379 41285
rect 11435 41229 11521 41285
rect 11577 41229 11663 41285
rect 11719 41229 11805 41285
rect 11861 41229 11947 41285
rect 12003 41229 12089 41285
rect 12145 41229 12231 41285
rect 12287 41229 12373 41285
rect 12429 41229 12515 41285
rect 12571 41229 12657 41285
rect 12713 41229 12799 41285
rect 12855 41229 12941 41285
rect 12997 41229 13083 41285
rect 13139 41229 13225 41285
rect 13281 41229 13367 41285
rect 13423 41229 13509 41285
rect 13565 41229 13651 41285
rect 13707 41229 13793 41285
rect 13849 41229 13935 41285
rect 13991 41229 14077 41285
rect 14133 41229 14219 41285
rect 14275 41229 14361 41285
rect 14417 41229 14503 41285
rect 14559 41229 14645 41285
rect 14701 41229 14787 41285
rect 14843 41229 15000 41285
rect 0 41200 15000 41229
rect 0 40963 15000 41000
rect 0 40907 161 40963
rect 217 40907 303 40963
rect 359 40907 445 40963
rect 501 40907 587 40963
rect 643 40907 729 40963
rect 785 40907 871 40963
rect 927 40907 1013 40963
rect 1069 40907 1155 40963
rect 1211 40907 1297 40963
rect 1353 40907 1439 40963
rect 1495 40907 1581 40963
rect 1637 40907 1723 40963
rect 1779 40907 1865 40963
rect 1921 40907 2007 40963
rect 2063 40907 2149 40963
rect 2205 40907 2291 40963
rect 2347 40907 2433 40963
rect 2489 40907 2575 40963
rect 2631 40907 2717 40963
rect 2773 40907 2859 40963
rect 2915 40907 3001 40963
rect 3057 40907 3143 40963
rect 3199 40907 3285 40963
rect 3341 40907 3427 40963
rect 3483 40907 3569 40963
rect 3625 40907 3711 40963
rect 3767 40907 3853 40963
rect 3909 40907 3995 40963
rect 4051 40907 4137 40963
rect 4193 40907 4279 40963
rect 4335 40907 4421 40963
rect 4477 40907 4563 40963
rect 4619 40907 4705 40963
rect 4761 40907 4847 40963
rect 4903 40907 4989 40963
rect 5045 40907 5131 40963
rect 5187 40907 5273 40963
rect 5329 40907 5415 40963
rect 5471 40907 5557 40963
rect 5613 40907 5699 40963
rect 5755 40907 5841 40963
rect 5897 40907 5983 40963
rect 6039 40907 6125 40963
rect 6181 40907 6267 40963
rect 6323 40907 6409 40963
rect 6465 40907 6551 40963
rect 6607 40907 6693 40963
rect 6749 40907 6835 40963
rect 6891 40907 6977 40963
rect 7033 40907 7119 40963
rect 7175 40907 7261 40963
rect 7317 40907 7403 40963
rect 7459 40907 7545 40963
rect 7601 40907 7687 40963
rect 7743 40907 7829 40963
rect 7885 40907 7971 40963
rect 8027 40907 8113 40963
rect 8169 40907 8255 40963
rect 8311 40907 8397 40963
rect 8453 40907 8539 40963
rect 8595 40907 8681 40963
rect 8737 40907 8823 40963
rect 8879 40907 8965 40963
rect 9021 40907 9107 40963
rect 9163 40907 9249 40963
rect 9305 40907 9391 40963
rect 9447 40907 9533 40963
rect 9589 40907 9675 40963
rect 9731 40907 9817 40963
rect 9873 40907 9959 40963
rect 10015 40907 10101 40963
rect 10157 40907 10243 40963
rect 10299 40907 10385 40963
rect 10441 40907 10527 40963
rect 10583 40907 10669 40963
rect 10725 40907 10811 40963
rect 10867 40907 10953 40963
rect 11009 40907 11095 40963
rect 11151 40907 11237 40963
rect 11293 40907 11379 40963
rect 11435 40907 11521 40963
rect 11577 40907 11663 40963
rect 11719 40907 11805 40963
rect 11861 40907 11947 40963
rect 12003 40907 12089 40963
rect 12145 40907 12231 40963
rect 12287 40907 12373 40963
rect 12429 40907 12515 40963
rect 12571 40907 12657 40963
rect 12713 40907 12799 40963
rect 12855 40907 12941 40963
rect 12997 40907 13083 40963
rect 13139 40907 13225 40963
rect 13281 40907 13367 40963
rect 13423 40907 13509 40963
rect 13565 40907 13651 40963
rect 13707 40907 13793 40963
rect 13849 40907 13935 40963
rect 13991 40907 14077 40963
rect 14133 40907 14219 40963
rect 14275 40907 14361 40963
rect 14417 40907 14503 40963
rect 14559 40907 14645 40963
rect 14701 40907 14787 40963
rect 14843 40907 15000 40963
rect 0 40821 15000 40907
rect 0 40765 161 40821
rect 217 40765 303 40821
rect 359 40765 445 40821
rect 501 40765 587 40821
rect 643 40765 729 40821
rect 785 40765 871 40821
rect 927 40765 1013 40821
rect 1069 40765 1155 40821
rect 1211 40765 1297 40821
rect 1353 40765 1439 40821
rect 1495 40765 1581 40821
rect 1637 40765 1723 40821
rect 1779 40765 1865 40821
rect 1921 40765 2007 40821
rect 2063 40765 2149 40821
rect 2205 40765 2291 40821
rect 2347 40765 2433 40821
rect 2489 40765 2575 40821
rect 2631 40765 2717 40821
rect 2773 40765 2859 40821
rect 2915 40765 3001 40821
rect 3057 40765 3143 40821
rect 3199 40765 3285 40821
rect 3341 40765 3427 40821
rect 3483 40765 3569 40821
rect 3625 40765 3711 40821
rect 3767 40765 3853 40821
rect 3909 40765 3995 40821
rect 4051 40765 4137 40821
rect 4193 40765 4279 40821
rect 4335 40765 4421 40821
rect 4477 40765 4563 40821
rect 4619 40765 4705 40821
rect 4761 40765 4847 40821
rect 4903 40765 4989 40821
rect 5045 40765 5131 40821
rect 5187 40765 5273 40821
rect 5329 40765 5415 40821
rect 5471 40765 5557 40821
rect 5613 40765 5699 40821
rect 5755 40765 5841 40821
rect 5897 40765 5983 40821
rect 6039 40765 6125 40821
rect 6181 40765 6267 40821
rect 6323 40765 6409 40821
rect 6465 40765 6551 40821
rect 6607 40765 6693 40821
rect 6749 40765 6835 40821
rect 6891 40765 6977 40821
rect 7033 40765 7119 40821
rect 7175 40765 7261 40821
rect 7317 40765 7403 40821
rect 7459 40765 7545 40821
rect 7601 40765 7687 40821
rect 7743 40765 7829 40821
rect 7885 40765 7971 40821
rect 8027 40765 8113 40821
rect 8169 40765 8255 40821
rect 8311 40765 8397 40821
rect 8453 40765 8539 40821
rect 8595 40765 8681 40821
rect 8737 40765 8823 40821
rect 8879 40765 8965 40821
rect 9021 40765 9107 40821
rect 9163 40765 9249 40821
rect 9305 40765 9391 40821
rect 9447 40765 9533 40821
rect 9589 40765 9675 40821
rect 9731 40765 9817 40821
rect 9873 40765 9959 40821
rect 10015 40765 10101 40821
rect 10157 40765 10243 40821
rect 10299 40765 10385 40821
rect 10441 40765 10527 40821
rect 10583 40765 10669 40821
rect 10725 40765 10811 40821
rect 10867 40765 10953 40821
rect 11009 40765 11095 40821
rect 11151 40765 11237 40821
rect 11293 40765 11379 40821
rect 11435 40765 11521 40821
rect 11577 40765 11663 40821
rect 11719 40765 11805 40821
rect 11861 40765 11947 40821
rect 12003 40765 12089 40821
rect 12145 40765 12231 40821
rect 12287 40765 12373 40821
rect 12429 40765 12515 40821
rect 12571 40765 12657 40821
rect 12713 40765 12799 40821
rect 12855 40765 12941 40821
rect 12997 40765 13083 40821
rect 13139 40765 13225 40821
rect 13281 40765 13367 40821
rect 13423 40765 13509 40821
rect 13565 40765 13651 40821
rect 13707 40765 13793 40821
rect 13849 40765 13935 40821
rect 13991 40765 14077 40821
rect 14133 40765 14219 40821
rect 14275 40765 14361 40821
rect 14417 40765 14503 40821
rect 14559 40765 14645 40821
rect 14701 40765 14787 40821
rect 14843 40765 15000 40821
rect 0 40679 15000 40765
rect 0 40623 161 40679
rect 217 40623 303 40679
rect 359 40623 445 40679
rect 501 40623 587 40679
rect 643 40623 729 40679
rect 785 40623 871 40679
rect 927 40623 1013 40679
rect 1069 40623 1155 40679
rect 1211 40623 1297 40679
rect 1353 40623 1439 40679
rect 1495 40623 1581 40679
rect 1637 40623 1723 40679
rect 1779 40623 1865 40679
rect 1921 40623 2007 40679
rect 2063 40623 2149 40679
rect 2205 40623 2291 40679
rect 2347 40623 2433 40679
rect 2489 40623 2575 40679
rect 2631 40623 2717 40679
rect 2773 40623 2859 40679
rect 2915 40623 3001 40679
rect 3057 40623 3143 40679
rect 3199 40623 3285 40679
rect 3341 40623 3427 40679
rect 3483 40623 3569 40679
rect 3625 40623 3711 40679
rect 3767 40623 3853 40679
rect 3909 40623 3995 40679
rect 4051 40623 4137 40679
rect 4193 40623 4279 40679
rect 4335 40623 4421 40679
rect 4477 40623 4563 40679
rect 4619 40623 4705 40679
rect 4761 40623 4847 40679
rect 4903 40623 4989 40679
rect 5045 40623 5131 40679
rect 5187 40623 5273 40679
rect 5329 40623 5415 40679
rect 5471 40623 5557 40679
rect 5613 40623 5699 40679
rect 5755 40623 5841 40679
rect 5897 40623 5983 40679
rect 6039 40623 6125 40679
rect 6181 40623 6267 40679
rect 6323 40623 6409 40679
rect 6465 40623 6551 40679
rect 6607 40623 6693 40679
rect 6749 40623 6835 40679
rect 6891 40623 6977 40679
rect 7033 40623 7119 40679
rect 7175 40623 7261 40679
rect 7317 40623 7403 40679
rect 7459 40623 7545 40679
rect 7601 40623 7687 40679
rect 7743 40623 7829 40679
rect 7885 40623 7971 40679
rect 8027 40623 8113 40679
rect 8169 40623 8255 40679
rect 8311 40623 8397 40679
rect 8453 40623 8539 40679
rect 8595 40623 8681 40679
rect 8737 40623 8823 40679
rect 8879 40623 8965 40679
rect 9021 40623 9107 40679
rect 9163 40623 9249 40679
rect 9305 40623 9391 40679
rect 9447 40623 9533 40679
rect 9589 40623 9675 40679
rect 9731 40623 9817 40679
rect 9873 40623 9959 40679
rect 10015 40623 10101 40679
rect 10157 40623 10243 40679
rect 10299 40623 10385 40679
rect 10441 40623 10527 40679
rect 10583 40623 10669 40679
rect 10725 40623 10811 40679
rect 10867 40623 10953 40679
rect 11009 40623 11095 40679
rect 11151 40623 11237 40679
rect 11293 40623 11379 40679
rect 11435 40623 11521 40679
rect 11577 40623 11663 40679
rect 11719 40623 11805 40679
rect 11861 40623 11947 40679
rect 12003 40623 12089 40679
rect 12145 40623 12231 40679
rect 12287 40623 12373 40679
rect 12429 40623 12515 40679
rect 12571 40623 12657 40679
rect 12713 40623 12799 40679
rect 12855 40623 12941 40679
rect 12997 40623 13083 40679
rect 13139 40623 13225 40679
rect 13281 40623 13367 40679
rect 13423 40623 13509 40679
rect 13565 40623 13651 40679
rect 13707 40623 13793 40679
rect 13849 40623 13935 40679
rect 13991 40623 14077 40679
rect 14133 40623 14219 40679
rect 14275 40623 14361 40679
rect 14417 40623 14503 40679
rect 14559 40623 14645 40679
rect 14701 40623 14787 40679
rect 14843 40623 15000 40679
rect 0 40537 15000 40623
rect 0 40481 161 40537
rect 217 40481 303 40537
rect 359 40481 445 40537
rect 501 40481 587 40537
rect 643 40481 729 40537
rect 785 40481 871 40537
rect 927 40481 1013 40537
rect 1069 40481 1155 40537
rect 1211 40481 1297 40537
rect 1353 40481 1439 40537
rect 1495 40481 1581 40537
rect 1637 40481 1723 40537
rect 1779 40481 1865 40537
rect 1921 40481 2007 40537
rect 2063 40481 2149 40537
rect 2205 40481 2291 40537
rect 2347 40481 2433 40537
rect 2489 40481 2575 40537
rect 2631 40481 2717 40537
rect 2773 40481 2859 40537
rect 2915 40481 3001 40537
rect 3057 40481 3143 40537
rect 3199 40481 3285 40537
rect 3341 40481 3427 40537
rect 3483 40481 3569 40537
rect 3625 40481 3711 40537
rect 3767 40481 3853 40537
rect 3909 40481 3995 40537
rect 4051 40481 4137 40537
rect 4193 40481 4279 40537
rect 4335 40481 4421 40537
rect 4477 40481 4563 40537
rect 4619 40481 4705 40537
rect 4761 40481 4847 40537
rect 4903 40481 4989 40537
rect 5045 40481 5131 40537
rect 5187 40481 5273 40537
rect 5329 40481 5415 40537
rect 5471 40481 5557 40537
rect 5613 40481 5699 40537
rect 5755 40481 5841 40537
rect 5897 40481 5983 40537
rect 6039 40481 6125 40537
rect 6181 40481 6267 40537
rect 6323 40481 6409 40537
rect 6465 40481 6551 40537
rect 6607 40481 6693 40537
rect 6749 40481 6835 40537
rect 6891 40481 6977 40537
rect 7033 40481 7119 40537
rect 7175 40481 7261 40537
rect 7317 40481 7403 40537
rect 7459 40481 7545 40537
rect 7601 40481 7687 40537
rect 7743 40481 7829 40537
rect 7885 40481 7971 40537
rect 8027 40481 8113 40537
rect 8169 40481 8255 40537
rect 8311 40481 8397 40537
rect 8453 40481 8539 40537
rect 8595 40481 8681 40537
rect 8737 40481 8823 40537
rect 8879 40481 8965 40537
rect 9021 40481 9107 40537
rect 9163 40481 9249 40537
rect 9305 40481 9391 40537
rect 9447 40481 9533 40537
rect 9589 40481 9675 40537
rect 9731 40481 9817 40537
rect 9873 40481 9959 40537
rect 10015 40481 10101 40537
rect 10157 40481 10243 40537
rect 10299 40481 10385 40537
rect 10441 40481 10527 40537
rect 10583 40481 10669 40537
rect 10725 40481 10811 40537
rect 10867 40481 10953 40537
rect 11009 40481 11095 40537
rect 11151 40481 11237 40537
rect 11293 40481 11379 40537
rect 11435 40481 11521 40537
rect 11577 40481 11663 40537
rect 11719 40481 11805 40537
rect 11861 40481 11947 40537
rect 12003 40481 12089 40537
rect 12145 40481 12231 40537
rect 12287 40481 12373 40537
rect 12429 40481 12515 40537
rect 12571 40481 12657 40537
rect 12713 40481 12799 40537
rect 12855 40481 12941 40537
rect 12997 40481 13083 40537
rect 13139 40481 13225 40537
rect 13281 40481 13367 40537
rect 13423 40481 13509 40537
rect 13565 40481 13651 40537
rect 13707 40481 13793 40537
rect 13849 40481 13935 40537
rect 13991 40481 14077 40537
rect 14133 40481 14219 40537
rect 14275 40481 14361 40537
rect 14417 40481 14503 40537
rect 14559 40481 14645 40537
rect 14701 40481 14787 40537
rect 14843 40481 15000 40537
rect 0 40395 15000 40481
rect 0 40339 161 40395
rect 217 40339 303 40395
rect 359 40339 445 40395
rect 501 40339 587 40395
rect 643 40339 729 40395
rect 785 40339 871 40395
rect 927 40339 1013 40395
rect 1069 40339 1155 40395
rect 1211 40339 1297 40395
rect 1353 40339 1439 40395
rect 1495 40339 1581 40395
rect 1637 40339 1723 40395
rect 1779 40339 1865 40395
rect 1921 40339 2007 40395
rect 2063 40339 2149 40395
rect 2205 40339 2291 40395
rect 2347 40339 2433 40395
rect 2489 40339 2575 40395
rect 2631 40339 2717 40395
rect 2773 40339 2859 40395
rect 2915 40339 3001 40395
rect 3057 40339 3143 40395
rect 3199 40339 3285 40395
rect 3341 40339 3427 40395
rect 3483 40339 3569 40395
rect 3625 40339 3711 40395
rect 3767 40339 3853 40395
rect 3909 40339 3995 40395
rect 4051 40339 4137 40395
rect 4193 40339 4279 40395
rect 4335 40339 4421 40395
rect 4477 40339 4563 40395
rect 4619 40339 4705 40395
rect 4761 40339 4847 40395
rect 4903 40339 4989 40395
rect 5045 40339 5131 40395
rect 5187 40339 5273 40395
rect 5329 40339 5415 40395
rect 5471 40339 5557 40395
rect 5613 40339 5699 40395
rect 5755 40339 5841 40395
rect 5897 40339 5983 40395
rect 6039 40339 6125 40395
rect 6181 40339 6267 40395
rect 6323 40339 6409 40395
rect 6465 40339 6551 40395
rect 6607 40339 6693 40395
rect 6749 40339 6835 40395
rect 6891 40339 6977 40395
rect 7033 40339 7119 40395
rect 7175 40339 7261 40395
rect 7317 40339 7403 40395
rect 7459 40339 7545 40395
rect 7601 40339 7687 40395
rect 7743 40339 7829 40395
rect 7885 40339 7971 40395
rect 8027 40339 8113 40395
rect 8169 40339 8255 40395
rect 8311 40339 8397 40395
rect 8453 40339 8539 40395
rect 8595 40339 8681 40395
rect 8737 40339 8823 40395
rect 8879 40339 8965 40395
rect 9021 40339 9107 40395
rect 9163 40339 9249 40395
rect 9305 40339 9391 40395
rect 9447 40339 9533 40395
rect 9589 40339 9675 40395
rect 9731 40339 9817 40395
rect 9873 40339 9959 40395
rect 10015 40339 10101 40395
rect 10157 40339 10243 40395
rect 10299 40339 10385 40395
rect 10441 40339 10527 40395
rect 10583 40339 10669 40395
rect 10725 40339 10811 40395
rect 10867 40339 10953 40395
rect 11009 40339 11095 40395
rect 11151 40339 11237 40395
rect 11293 40339 11379 40395
rect 11435 40339 11521 40395
rect 11577 40339 11663 40395
rect 11719 40339 11805 40395
rect 11861 40339 11947 40395
rect 12003 40339 12089 40395
rect 12145 40339 12231 40395
rect 12287 40339 12373 40395
rect 12429 40339 12515 40395
rect 12571 40339 12657 40395
rect 12713 40339 12799 40395
rect 12855 40339 12941 40395
rect 12997 40339 13083 40395
rect 13139 40339 13225 40395
rect 13281 40339 13367 40395
rect 13423 40339 13509 40395
rect 13565 40339 13651 40395
rect 13707 40339 13793 40395
rect 13849 40339 13935 40395
rect 13991 40339 14077 40395
rect 14133 40339 14219 40395
rect 14275 40339 14361 40395
rect 14417 40339 14503 40395
rect 14559 40339 14645 40395
rect 14701 40339 14787 40395
rect 14843 40339 15000 40395
rect 0 40253 15000 40339
rect 0 40197 161 40253
rect 217 40197 303 40253
rect 359 40197 445 40253
rect 501 40197 587 40253
rect 643 40197 729 40253
rect 785 40197 871 40253
rect 927 40197 1013 40253
rect 1069 40197 1155 40253
rect 1211 40197 1297 40253
rect 1353 40197 1439 40253
rect 1495 40197 1581 40253
rect 1637 40197 1723 40253
rect 1779 40197 1865 40253
rect 1921 40197 2007 40253
rect 2063 40197 2149 40253
rect 2205 40197 2291 40253
rect 2347 40197 2433 40253
rect 2489 40197 2575 40253
rect 2631 40197 2717 40253
rect 2773 40197 2859 40253
rect 2915 40197 3001 40253
rect 3057 40197 3143 40253
rect 3199 40197 3285 40253
rect 3341 40197 3427 40253
rect 3483 40197 3569 40253
rect 3625 40197 3711 40253
rect 3767 40197 3853 40253
rect 3909 40197 3995 40253
rect 4051 40197 4137 40253
rect 4193 40197 4279 40253
rect 4335 40197 4421 40253
rect 4477 40197 4563 40253
rect 4619 40197 4705 40253
rect 4761 40197 4847 40253
rect 4903 40197 4989 40253
rect 5045 40197 5131 40253
rect 5187 40197 5273 40253
rect 5329 40197 5415 40253
rect 5471 40197 5557 40253
rect 5613 40197 5699 40253
rect 5755 40197 5841 40253
rect 5897 40197 5983 40253
rect 6039 40197 6125 40253
rect 6181 40197 6267 40253
rect 6323 40197 6409 40253
rect 6465 40197 6551 40253
rect 6607 40197 6693 40253
rect 6749 40197 6835 40253
rect 6891 40197 6977 40253
rect 7033 40197 7119 40253
rect 7175 40197 7261 40253
rect 7317 40197 7403 40253
rect 7459 40197 7545 40253
rect 7601 40197 7687 40253
rect 7743 40197 7829 40253
rect 7885 40197 7971 40253
rect 8027 40197 8113 40253
rect 8169 40197 8255 40253
rect 8311 40197 8397 40253
rect 8453 40197 8539 40253
rect 8595 40197 8681 40253
rect 8737 40197 8823 40253
rect 8879 40197 8965 40253
rect 9021 40197 9107 40253
rect 9163 40197 9249 40253
rect 9305 40197 9391 40253
rect 9447 40197 9533 40253
rect 9589 40197 9675 40253
rect 9731 40197 9817 40253
rect 9873 40197 9959 40253
rect 10015 40197 10101 40253
rect 10157 40197 10243 40253
rect 10299 40197 10385 40253
rect 10441 40197 10527 40253
rect 10583 40197 10669 40253
rect 10725 40197 10811 40253
rect 10867 40197 10953 40253
rect 11009 40197 11095 40253
rect 11151 40197 11237 40253
rect 11293 40197 11379 40253
rect 11435 40197 11521 40253
rect 11577 40197 11663 40253
rect 11719 40197 11805 40253
rect 11861 40197 11947 40253
rect 12003 40197 12089 40253
rect 12145 40197 12231 40253
rect 12287 40197 12373 40253
rect 12429 40197 12515 40253
rect 12571 40197 12657 40253
rect 12713 40197 12799 40253
rect 12855 40197 12941 40253
rect 12997 40197 13083 40253
rect 13139 40197 13225 40253
rect 13281 40197 13367 40253
rect 13423 40197 13509 40253
rect 13565 40197 13651 40253
rect 13707 40197 13793 40253
rect 13849 40197 13935 40253
rect 13991 40197 14077 40253
rect 14133 40197 14219 40253
rect 14275 40197 14361 40253
rect 14417 40197 14503 40253
rect 14559 40197 14645 40253
rect 14701 40197 14787 40253
rect 14843 40197 15000 40253
rect 0 40111 15000 40197
rect 0 40055 161 40111
rect 217 40055 303 40111
rect 359 40055 445 40111
rect 501 40055 587 40111
rect 643 40055 729 40111
rect 785 40055 871 40111
rect 927 40055 1013 40111
rect 1069 40055 1155 40111
rect 1211 40055 1297 40111
rect 1353 40055 1439 40111
rect 1495 40055 1581 40111
rect 1637 40055 1723 40111
rect 1779 40055 1865 40111
rect 1921 40055 2007 40111
rect 2063 40055 2149 40111
rect 2205 40055 2291 40111
rect 2347 40055 2433 40111
rect 2489 40055 2575 40111
rect 2631 40055 2717 40111
rect 2773 40055 2859 40111
rect 2915 40055 3001 40111
rect 3057 40055 3143 40111
rect 3199 40055 3285 40111
rect 3341 40055 3427 40111
rect 3483 40055 3569 40111
rect 3625 40055 3711 40111
rect 3767 40055 3853 40111
rect 3909 40055 3995 40111
rect 4051 40055 4137 40111
rect 4193 40055 4279 40111
rect 4335 40055 4421 40111
rect 4477 40055 4563 40111
rect 4619 40055 4705 40111
rect 4761 40055 4847 40111
rect 4903 40055 4989 40111
rect 5045 40055 5131 40111
rect 5187 40055 5273 40111
rect 5329 40055 5415 40111
rect 5471 40055 5557 40111
rect 5613 40055 5699 40111
rect 5755 40055 5841 40111
rect 5897 40055 5983 40111
rect 6039 40055 6125 40111
rect 6181 40055 6267 40111
rect 6323 40055 6409 40111
rect 6465 40055 6551 40111
rect 6607 40055 6693 40111
rect 6749 40055 6835 40111
rect 6891 40055 6977 40111
rect 7033 40055 7119 40111
rect 7175 40055 7261 40111
rect 7317 40055 7403 40111
rect 7459 40055 7545 40111
rect 7601 40055 7687 40111
rect 7743 40055 7829 40111
rect 7885 40055 7971 40111
rect 8027 40055 8113 40111
rect 8169 40055 8255 40111
rect 8311 40055 8397 40111
rect 8453 40055 8539 40111
rect 8595 40055 8681 40111
rect 8737 40055 8823 40111
rect 8879 40055 8965 40111
rect 9021 40055 9107 40111
rect 9163 40055 9249 40111
rect 9305 40055 9391 40111
rect 9447 40055 9533 40111
rect 9589 40055 9675 40111
rect 9731 40055 9817 40111
rect 9873 40055 9959 40111
rect 10015 40055 10101 40111
rect 10157 40055 10243 40111
rect 10299 40055 10385 40111
rect 10441 40055 10527 40111
rect 10583 40055 10669 40111
rect 10725 40055 10811 40111
rect 10867 40055 10953 40111
rect 11009 40055 11095 40111
rect 11151 40055 11237 40111
rect 11293 40055 11379 40111
rect 11435 40055 11521 40111
rect 11577 40055 11663 40111
rect 11719 40055 11805 40111
rect 11861 40055 11947 40111
rect 12003 40055 12089 40111
rect 12145 40055 12231 40111
rect 12287 40055 12373 40111
rect 12429 40055 12515 40111
rect 12571 40055 12657 40111
rect 12713 40055 12799 40111
rect 12855 40055 12941 40111
rect 12997 40055 13083 40111
rect 13139 40055 13225 40111
rect 13281 40055 13367 40111
rect 13423 40055 13509 40111
rect 13565 40055 13651 40111
rect 13707 40055 13793 40111
rect 13849 40055 13935 40111
rect 13991 40055 14077 40111
rect 14133 40055 14219 40111
rect 14275 40055 14361 40111
rect 14417 40055 14503 40111
rect 14559 40055 14645 40111
rect 14701 40055 14787 40111
rect 14843 40055 15000 40111
rect 0 39969 15000 40055
rect 0 39913 161 39969
rect 217 39913 303 39969
rect 359 39913 445 39969
rect 501 39913 587 39969
rect 643 39913 729 39969
rect 785 39913 871 39969
rect 927 39913 1013 39969
rect 1069 39913 1155 39969
rect 1211 39913 1297 39969
rect 1353 39913 1439 39969
rect 1495 39913 1581 39969
rect 1637 39913 1723 39969
rect 1779 39913 1865 39969
rect 1921 39913 2007 39969
rect 2063 39913 2149 39969
rect 2205 39913 2291 39969
rect 2347 39913 2433 39969
rect 2489 39913 2575 39969
rect 2631 39913 2717 39969
rect 2773 39913 2859 39969
rect 2915 39913 3001 39969
rect 3057 39913 3143 39969
rect 3199 39913 3285 39969
rect 3341 39913 3427 39969
rect 3483 39913 3569 39969
rect 3625 39913 3711 39969
rect 3767 39913 3853 39969
rect 3909 39913 3995 39969
rect 4051 39913 4137 39969
rect 4193 39913 4279 39969
rect 4335 39913 4421 39969
rect 4477 39913 4563 39969
rect 4619 39913 4705 39969
rect 4761 39913 4847 39969
rect 4903 39913 4989 39969
rect 5045 39913 5131 39969
rect 5187 39913 5273 39969
rect 5329 39913 5415 39969
rect 5471 39913 5557 39969
rect 5613 39913 5699 39969
rect 5755 39913 5841 39969
rect 5897 39913 5983 39969
rect 6039 39913 6125 39969
rect 6181 39913 6267 39969
rect 6323 39913 6409 39969
rect 6465 39913 6551 39969
rect 6607 39913 6693 39969
rect 6749 39913 6835 39969
rect 6891 39913 6977 39969
rect 7033 39913 7119 39969
rect 7175 39913 7261 39969
rect 7317 39913 7403 39969
rect 7459 39913 7545 39969
rect 7601 39913 7687 39969
rect 7743 39913 7829 39969
rect 7885 39913 7971 39969
rect 8027 39913 8113 39969
rect 8169 39913 8255 39969
rect 8311 39913 8397 39969
rect 8453 39913 8539 39969
rect 8595 39913 8681 39969
rect 8737 39913 8823 39969
rect 8879 39913 8965 39969
rect 9021 39913 9107 39969
rect 9163 39913 9249 39969
rect 9305 39913 9391 39969
rect 9447 39913 9533 39969
rect 9589 39913 9675 39969
rect 9731 39913 9817 39969
rect 9873 39913 9959 39969
rect 10015 39913 10101 39969
rect 10157 39913 10243 39969
rect 10299 39913 10385 39969
rect 10441 39913 10527 39969
rect 10583 39913 10669 39969
rect 10725 39913 10811 39969
rect 10867 39913 10953 39969
rect 11009 39913 11095 39969
rect 11151 39913 11237 39969
rect 11293 39913 11379 39969
rect 11435 39913 11521 39969
rect 11577 39913 11663 39969
rect 11719 39913 11805 39969
rect 11861 39913 11947 39969
rect 12003 39913 12089 39969
rect 12145 39913 12231 39969
rect 12287 39913 12373 39969
rect 12429 39913 12515 39969
rect 12571 39913 12657 39969
rect 12713 39913 12799 39969
rect 12855 39913 12941 39969
rect 12997 39913 13083 39969
rect 13139 39913 13225 39969
rect 13281 39913 13367 39969
rect 13423 39913 13509 39969
rect 13565 39913 13651 39969
rect 13707 39913 13793 39969
rect 13849 39913 13935 39969
rect 13991 39913 14077 39969
rect 14133 39913 14219 39969
rect 14275 39913 14361 39969
rect 14417 39913 14503 39969
rect 14559 39913 14645 39969
rect 14701 39913 14787 39969
rect 14843 39913 15000 39969
rect 0 39827 15000 39913
rect 0 39771 161 39827
rect 217 39771 303 39827
rect 359 39771 445 39827
rect 501 39771 587 39827
rect 643 39771 729 39827
rect 785 39771 871 39827
rect 927 39771 1013 39827
rect 1069 39771 1155 39827
rect 1211 39771 1297 39827
rect 1353 39771 1439 39827
rect 1495 39771 1581 39827
rect 1637 39771 1723 39827
rect 1779 39771 1865 39827
rect 1921 39771 2007 39827
rect 2063 39771 2149 39827
rect 2205 39771 2291 39827
rect 2347 39771 2433 39827
rect 2489 39771 2575 39827
rect 2631 39771 2717 39827
rect 2773 39771 2859 39827
rect 2915 39771 3001 39827
rect 3057 39771 3143 39827
rect 3199 39771 3285 39827
rect 3341 39771 3427 39827
rect 3483 39771 3569 39827
rect 3625 39771 3711 39827
rect 3767 39771 3853 39827
rect 3909 39771 3995 39827
rect 4051 39771 4137 39827
rect 4193 39771 4279 39827
rect 4335 39771 4421 39827
rect 4477 39771 4563 39827
rect 4619 39771 4705 39827
rect 4761 39771 4847 39827
rect 4903 39771 4989 39827
rect 5045 39771 5131 39827
rect 5187 39771 5273 39827
rect 5329 39771 5415 39827
rect 5471 39771 5557 39827
rect 5613 39771 5699 39827
rect 5755 39771 5841 39827
rect 5897 39771 5983 39827
rect 6039 39771 6125 39827
rect 6181 39771 6267 39827
rect 6323 39771 6409 39827
rect 6465 39771 6551 39827
rect 6607 39771 6693 39827
rect 6749 39771 6835 39827
rect 6891 39771 6977 39827
rect 7033 39771 7119 39827
rect 7175 39771 7261 39827
rect 7317 39771 7403 39827
rect 7459 39771 7545 39827
rect 7601 39771 7687 39827
rect 7743 39771 7829 39827
rect 7885 39771 7971 39827
rect 8027 39771 8113 39827
rect 8169 39771 8255 39827
rect 8311 39771 8397 39827
rect 8453 39771 8539 39827
rect 8595 39771 8681 39827
rect 8737 39771 8823 39827
rect 8879 39771 8965 39827
rect 9021 39771 9107 39827
rect 9163 39771 9249 39827
rect 9305 39771 9391 39827
rect 9447 39771 9533 39827
rect 9589 39771 9675 39827
rect 9731 39771 9817 39827
rect 9873 39771 9959 39827
rect 10015 39771 10101 39827
rect 10157 39771 10243 39827
rect 10299 39771 10385 39827
rect 10441 39771 10527 39827
rect 10583 39771 10669 39827
rect 10725 39771 10811 39827
rect 10867 39771 10953 39827
rect 11009 39771 11095 39827
rect 11151 39771 11237 39827
rect 11293 39771 11379 39827
rect 11435 39771 11521 39827
rect 11577 39771 11663 39827
rect 11719 39771 11805 39827
rect 11861 39771 11947 39827
rect 12003 39771 12089 39827
rect 12145 39771 12231 39827
rect 12287 39771 12373 39827
rect 12429 39771 12515 39827
rect 12571 39771 12657 39827
rect 12713 39771 12799 39827
rect 12855 39771 12941 39827
rect 12997 39771 13083 39827
rect 13139 39771 13225 39827
rect 13281 39771 13367 39827
rect 13423 39771 13509 39827
rect 13565 39771 13651 39827
rect 13707 39771 13793 39827
rect 13849 39771 13935 39827
rect 13991 39771 14077 39827
rect 14133 39771 14219 39827
rect 14275 39771 14361 39827
rect 14417 39771 14503 39827
rect 14559 39771 14645 39827
rect 14701 39771 14787 39827
rect 14843 39771 15000 39827
rect 0 39685 15000 39771
rect 0 39629 161 39685
rect 217 39629 303 39685
rect 359 39629 445 39685
rect 501 39629 587 39685
rect 643 39629 729 39685
rect 785 39629 871 39685
rect 927 39629 1013 39685
rect 1069 39629 1155 39685
rect 1211 39629 1297 39685
rect 1353 39629 1439 39685
rect 1495 39629 1581 39685
rect 1637 39629 1723 39685
rect 1779 39629 1865 39685
rect 1921 39629 2007 39685
rect 2063 39629 2149 39685
rect 2205 39629 2291 39685
rect 2347 39629 2433 39685
rect 2489 39629 2575 39685
rect 2631 39629 2717 39685
rect 2773 39629 2859 39685
rect 2915 39629 3001 39685
rect 3057 39629 3143 39685
rect 3199 39629 3285 39685
rect 3341 39629 3427 39685
rect 3483 39629 3569 39685
rect 3625 39629 3711 39685
rect 3767 39629 3853 39685
rect 3909 39629 3995 39685
rect 4051 39629 4137 39685
rect 4193 39629 4279 39685
rect 4335 39629 4421 39685
rect 4477 39629 4563 39685
rect 4619 39629 4705 39685
rect 4761 39629 4847 39685
rect 4903 39629 4989 39685
rect 5045 39629 5131 39685
rect 5187 39629 5273 39685
rect 5329 39629 5415 39685
rect 5471 39629 5557 39685
rect 5613 39629 5699 39685
rect 5755 39629 5841 39685
rect 5897 39629 5983 39685
rect 6039 39629 6125 39685
rect 6181 39629 6267 39685
rect 6323 39629 6409 39685
rect 6465 39629 6551 39685
rect 6607 39629 6693 39685
rect 6749 39629 6835 39685
rect 6891 39629 6977 39685
rect 7033 39629 7119 39685
rect 7175 39629 7261 39685
rect 7317 39629 7403 39685
rect 7459 39629 7545 39685
rect 7601 39629 7687 39685
rect 7743 39629 7829 39685
rect 7885 39629 7971 39685
rect 8027 39629 8113 39685
rect 8169 39629 8255 39685
rect 8311 39629 8397 39685
rect 8453 39629 8539 39685
rect 8595 39629 8681 39685
rect 8737 39629 8823 39685
rect 8879 39629 8965 39685
rect 9021 39629 9107 39685
rect 9163 39629 9249 39685
rect 9305 39629 9391 39685
rect 9447 39629 9533 39685
rect 9589 39629 9675 39685
rect 9731 39629 9817 39685
rect 9873 39629 9959 39685
rect 10015 39629 10101 39685
rect 10157 39629 10243 39685
rect 10299 39629 10385 39685
rect 10441 39629 10527 39685
rect 10583 39629 10669 39685
rect 10725 39629 10811 39685
rect 10867 39629 10953 39685
rect 11009 39629 11095 39685
rect 11151 39629 11237 39685
rect 11293 39629 11379 39685
rect 11435 39629 11521 39685
rect 11577 39629 11663 39685
rect 11719 39629 11805 39685
rect 11861 39629 11947 39685
rect 12003 39629 12089 39685
rect 12145 39629 12231 39685
rect 12287 39629 12373 39685
rect 12429 39629 12515 39685
rect 12571 39629 12657 39685
rect 12713 39629 12799 39685
rect 12855 39629 12941 39685
rect 12997 39629 13083 39685
rect 13139 39629 13225 39685
rect 13281 39629 13367 39685
rect 13423 39629 13509 39685
rect 13565 39629 13651 39685
rect 13707 39629 13793 39685
rect 13849 39629 13935 39685
rect 13991 39629 14077 39685
rect 14133 39629 14219 39685
rect 14275 39629 14361 39685
rect 14417 39629 14503 39685
rect 14559 39629 14645 39685
rect 14701 39629 14787 39685
rect 14843 39629 15000 39685
rect 0 39600 15000 39629
rect 0 39342 15000 39400
rect 0 39286 161 39342
rect 217 39286 303 39342
rect 359 39286 445 39342
rect 501 39286 587 39342
rect 643 39286 729 39342
rect 785 39286 871 39342
rect 927 39286 1013 39342
rect 1069 39286 1155 39342
rect 1211 39286 1297 39342
rect 1353 39286 1439 39342
rect 1495 39286 1581 39342
rect 1637 39286 1723 39342
rect 1779 39286 1865 39342
rect 1921 39286 2007 39342
rect 2063 39286 2149 39342
rect 2205 39286 2291 39342
rect 2347 39286 2433 39342
rect 2489 39286 2575 39342
rect 2631 39286 2717 39342
rect 2773 39286 2859 39342
rect 2915 39286 3001 39342
rect 3057 39286 3143 39342
rect 3199 39286 3285 39342
rect 3341 39286 3427 39342
rect 3483 39286 3569 39342
rect 3625 39286 3711 39342
rect 3767 39286 3853 39342
rect 3909 39286 3995 39342
rect 4051 39286 4137 39342
rect 4193 39286 4279 39342
rect 4335 39286 4421 39342
rect 4477 39286 4563 39342
rect 4619 39286 4705 39342
rect 4761 39286 4847 39342
rect 4903 39286 4989 39342
rect 5045 39286 5131 39342
rect 5187 39286 5273 39342
rect 5329 39286 5415 39342
rect 5471 39286 5557 39342
rect 5613 39286 5699 39342
rect 5755 39286 5841 39342
rect 5897 39286 5983 39342
rect 6039 39286 6125 39342
rect 6181 39286 6267 39342
rect 6323 39286 6409 39342
rect 6465 39286 6551 39342
rect 6607 39286 6693 39342
rect 6749 39286 6835 39342
rect 6891 39286 6977 39342
rect 7033 39286 7119 39342
rect 7175 39286 7261 39342
rect 7317 39286 7403 39342
rect 7459 39286 7545 39342
rect 7601 39286 7687 39342
rect 7743 39286 7829 39342
rect 7885 39286 7971 39342
rect 8027 39286 8113 39342
rect 8169 39286 8255 39342
rect 8311 39286 8397 39342
rect 8453 39286 8539 39342
rect 8595 39286 8681 39342
rect 8737 39286 8823 39342
rect 8879 39286 8965 39342
rect 9021 39286 9107 39342
rect 9163 39286 9249 39342
rect 9305 39286 9391 39342
rect 9447 39286 9533 39342
rect 9589 39286 9675 39342
rect 9731 39286 9817 39342
rect 9873 39286 9959 39342
rect 10015 39286 10101 39342
rect 10157 39286 10243 39342
rect 10299 39286 10385 39342
rect 10441 39286 10527 39342
rect 10583 39286 10669 39342
rect 10725 39286 10811 39342
rect 10867 39286 10953 39342
rect 11009 39286 11095 39342
rect 11151 39286 11237 39342
rect 11293 39286 11379 39342
rect 11435 39286 11521 39342
rect 11577 39286 11663 39342
rect 11719 39286 11805 39342
rect 11861 39286 11947 39342
rect 12003 39286 12089 39342
rect 12145 39286 12231 39342
rect 12287 39286 12373 39342
rect 12429 39286 12515 39342
rect 12571 39286 12657 39342
rect 12713 39286 12799 39342
rect 12855 39286 12941 39342
rect 12997 39286 13083 39342
rect 13139 39286 13225 39342
rect 13281 39286 13367 39342
rect 13423 39286 13509 39342
rect 13565 39286 13651 39342
rect 13707 39286 13793 39342
rect 13849 39286 13935 39342
rect 13991 39286 14077 39342
rect 14133 39286 14219 39342
rect 14275 39286 14361 39342
rect 14417 39286 14503 39342
rect 14559 39286 14645 39342
rect 14701 39286 14787 39342
rect 14843 39286 15000 39342
rect 0 39200 15000 39286
rect 0 39144 161 39200
rect 217 39144 303 39200
rect 359 39144 445 39200
rect 501 39144 587 39200
rect 643 39144 729 39200
rect 785 39144 871 39200
rect 927 39144 1013 39200
rect 1069 39144 1155 39200
rect 1211 39144 1297 39200
rect 1353 39144 1439 39200
rect 1495 39144 1581 39200
rect 1637 39144 1723 39200
rect 1779 39144 1865 39200
rect 1921 39144 2007 39200
rect 2063 39144 2149 39200
rect 2205 39144 2291 39200
rect 2347 39144 2433 39200
rect 2489 39144 2575 39200
rect 2631 39144 2717 39200
rect 2773 39144 2859 39200
rect 2915 39144 3001 39200
rect 3057 39144 3143 39200
rect 3199 39144 3285 39200
rect 3341 39144 3427 39200
rect 3483 39144 3569 39200
rect 3625 39144 3711 39200
rect 3767 39144 3853 39200
rect 3909 39144 3995 39200
rect 4051 39144 4137 39200
rect 4193 39144 4279 39200
rect 4335 39144 4421 39200
rect 4477 39144 4563 39200
rect 4619 39144 4705 39200
rect 4761 39144 4847 39200
rect 4903 39144 4989 39200
rect 5045 39144 5131 39200
rect 5187 39144 5273 39200
rect 5329 39144 5415 39200
rect 5471 39144 5557 39200
rect 5613 39144 5699 39200
rect 5755 39144 5841 39200
rect 5897 39144 5983 39200
rect 6039 39144 6125 39200
rect 6181 39144 6267 39200
rect 6323 39144 6409 39200
rect 6465 39144 6551 39200
rect 6607 39144 6693 39200
rect 6749 39144 6835 39200
rect 6891 39144 6977 39200
rect 7033 39144 7119 39200
rect 7175 39144 7261 39200
rect 7317 39144 7403 39200
rect 7459 39144 7545 39200
rect 7601 39144 7687 39200
rect 7743 39144 7829 39200
rect 7885 39144 7971 39200
rect 8027 39144 8113 39200
rect 8169 39144 8255 39200
rect 8311 39144 8397 39200
rect 8453 39144 8539 39200
rect 8595 39144 8681 39200
rect 8737 39144 8823 39200
rect 8879 39144 8965 39200
rect 9021 39144 9107 39200
rect 9163 39144 9249 39200
rect 9305 39144 9391 39200
rect 9447 39144 9533 39200
rect 9589 39144 9675 39200
rect 9731 39144 9817 39200
rect 9873 39144 9959 39200
rect 10015 39144 10101 39200
rect 10157 39144 10243 39200
rect 10299 39144 10385 39200
rect 10441 39144 10527 39200
rect 10583 39144 10669 39200
rect 10725 39144 10811 39200
rect 10867 39144 10953 39200
rect 11009 39144 11095 39200
rect 11151 39144 11237 39200
rect 11293 39144 11379 39200
rect 11435 39144 11521 39200
rect 11577 39144 11663 39200
rect 11719 39144 11805 39200
rect 11861 39144 11947 39200
rect 12003 39144 12089 39200
rect 12145 39144 12231 39200
rect 12287 39144 12373 39200
rect 12429 39144 12515 39200
rect 12571 39144 12657 39200
rect 12713 39144 12799 39200
rect 12855 39144 12941 39200
rect 12997 39144 13083 39200
rect 13139 39144 13225 39200
rect 13281 39144 13367 39200
rect 13423 39144 13509 39200
rect 13565 39144 13651 39200
rect 13707 39144 13793 39200
rect 13849 39144 13935 39200
rect 13991 39144 14077 39200
rect 14133 39144 14219 39200
rect 14275 39144 14361 39200
rect 14417 39144 14503 39200
rect 14559 39144 14645 39200
rect 14701 39144 14787 39200
rect 14843 39144 15000 39200
rect 0 39058 15000 39144
rect 0 39002 161 39058
rect 217 39002 303 39058
rect 359 39002 445 39058
rect 501 39002 587 39058
rect 643 39002 729 39058
rect 785 39002 871 39058
rect 927 39002 1013 39058
rect 1069 39002 1155 39058
rect 1211 39002 1297 39058
rect 1353 39002 1439 39058
rect 1495 39002 1581 39058
rect 1637 39002 1723 39058
rect 1779 39002 1865 39058
rect 1921 39002 2007 39058
rect 2063 39002 2149 39058
rect 2205 39002 2291 39058
rect 2347 39002 2433 39058
rect 2489 39002 2575 39058
rect 2631 39002 2717 39058
rect 2773 39002 2859 39058
rect 2915 39002 3001 39058
rect 3057 39002 3143 39058
rect 3199 39002 3285 39058
rect 3341 39002 3427 39058
rect 3483 39002 3569 39058
rect 3625 39002 3711 39058
rect 3767 39002 3853 39058
rect 3909 39002 3995 39058
rect 4051 39002 4137 39058
rect 4193 39002 4279 39058
rect 4335 39002 4421 39058
rect 4477 39002 4563 39058
rect 4619 39002 4705 39058
rect 4761 39002 4847 39058
rect 4903 39002 4989 39058
rect 5045 39002 5131 39058
rect 5187 39002 5273 39058
rect 5329 39002 5415 39058
rect 5471 39002 5557 39058
rect 5613 39002 5699 39058
rect 5755 39002 5841 39058
rect 5897 39002 5983 39058
rect 6039 39002 6125 39058
rect 6181 39002 6267 39058
rect 6323 39002 6409 39058
rect 6465 39002 6551 39058
rect 6607 39002 6693 39058
rect 6749 39002 6835 39058
rect 6891 39002 6977 39058
rect 7033 39002 7119 39058
rect 7175 39002 7261 39058
rect 7317 39002 7403 39058
rect 7459 39002 7545 39058
rect 7601 39002 7687 39058
rect 7743 39002 7829 39058
rect 7885 39002 7971 39058
rect 8027 39002 8113 39058
rect 8169 39002 8255 39058
rect 8311 39002 8397 39058
rect 8453 39002 8539 39058
rect 8595 39002 8681 39058
rect 8737 39002 8823 39058
rect 8879 39002 8965 39058
rect 9021 39002 9107 39058
rect 9163 39002 9249 39058
rect 9305 39002 9391 39058
rect 9447 39002 9533 39058
rect 9589 39002 9675 39058
rect 9731 39002 9817 39058
rect 9873 39002 9959 39058
rect 10015 39002 10101 39058
rect 10157 39002 10243 39058
rect 10299 39002 10385 39058
rect 10441 39002 10527 39058
rect 10583 39002 10669 39058
rect 10725 39002 10811 39058
rect 10867 39002 10953 39058
rect 11009 39002 11095 39058
rect 11151 39002 11237 39058
rect 11293 39002 11379 39058
rect 11435 39002 11521 39058
rect 11577 39002 11663 39058
rect 11719 39002 11805 39058
rect 11861 39002 11947 39058
rect 12003 39002 12089 39058
rect 12145 39002 12231 39058
rect 12287 39002 12373 39058
rect 12429 39002 12515 39058
rect 12571 39002 12657 39058
rect 12713 39002 12799 39058
rect 12855 39002 12941 39058
rect 12997 39002 13083 39058
rect 13139 39002 13225 39058
rect 13281 39002 13367 39058
rect 13423 39002 13509 39058
rect 13565 39002 13651 39058
rect 13707 39002 13793 39058
rect 13849 39002 13935 39058
rect 13991 39002 14077 39058
rect 14133 39002 14219 39058
rect 14275 39002 14361 39058
rect 14417 39002 14503 39058
rect 14559 39002 14645 39058
rect 14701 39002 14787 39058
rect 14843 39002 15000 39058
rect 0 38916 15000 39002
rect 0 38860 161 38916
rect 217 38860 303 38916
rect 359 38860 445 38916
rect 501 38860 587 38916
rect 643 38860 729 38916
rect 785 38860 871 38916
rect 927 38860 1013 38916
rect 1069 38860 1155 38916
rect 1211 38860 1297 38916
rect 1353 38860 1439 38916
rect 1495 38860 1581 38916
rect 1637 38860 1723 38916
rect 1779 38860 1865 38916
rect 1921 38860 2007 38916
rect 2063 38860 2149 38916
rect 2205 38860 2291 38916
rect 2347 38860 2433 38916
rect 2489 38860 2575 38916
rect 2631 38860 2717 38916
rect 2773 38860 2859 38916
rect 2915 38860 3001 38916
rect 3057 38860 3143 38916
rect 3199 38860 3285 38916
rect 3341 38860 3427 38916
rect 3483 38860 3569 38916
rect 3625 38860 3711 38916
rect 3767 38860 3853 38916
rect 3909 38860 3995 38916
rect 4051 38860 4137 38916
rect 4193 38860 4279 38916
rect 4335 38860 4421 38916
rect 4477 38860 4563 38916
rect 4619 38860 4705 38916
rect 4761 38860 4847 38916
rect 4903 38860 4989 38916
rect 5045 38860 5131 38916
rect 5187 38860 5273 38916
rect 5329 38860 5415 38916
rect 5471 38860 5557 38916
rect 5613 38860 5699 38916
rect 5755 38860 5841 38916
rect 5897 38860 5983 38916
rect 6039 38860 6125 38916
rect 6181 38860 6267 38916
rect 6323 38860 6409 38916
rect 6465 38860 6551 38916
rect 6607 38860 6693 38916
rect 6749 38860 6835 38916
rect 6891 38860 6977 38916
rect 7033 38860 7119 38916
rect 7175 38860 7261 38916
rect 7317 38860 7403 38916
rect 7459 38860 7545 38916
rect 7601 38860 7687 38916
rect 7743 38860 7829 38916
rect 7885 38860 7971 38916
rect 8027 38860 8113 38916
rect 8169 38860 8255 38916
rect 8311 38860 8397 38916
rect 8453 38860 8539 38916
rect 8595 38860 8681 38916
rect 8737 38860 8823 38916
rect 8879 38860 8965 38916
rect 9021 38860 9107 38916
rect 9163 38860 9249 38916
rect 9305 38860 9391 38916
rect 9447 38860 9533 38916
rect 9589 38860 9675 38916
rect 9731 38860 9817 38916
rect 9873 38860 9959 38916
rect 10015 38860 10101 38916
rect 10157 38860 10243 38916
rect 10299 38860 10385 38916
rect 10441 38860 10527 38916
rect 10583 38860 10669 38916
rect 10725 38860 10811 38916
rect 10867 38860 10953 38916
rect 11009 38860 11095 38916
rect 11151 38860 11237 38916
rect 11293 38860 11379 38916
rect 11435 38860 11521 38916
rect 11577 38860 11663 38916
rect 11719 38860 11805 38916
rect 11861 38860 11947 38916
rect 12003 38860 12089 38916
rect 12145 38860 12231 38916
rect 12287 38860 12373 38916
rect 12429 38860 12515 38916
rect 12571 38860 12657 38916
rect 12713 38860 12799 38916
rect 12855 38860 12941 38916
rect 12997 38860 13083 38916
rect 13139 38860 13225 38916
rect 13281 38860 13367 38916
rect 13423 38860 13509 38916
rect 13565 38860 13651 38916
rect 13707 38860 13793 38916
rect 13849 38860 13935 38916
rect 13991 38860 14077 38916
rect 14133 38860 14219 38916
rect 14275 38860 14361 38916
rect 14417 38860 14503 38916
rect 14559 38860 14645 38916
rect 14701 38860 14787 38916
rect 14843 38860 15000 38916
rect 0 38774 15000 38860
rect 0 38718 161 38774
rect 217 38718 303 38774
rect 359 38718 445 38774
rect 501 38718 587 38774
rect 643 38718 729 38774
rect 785 38718 871 38774
rect 927 38718 1013 38774
rect 1069 38718 1155 38774
rect 1211 38718 1297 38774
rect 1353 38718 1439 38774
rect 1495 38718 1581 38774
rect 1637 38718 1723 38774
rect 1779 38718 1865 38774
rect 1921 38718 2007 38774
rect 2063 38718 2149 38774
rect 2205 38718 2291 38774
rect 2347 38718 2433 38774
rect 2489 38718 2575 38774
rect 2631 38718 2717 38774
rect 2773 38718 2859 38774
rect 2915 38718 3001 38774
rect 3057 38718 3143 38774
rect 3199 38718 3285 38774
rect 3341 38718 3427 38774
rect 3483 38718 3569 38774
rect 3625 38718 3711 38774
rect 3767 38718 3853 38774
rect 3909 38718 3995 38774
rect 4051 38718 4137 38774
rect 4193 38718 4279 38774
rect 4335 38718 4421 38774
rect 4477 38718 4563 38774
rect 4619 38718 4705 38774
rect 4761 38718 4847 38774
rect 4903 38718 4989 38774
rect 5045 38718 5131 38774
rect 5187 38718 5273 38774
rect 5329 38718 5415 38774
rect 5471 38718 5557 38774
rect 5613 38718 5699 38774
rect 5755 38718 5841 38774
rect 5897 38718 5983 38774
rect 6039 38718 6125 38774
rect 6181 38718 6267 38774
rect 6323 38718 6409 38774
rect 6465 38718 6551 38774
rect 6607 38718 6693 38774
rect 6749 38718 6835 38774
rect 6891 38718 6977 38774
rect 7033 38718 7119 38774
rect 7175 38718 7261 38774
rect 7317 38718 7403 38774
rect 7459 38718 7545 38774
rect 7601 38718 7687 38774
rect 7743 38718 7829 38774
rect 7885 38718 7971 38774
rect 8027 38718 8113 38774
rect 8169 38718 8255 38774
rect 8311 38718 8397 38774
rect 8453 38718 8539 38774
rect 8595 38718 8681 38774
rect 8737 38718 8823 38774
rect 8879 38718 8965 38774
rect 9021 38718 9107 38774
rect 9163 38718 9249 38774
rect 9305 38718 9391 38774
rect 9447 38718 9533 38774
rect 9589 38718 9675 38774
rect 9731 38718 9817 38774
rect 9873 38718 9959 38774
rect 10015 38718 10101 38774
rect 10157 38718 10243 38774
rect 10299 38718 10385 38774
rect 10441 38718 10527 38774
rect 10583 38718 10669 38774
rect 10725 38718 10811 38774
rect 10867 38718 10953 38774
rect 11009 38718 11095 38774
rect 11151 38718 11237 38774
rect 11293 38718 11379 38774
rect 11435 38718 11521 38774
rect 11577 38718 11663 38774
rect 11719 38718 11805 38774
rect 11861 38718 11947 38774
rect 12003 38718 12089 38774
rect 12145 38718 12231 38774
rect 12287 38718 12373 38774
rect 12429 38718 12515 38774
rect 12571 38718 12657 38774
rect 12713 38718 12799 38774
rect 12855 38718 12941 38774
rect 12997 38718 13083 38774
rect 13139 38718 13225 38774
rect 13281 38718 13367 38774
rect 13423 38718 13509 38774
rect 13565 38718 13651 38774
rect 13707 38718 13793 38774
rect 13849 38718 13935 38774
rect 13991 38718 14077 38774
rect 14133 38718 14219 38774
rect 14275 38718 14361 38774
rect 14417 38718 14503 38774
rect 14559 38718 14645 38774
rect 14701 38718 14787 38774
rect 14843 38718 15000 38774
rect 0 38632 15000 38718
rect 0 38576 161 38632
rect 217 38576 303 38632
rect 359 38576 445 38632
rect 501 38576 587 38632
rect 643 38576 729 38632
rect 785 38576 871 38632
rect 927 38576 1013 38632
rect 1069 38576 1155 38632
rect 1211 38576 1297 38632
rect 1353 38576 1439 38632
rect 1495 38576 1581 38632
rect 1637 38576 1723 38632
rect 1779 38576 1865 38632
rect 1921 38576 2007 38632
rect 2063 38576 2149 38632
rect 2205 38576 2291 38632
rect 2347 38576 2433 38632
rect 2489 38576 2575 38632
rect 2631 38576 2717 38632
rect 2773 38576 2859 38632
rect 2915 38576 3001 38632
rect 3057 38576 3143 38632
rect 3199 38576 3285 38632
rect 3341 38576 3427 38632
rect 3483 38576 3569 38632
rect 3625 38576 3711 38632
rect 3767 38576 3853 38632
rect 3909 38576 3995 38632
rect 4051 38576 4137 38632
rect 4193 38576 4279 38632
rect 4335 38576 4421 38632
rect 4477 38576 4563 38632
rect 4619 38576 4705 38632
rect 4761 38576 4847 38632
rect 4903 38576 4989 38632
rect 5045 38576 5131 38632
rect 5187 38576 5273 38632
rect 5329 38576 5415 38632
rect 5471 38576 5557 38632
rect 5613 38576 5699 38632
rect 5755 38576 5841 38632
rect 5897 38576 5983 38632
rect 6039 38576 6125 38632
rect 6181 38576 6267 38632
rect 6323 38576 6409 38632
rect 6465 38576 6551 38632
rect 6607 38576 6693 38632
rect 6749 38576 6835 38632
rect 6891 38576 6977 38632
rect 7033 38576 7119 38632
rect 7175 38576 7261 38632
rect 7317 38576 7403 38632
rect 7459 38576 7545 38632
rect 7601 38576 7687 38632
rect 7743 38576 7829 38632
rect 7885 38576 7971 38632
rect 8027 38576 8113 38632
rect 8169 38576 8255 38632
rect 8311 38576 8397 38632
rect 8453 38576 8539 38632
rect 8595 38576 8681 38632
rect 8737 38576 8823 38632
rect 8879 38576 8965 38632
rect 9021 38576 9107 38632
rect 9163 38576 9249 38632
rect 9305 38576 9391 38632
rect 9447 38576 9533 38632
rect 9589 38576 9675 38632
rect 9731 38576 9817 38632
rect 9873 38576 9959 38632
rect 10015 38576 10101 38632
rect 10157 38576 10243 38632
rect 10299 38576 10385 38632
rect 10441 38576 10527 38632
rect 10583 38576 10669 38632
rect 10725 38576 10811 38632
rect 10867 38576 10953 38632
rect 11009 38576 11095 38632
rect 11151 38576 11237 38632
rect 11293 38576 11379 38632
rect 11435 38576 11521 38632
rect 11577 38576 11663 38632
rect 11719 38576 11805 38632
rect 11861 38576 11947 38632
rect 12003 38576 12089 38632
rect 12145 38576 12231 38632
rect 12287 38576 12373 38632
rect 12429 38576 12515 38632
rect 12571 38576 12657 38632
rect 12713 38576 12799 38632
rect 12855 38576 12941 38632
rect 12997 38576 13083 38632
rect 13139 38576 13225 38632
rect 13281 38576 13367 38632
rect 13423 38576 13509 38632
rect 13565 38576 13651 38632
rect 13707 38576 13793 38632
rect 13849 38576 13935 38632
rect 13991 38576 14077 38632
rect 14133 38576 14219 38632
rect 14275 38576 14361 38632
rect 14417 38576 14503 38632
rect 14559 38576 14645 38632
rect 14701 38576 14787 38632
rect 14843 38576 15000 38632
rect 0 38490 15000 38576
rect 0 38434 161 38490
rect 217 38434 303 38490
rect 359 38434 445 38490
rect 501 38434 587 38490
rect 643 38434 729 38490
rect 785 38434 871 38490
rect 927 38434 1013 38490
rect 1069 38434 1155 38490
rect 1211 38434 1297 38490
rect 1353 38434 1439 38490
rect 1495 38434 1581 38490
rect 1637 38434 1723 38490
rect 1779 38434 1865 38490
rect 1921 38434 2007 38490
rect 2063 38434 2149 38490
rect 2205 38434 2291 38490
rect 2347 38434 2433 38490
rect 2489 38434 2575 38490
rect 2631 38434 2717 38490
rect 2773 38434 2859 38490
rect 2915 38434 3001 38490
rect 3057 38434 3143 38490
rect 3199 38434 3285 38490
rect 3341 38434 3427 38490
rect 3483 38434 3569 38490
rect 3625 38434 3711 38490
rect 3767 38434 3853 38490
rect 3909 38434 3995 38490
rect 4051 38434 4137 38490
rect 4193 38434 4279 38490
rect 4335 38434 4421 38490
rect 4477 38434 4563 38490
rect 4619 38434 4705 38490
rect 4761 38434 4847 38490
rect 4903 38434 4989 38490
rect 5045 38434 5131 38490
rect 5187 38434 5273 38490
rect 5329 38434 5415 38490
rect 5471 38434 5557 38490
rect 5613 38434 5699 38490
rect 5755 38434 5841 38490
rect 5897 38434 5983 38490
rect 6039 38434 6125 38490
rect 6181 38434 6267 38490
rect 6323 38434 6409 38490
rect 6465 38434 6551 38490
rect 6607 38434 6693 38490
rect 6749 38434 6835 38490
rect 6891 38434 6977 38490
rect 7033 38434 7119 38490
rect 7175 38434 7261 38490
rect 7317 38434 7403 38490
rect 7459 38434 7545 38490
rect 7601 38434 7687 38490
rect 7743 38434 7829 38490
rect 7885 38434 7971 38490
rect 8027 38434 8113 38490
rect 8169 38434 8255 38490
rect 8311 38434 8397 38490
rect 8453 38434 8539 38490
rect 8595 38434 8681 38490
rect 8737 38434 8823 38490
rect 8879 38434 8965 38490
rect 9021 38434 9107 38490
rect 9163 38434 9249 38490
rect 9305 38434 9391 38490
rect 9447 38434 9533 38490
rect 9589 38434 9675 38490
rect 9731 38434 9817 38490
rect 9873 38434 9959 38490
rect 10015 38434 10101 38490
rect 10157 38434 10243 38490
rect 10299 38434 10385 38490
rect 10441 38434 10527 38490
rect 10583 38434 10669 38490
rect 10725 38434 10811 38490
rect 10867 38434 10953 38490
rect 11009 38434 11095 38490
rect 11151 38434 11237 38490
rect 11293 38434 11379 38490
rect 11435 38434 11521 38490
rect 11577 38434 11663 38490
rect 11719 38434 11805 38490
rect 11861 38434 11947 38490
rect 12003 38434 12089 38490
rect 12145 38434 12231 38490
rect 12287 38434 12373 38490
rect 12429 38434 12515 38490
rect 12571 38434 12657 38490
rect 12713 38434 12799 38490
rect 12855 38434 12941 38490
rect 12997 38434 13083 38490
rect 13139 38434 13225 38490
rect 13281 38434 13367 38490
rect 13423 38434 13509 38490
rect 13565 38434 13651 38490
rect 13707 38434 13793 38490
rect 13849 38434 13935 38490
rect 13991 38434 14077 38490
rect 14133 38434 14219 38490
rect 14275 38434 14361 38490
rect 14417 38434 14503 38490
rect 14559 38434 14645 38490
rect 14701 38434 14787 38490
rect 14843 38434 15000 38490
rect 0 38348 15000 38434
rect 0 38292 161 38348
rect 217 38292 303 38348
rect 359 38292 445 38348
rect 501 38292 587 38348
rect 643 38292 729 38348
rect 785 38292 871 38348
rect 927 38292 1013 38348
rect 1069 38292 1155 38348
rect 1211 38292 1297 38348
rect 1353 38292 1439 38348
rect 1495 38292 1581 38348
rect 1637 38292 1723 38348
rect 1779 38292 1865 38348
rect 1921 38292 2007 38348
rect 2063 38292 2149 38348
rect 2205 38292 2291 38348
rect 2347 38292 2433 38348
rect 2489 38292 2575 38348
rect 2631 38292 2717 38348
rect 2773 38292 2859 38348
rect 2915 38292 3001 38348
rect 3057 38292 3143 38348
rect 3199 38292 3285 38348
rect 3341 38292 3427 38348
rect 3483 38292 3569 38348
rect 3625 38292 3711 38348
rect 3767 38292 3853 38348
rect 3909 38292 3995 38348
rect 4051 38292 4137 38348
rect 4193 38292 4279 38348
rect 4335 38292 4421 38348
rect 4477 38292 4563 38348
rect 4619 38292 4705 38348
rect 4761 38292 4847 38348
rect 4903 38292 4989 38348
rect 5045 38292 5131 38348
rect 5187 38292 5273 38348
rect 5329 38292 5415 38348
rect 5471 38292 5557 38348
rect 5613 38292 5699 38348
rect 5755 38292 5841 38348
rect 5897 38292 5983 38348
rect 6039 38292 6125 38348
rect 6181 38292 6267 38348
rect 6323 38292 6409 38348
rect 6465 38292 6551 38348
rect 6607 38292 6693 38348
rect 6749 38292 6835 38348
rect 6891 38292 6977 38348
rect 7033 38292 7119 38348
rect 7175 38292 7261 38348
rect 7317 38292 7403 38348
rect 7459 38292 7545 38348
rect 7601 38292 7687 38348
rect 7743 38292 7829 38348
rect 7885 38292 7971 38348
rect 8027 38292 8113 38348
rect 8169 38292 8255 38348
rect 8311 38292 8397 38348
rect 8453 38292 8539 38348
rect 8595 38292 8681 38348
rect 8737 38292 8823 38348
rect 8879 38292 8965 38348
rect 9021 38292 9107 38348
rect 9163 38292 9249 38348
rect 9305 38292 9391 38348
rect 9447 38292 9533 38348
rect 9589 38292 9675 38348
rect 9731 38292 9817 38348
rect 9873 38292 9959 38348
rect 10015 38292 10101 38348
rect 10157 38292 10243 38348
rect 10299 38292 10385 38348
rect 10441 38292 10527 38348
rect 10583 38292 10669 38348
rect 10725 38292 10811 38348
rect 10867 38292 10953 38348
rect 11009 38292 11095 38348
rect 11151 38292 11237 38348
rect 11293 38292 11379 38348
rect 11435 38292 11521 38348
rect 11577 38292 11663 38348
rect 11719 38292 11805 38348
rect 11861 38292 11947 38348
rect 12003 38292 12089 38348
rect 12145 38292 12231 38348
rect 12287 38292 12373 38348
rect 12429 38292 12515 38348
rect 12571 38292 12657 38348
rect 12713 38292 12799 38348
rect 12855 38292 12941 38348
rect 12997 38292 13083 38348
rect 13139 38292 13225 38348
rect 13281 38292 13367 38348
rect 13423 38292 13509 38348
rect 13565 38292 13651 38348
rect 13707 38292 13793 38348
rect 13849 38292 13935 38348
rect 13991 38292 14077 38348
rect 14133 38292 14219 38348
rect 14275 38292 14361 38348
rect 14417 38292 14503 38348
rect 14559 38292 14645 38348
rect 14701 38292 14787 38348
rect 14843 38292 15000 38348
rect 0 38206 15000 38292
rect 0 38150 161 38206
rect 217 38150 303 38206
rect 359 38150 445 38206
rect 501 38150 587 38206
rect 643 38150 729 38206
rect 785 38150 871 38206
rect 927 38150 1013 38206
rect 1069 38150 1155 38206
rect 1211 38150 1297 38206
rect 1353 38150 1439 38206
rect 1495 38150 1581 38206
rect 1637 38150 1723 38206
rect 1779 38150 1865 38206
rect 1921 38150 2007 38206
rect 2063 38150 2149 38206
rect 2205 38150 2291 38206
rect 2347 38150 2433 38206
rect 2489 38150 2575 38206
rect 2631 38150 2717 38206
rect 2773 38150 2859 38206
rect 2915 38150 3001 38206
rect 3057 38150 3143 38206
rect 3199 38150 3285 38206
rect 3341 38150 3427 38206
rect 3483 38150 3569 38206
rect 3625 38150 3711 38206
rect 3767 38150 3853 38206
rect 3909 38150 3995 38206
rect 4051 38150 4137 38206
rect 4193 38150 4279 38206
rect 4335 38150 4421 38206
rect 4477 38150 4563 38206
rect 4619 38150 4705 38206
rect 4761 38150 4847 38206
rect 4903 38150 4989 38206
rect 5045 38150 5131 38206
rect 5187 38150 5273 38206
rect 5329 38150 5415 38206
rect 5471 38150 5557 38206
rect 5613 38150 5699 38206
rect 5755 38150 5841 38206
rect 5897 38150 5983 38206
rect 6039 38150 6125 38206
rect 6181 38150 6267 38206
rect 6323 38150 6409 38206
rect 6465 38150 6551 38206
rect 6607 38150 6693 38206
rect 6749 38150 6835 38206
rect 6891 38150 6977 38206
rect 7033 38150 7119 38206
rect 7175 38150 7261 38206
rect 7317 38150 7403 38206
rect 7459 38150 7545 38206
rect 7601 38150 7687 38206
rect 7743 38150 7829 38206
rect 7885 38150 7971 38206
rect 8027 38150 8113 38206
rect 8169 38150 8255 38206
rect 8311 38150 8397 38206
rect 8453 38150 8539 38206
rect 8595 38150 8681 38206
rect 8737 38150 8823 38206
rect 8879 38150 8965 38206
rect 9021 38150 9107 38206
rect 9163 38150 9249 38206
rect 9305 38150 9391 38206
rect 9447 38150 9533 38206
rect 9589 38150 9675 38206
rect 9731 38150 9817 38206
rect 9873 38150 9959 38206
rect 10015 38150 10101 38206
rect 10157 38150 10243 38206
rect 10299 38150 10385 38206
rect 10441 38150 10527 38206
rect 10583 38150 10669 38206
rect 10725 38150 10811 38206
rect 10867 38150 10953 38206
rect 11009 38150 11095 38206
rect 11151 38150 11237 38206
rect 11293 38150 11379 38206
rect 11435 38150 11521 38206
rect 11577 38150 11663 38206
rect 11719 38150 11805 38206
rect 11861 38150 11947 38206
rect 12003 38150 12089 38206
rect 12145 38150 12231 38206
rect 12287 38150 12373 38206
rect 12429 38150 12515 38206
rect 12571 38150 12657 38206
rect 12713 38150 12799 38206
rect 12855 38150 12941 38206
rect 12997 38150 13083 38206
rect 13139 38150 13225 38206
rect 13281 38150 13367 38206
rect 13423 38150 13509 38206
rect 13565 38150 13651 38206
rect 13707 38150 13793 38206
rect 13849 38150 13935 38206
rect 13991 38150 14077 38206
rect 14133 38150 14219 38206
rect 14275 38150 14361 38206
rect 14417 38150 14503 38206
rect 14559 38150 14645 38206
rect 14701 38150 14787 38206
rect 14843 38150 15000 38206
rect 0 38064 15000 38150
rect 0 38008 161 38064
rect 217 38008 303 38064
rect 359 38008 445 38064
rect 501 38008 587 38064
rect 643 38008 729 38064
rect 785 38008 871 38064
rect 927 38008 1013 38064
rect 1069 38008 1155 38064
rect 1211 38008 1297 38064
rect 1353 38008 1439 38064
rect 1495 38008 1581 38064
rect 1637 38008 1723 38064
rect 1779 38008 1865 38064
rect 1921 38008 2007 38064
rect 2063 38008 2149 38064
rect 2205 38008 2291 38064
rect 2347 38008 2433 38064
rect 2489 38008 2575 38064
rect 2631 38008 2717 38064
rect 2773 38008 2859 38064
rect 2915 38008 3001 38064
rect 3057 38008 3143 38064
rect 3199 38008 3285 38064
rect 3341 38008 3427 38064
rect 3483 38008 3569 38064
rect 3625 38008 3711 38064
rect 3767 38008 3853 38064
rect 3909 38008 3995 38064
rect 4051 38008 4137 38064
rect 4193 38008 4279 38064
rect 4335 38008 4421 38064
rect 4477 38008 4563 38064
rect 4619 38008 4705 38064
rect 4761 38008 4847 38064
rect 4903 38008 4989 38064
rect 5045 38008 5131 38064
rect 5187 38008 5273 38064
rect 5329 38008 5415 38064
rect 5471 38008 5557 38064
rect 5613 38008 5699 38064
rect 5755 38008 5841 38064
rect 5897 38008 5983 38064
rect 6039 38008 6125 38064
rect 6181 38008 6267 38064
rect 6323 38008 6409 38064
rect 6465 38008 6551 38064
rect 6607 38008 6693 38064
rect 6749 38008 6835 38064
rect 6891 38008 6977 38064
rect 7033 38008 7119 38064
rect 7175 38008 7261 38064
rect 7317 38008 7403 38064
rect 7459 38008 7545 38064
rect 7601 38008 7687 38064
rect 7743 38008 7829 38064
rect 7885 38008 7971 38064
rect 8027 38008 8113 38064
rect 8169 38008 8255 38064
rect 8311 38008 8397 38064
rect 8453 38008 8539 38064
rect 8595 38008 8681 38064
rect 8737 38008 8823 38064
rect 8879 38008 8965 38064
rect 9021 38008 9107 38064
rect 9163 38008 9249 38064
rect 9305 38008 9391 38064
rect 9447 38008 9533 38064
rect 9589 38008 9675 38064
rect 9731 38008 9817 38064
rect 9873 38008 9959 38064
rect 10015 38008 10101 38064
rect 10157 38008 10243 38064
rect 10299 38008 10385 38064
rect 10441 38008 10527 38064
rect 10583 38008 10669 38064
rect 10725 38008 10811 38064
rect 10867 38008 10953 38064
rect 11009 38008 11095 38064
rect 11151 38008 11237 38064
rect 11293 38008 11379 38064
rect 11435 38008 11521 38064
rect 11577 38008 11663 38064
rect 11719 38008 11805 38064
rect 11861 38008 11947 38064
rect 12003 38008 12089 38064
rect 12145 38008 12231 38064
rect 12287 38008 12373 38064
rect 12429 38008 12515 38064
rect 12571 38008 12657 38064
rect 12713 38008 12799 38064
rect 12855 38008 12941 38064
rect 12997 38008 13083 38064
rect 13139 38008 13225 38064
rect 13281 38008 13367 38064
rect 13423 38008 13509 38064
rect 13565 38008 13651 38064
rect 13707 38008 13793 38064
rect 13849 38008 13935 38064
rect 13991 38008 14077 38064
rect 14133 38008 14219 38064
rect 14275 38008 14361 38064
rect 14417 38008 14503 38064
rect 14559 38008 14645 38064
rect 14701 38008 14787 38064
rect 14843 38008 15000 38064
rect 0 37922 15000 38008
rect 0 37866 161 37922
rect 217 37866 303 37922
rect 359 37866 445 37922
rect 501 37866 587 37922
rect 643 37866 729 37922
rect 785 37866 871 37922
rect 927 37866 1013 37922
rect 1069 37866 1155 37922
rect 1211 37866 1297 37922
rect 1353 37866 1439 37922
rect 1495 37866 1581 37922
rect 1637 37866 1723 37922
rect 1779 37866 1865 37922
rect 1921 37866 2007 37922
rect 2063 37866 2149 37922
rect 2205 37866 2291 37922
rect 2347 37866 2433 37922
rect 2489 37866 2575 37922
rect 2631 37866 2717 37922
rect 2773 37866 2859 37922
rect 2915 37866 3001 37922
rect 3057 37866 3143 37922
rect 3199 37866 3285 37922
rect 3341 37866 3427 37922
rect 3483 37866 3569 37922
rect 3625 37866 3711 37922
rect 3767 37866 3853 37922
rect 3909 37866 3995 37922
rect 4051 37866 4137 37922
rect 4193 37866 4279 37922
rect 4335 37866 4421 37922
rect 4477 37866 4563 37922
rect 4619 37866 4705 37922
rect 4761 37866 4847 37922
rect 4903 37866 4989 37922
rect 5045 37866 5131 37922
rect 5187 37866 5273 37922
rect 5329 37866 5415 37922
rect 5471 37866 5557 37922
rect 5613 37866 5699 37922
rect 5755 37866 5841 37922
rect 5897 37866 5983 37922
rect 6039 37866 6125 37922
rect 6181 37866 6267 37922
rect 6323 37866 6409 37922
rect 6465 37866 6551 37922
rect 6607 37866 6693 37922
rect 6749 37866 6835 37922
rect 6891 37866 6977 37922
rect 7033 37866 7119 37922
rect 7175 37866 7261 37922
rect 7317 37866 7403 37922
rect 7459 37866 7545 37922
rect 7601 37866 7687 37922
rect 7743 37866 7829 37922
rect 7885 37866 7971 37922
rect 8027 37866 8113 37922
rect 8169 37866 8255 37922
rect 8311 37866 8397 37922
rect 8453 37866 8539 37922
rect 8595 37866 8681 37922
rect 8737 37866 8823 37922
rect 8879 37866 8965 37922
rect 9021 37866 9107 37922
rect 9163 37866 9249 37922
rect 9305 37866 9391 37922
rect 9447 37866 9533 37922
rect 9589 37866 9675 37922
rect 9731 37866 9817 37922
rect 9873 37866 9959 37922
rect 10015 37866 10101 37922
rect 10157 37866 10243 37922
rect 10299 37866 10385 37922
rect 10441 37866 10527 37922
rect 10583 37866 10669 37922
rect 10725 37866 10811 37922
rect 10867 37866 10953 37922
rect 11009 37866 11095 37922
rect 11151 37866 11237 37922
rect 11293 37866 11379 37922
rect 11435 37866 11521 37922
rect 11577 37866 11663 37922
rect 11719 37866 11805 37922
rect 11861 37866 11947 37922
rect 12003 37866 12089 37922
rect 12145 37866 12231 37922
rect 12287 37866 12373 37922
rect 12429 37866 12515 37922
rect 12571 37866 12657 37922
rect 12713 37866 12799 37922
rect 12855 37866 12941 37922
rect 12997 37866 13083 37922
rect 13139 37866 13225 37922
rect 13281 37866 13367 37922
rect 13423 37866 13509 37922
rect 13565 37866 13651 37922
rect 13707 37866 13793 37922
rect 13849 37866 13935 37922
rect 13991 37866 14077 37922
rect 14133 37866 14219 37922
rect 14275 37866 14361 37922
rect 14417 37866 14503 37922
rect 14559 37866 14645 37922
rect 14701 37866 14787 37922
rect 14843 37866 15000 37922
rect 0 37780 15000 37866
rect 0 37724 161 37780
rect 217 37724 303 37780
rect 359 37724 445 37780
rect 501 37724 587 37780
rect 643 37724 729 37780
rect 785 37724 871 37780
rect 927 37724 1013 37780
rect 1069 37724 1155 37780
rect 1211 37724 1297 37780
rect 1353 37724 1439 37780
rect 1495 37724 1581 37780
rect 1637 37724 1723 37780
rect 1779 37724 1865 37780
rect 1921 37724 2007 37780
rect 2063 37724 2149 37780
rect 2205 37724 2291 37780
rect 2347 37724 2433 37780
rect 2489 37724 2575 37780
rect 2631 37724 2717 37780
rect 2773 37724 2859 37780
rect 2915 37724 3001 37780
rect 3057 37724 3143 37780
rect 3199 37724 3285 37780
rect 3341 37724 3427 37780
rect 3483 37724 3569 37780
rect 3625 37724 3711 37780
rect 3767 37724 3853 37780
rect 3909 37724 3995 37780
rect 4051 37724 4137 37780
rect 4193 37724 4279 37780
rect 4335 37724 4421 37780
rect 4477 37724 4563 37780
rect 4619 37724 4705 37780
rect 4761 37724 4847 37780
rect 4903 37724 4989 37780
rect 5045 37724 5131 37780
rect 5187 37724 5273 37780
rect 5329 37724 5415 37780
rect 5471 37724 5557 37780
rect 5613 37724 5699 37780
rect 5755 37724 5841 37780
rect 5897 37724 5983 37780
rect 6039 37724 6125 37780
rect 6181 37724 6267 37780
rect 6323 37724 6409 37780
rect 6465 37724 6551 37780
rect 6607 37724 6693 37780
rect 6749 37724 6835 37780
rect 6891 37724 6977 37780
rect 7033 37724 7119 37780
rect 7175 37724 7261 37780
rect 7317 37724 7403 37780
rect 7459 37724 7545 37780
rect 7601 37724 7687 37780
rect 7743 37724 7829 37780
rect 7885 37724 7971 37780
rect 8027 37724 8113 37780
rect 8169 37724 8255 37780
rect 8311 37724 8397 37780
rect 8453 37724 8539 37780
rect 8595 37724 8681 37780
rect 8737 37724 8823 37780
rect 8879 37724 8965 37780
rect 9021 37724 9107 37780
rect 9163 37724 9249 37780
rect 9305 37724 9391 37780
rect 9447 37724 9533 37780
rect 9589 37724 9675 37780
rect 9731 37724 9817 37780
rect 9873 37724 9959 37780
rect 10015 37724 10101 37780
rect 10157 37724 10243 37780
rect 10299 37724 10385 37780
rect 10441 37724 10527 37780
rect 10583 37724 10669 37780
rect 10725 37724 10811 37780
rect 10867 37724 10953 37780
rect 11009 37724 11095 37780
rect 11151 37724 11237 37780
rect 11293 37724 11379 37780
rect 11435 37724 11521 37780
rect 11577 37724 11663 37780
rect 11719 37724 11805 37780
rect 11861 37724 11947 37780
rect 12003 37724 12089 37780
rect 12145 37724 12231 37780
rect 12287 37724 12373 37780
rect 12429 37724 12515 37780
rect 12571 37724 12657 37780
rect 12713 37724 12799 37780
rect 12855 37724 12941 37780
rect 12997 37724 13083 37780
rect 13139 37724 13225 37780
rect 13281 37724 13367 37780
rect 13423 37724 13509 37780
rect 13565 37724 13651 37780
rect 13707 37724 13793 37780
rect 13849 37724 13935 37780
rect 13991 37724 14077 37780
rect 14133 37724 14219 37780
rect 14275 37724 14361 37780
rect 14417 37724 14503 37780
rect 14559 37724 14645 37780
rect 14701 37724 14787 37780
rect 14843 37724 15000 37780
rect 0 37638 15000 37724
rect 0 37582 161 37638
rect 217 37582 303 37638
rect 359 37582 445 37638
rect 501 37582 587 37638
rect 643 37582 729 37638
rect 785 37582 871 37638
rect 927 37582 1013 37638
rect 1069 37582 1155 37638
rect 1211 37582 1297 37638
rect 1353 37582 1439 37638
rect 1495 37582 1581 37638
rect 1637 37582 1723 37638
rect 1779 37582 1865 37638
rect 1921 37582 2007 37638
rect 2063 37582 2149 37638
rect 2205 37582 2291 37638
rect 2347 37582 2433 37638
rect 2489 37582 2575 37638
rect 2631 37582 2717 37638
rect 2773 37582 2859 37638
rect 2915 37582 3001 37638
rect 3057 37582 3143 37638
rect 3199 37582 3285 37638
rect 3341 37582 3427 37638
rect 3483 37582 3569 37638
rect 3625 37582 3711 37638
rect 3767 37582 3853 37638
rect 3909 37582 3995 37638
rect 4051 37582 4137 37638
rect 4193 37582 4279 37638
rect 4335 37582 4421 37638
rect 4477 37582 4563 37638
rect 4619 37582 4705 37638
rect 4761 37582 4847 37638
rect 4903 37582 4989 37638
rect 5045 37582 5131 37638
rect 5187 37582 5273 37638
rect 5329 37582 5415 37638
rect 5471 37582 5557 37638
rect 5613 37582 5699 37638
rect 5755 37582 5841 37638
rect 5897 37582 5983 37638
rect 6039 37582 6125 37638
rect 6181 37582 6267 37638
rect 6323 37582 6409 37638
rect 6465 37582 6551 37638
rect 6607 37582 6693 37638
rect 6749 37582 6835 37638
rect 6891 37582 6977 37638
rect 7033 37582 7119 37638
rect 7175 37582 7261 37638
rect 7317 37582 7403 37638
rect 7459 37582 7545 37638
rect 7601 37582 7687 37638
rect 7743 37582 7829 37638
rect 7885 37582 7971 37638
rect 8027 37582 8113 37638
rect 8169 37582 8255 37638
rect 8311 37582 8397 37638
rect 8453 37582 8539 37638
rect 8595 37582 8681 37638
rect 8737 37582 8823 37638
rect 8879 37582 8965 37638
rect 9021 37582 9107 37638
rect 9163 37582 9249 37638
rect 9305 37582 9391 37638
rect 9447 37582 9533 37638
rect 9589 37582 9675 37638
rect 9731 37582 9817 37638
rect 9873 37582 9959 37638
rect 10015 37582 10101 37638
rect 10157 37582 10243 37638
rect 10299 37582 10385 37638
rect 10441 37582 10527 37638
rect 10583 37582 10669 37638
rect 10725 37582 10811 37638
rect 10867 37582 10953 37638
rect 11009 37582 11095 37638
rect 11151 37582 11237 37638
rect 11293 37582 11379 37638
rect 11435 37582 11521 37638
rect 11577 37582 11663 37638
rect 11719 37582 11805 37638
rect 11861 37582 11947 37638
rect 12003 37582 12089 37638
rect 12145 37582 12231 37638
rect 12287 37582 12373 37638
rect 12429 37582 12515 37638
rect 12571 37582 12657 37638
rect 12713 37582 12799 37638
rect 12855 37582 12941 37638
rect 12997 37582 13083 37638
rect 13139 37582 13225 37638
rect 13281 37582 13367 37638
rect 13423 37582 13509 37638
rect 13565 37582 13651 37638
rect 13707 37582 13793 37638
rect 13849 37582 13935 37638
rect 13991 37582 14077 37638
rect 14133 37582 14219 37638
rect 14275 37582 14361 37638
rect 14417 37582 14503 37638
rect 14559 37582 14645 37638
rect 14701 37582 14787 37638
rect 14843 37582 15000 37638
rect 0 37496 15000 37582
rect 0 37440 161 37496
rect 217 37440 303 37496
rect 359 37440 445 37496
rect 501 37440 587 37496
rect 643 37440 729 37496
rect 785 37440 871 37496
rect 927 37440 1013 37496
rect 1069 37440 1155 37496
rect 1211 37440 1297 37496
rect 1353 37440 1439 37496
rect 1495 37440 1581 37496
rect 1637 37440 1723 37496
rect 1779 37440 1865 37496
rect 1921 37440 2007 37496
rect 2063 37440 2149 37496
rect 2205 37440 2291 37496
rect 2347 37440 2433 37496
rect 2489 37440 2575 37496
rect 2631 37440 2717 37496
rect 2773 37440 2859 37496
rect 2915 37440 3001 37496
rect 3057 37440 3143 37496
rect 3199 37440 3285 37496
rect 3341 37440 3427 37496
rect 3483 37440 3569 37496
rect 3625 37440 3711 37496
rect 3767 37440 3853 37496
rect 3909 37440 3995 37496
rect 4051 37440 4137 37496
rect 4193 37440 4279 37496
rect 4335 37440 4421 37496
rect 4477 37440 4563 37496
rect 4619 37440 4705 37496
rect 4761 37440 4847 37496
rect 4903 37440 4989 37496
rect 5045 37440 5131 37496
rect 5187 37440 5273 37496
rect 5329 37440 5415 37496
rect 5471 37440 5557 37496
rect 5613 37440 5699 37496
rect 5755 37440 5841 37496
rect 5897 37440 5983 37496
rect 6039 37440 6125 37496
rect 6181 37440 6267 37496
rect 6323 37440 6409 37496
rect 6465 37440 6551 37496
rect 6607 37440 6693 37496
rect 6749 37440 6835 37496
rect 6891 37440 6977 37496
rect 7033 37440 7119 37496
rect 7175 37440 7261 37496
rect 7317 37440 7403 37496
rect 7459 37440 7545 37496
rect 7601 37440 7687 37496
rect 7743 37440 7829 37496
rect 7885 37440 7971 37496
rect 8027 37440 8113 37496
rect 8169 37440 8255 37496
rect 8311 37440 8397 37496
rect 8453 37440 8539 37496
rect 8595 37440 8681 37496
rect 8737 37440 8823 37496
rect 8879 37440 8965 37496
rect 9021 37440 9107 37496
rect 9163 37440 9249 37496
rect 9305 37440 9391 37496
rect 9447 37440 9533 37496
rect 9589 37440 9675 37496
rect 9731 37440 9817 37496
rect 9873 37440 9959 37496
rect 10015 37440 10101 37496
rect 10157 37440 10243 37496
rect 10299 37440 10385 37496
rect 10441 37440 10527 37496
rect 10583 37440 10669 37496
rect 10725 37440 10811 37496
rect 10867 37440 10953 37496
rect 11009 37440 11095 37496
rect 11151 37440 11237 37496
rect 11293 37440 11379 37496
rect 11435 37440 11521 37496
rect 11577 37440 11663 37496
rect 11719 37440 11805 37496
rect 11861 37440 11947 37496
rect 12003 37440 12089 37496
rect 12145 37440 12231 37496
rect 12287 37440 12373 37496
rect 12429 37440 12515 37496
rect 12571 37440 12657 37496
rect 12713 37440 12799 37496
rect 12855 37440 12941 37496
rect 12997 37440 13083 37496
rect 13139 37440 13225 37496
rect 13281 37440 13367 37496
rect 13423 37440 13509 37496
rect 13565 37440 13651 37496
rect 13707 37440 13793 37496
rect 13849 37440 13935 37496
rect 13991 37440 14077 37496
rect 14133 37440 14219 37496
rect 14275 37440 14361 37496
rect 14417 37440 14503 37496
rect 14559 37440 14645 37496
rect 14701 37440 14787 37496
rect 14843 37440 15000 37496
rect 0 37354 15000 37440
rect 0 37298 161 37354
rect 217 37298 303 37354
rect 359 37298 445 37354
rect 501 37298 587 37354
rect 643 37298 729 37354
rect 785 37298 871 37354
rect 927 37298 1013 37354
rect 1069 37298 1155 37354
rect 1211 37298 1297 37354
rect 1353 37298 1439 37354
rect 1495 37298 1581 37354
rect 1637 37298 1723 37354
rect 1779 37298 1865 37354
rect 1921 37298 2007 37354
rect 2063 37298 2149 37354
rect 2205 37298 2291 37354
rect 2347 37298 2433 37354
rect 2489 37298 2575 37354
rect 2631 37298 2717 37354
rect 2773 37298 2859 37354
rect 2915 37298 3001 37354
rect 3057 37298 3143 37354
rect 3199 37298 3285 37354
rect 3341 37298 3427 37354
rect 3483 37298 3569 37354
rect 3625 37298 3711 37354
rect 3767 37298 3853 37354
rect 3909 37298 3995 37354
rect 4051 37298 4137 37354
rect 4193 37298 4279 37354
rect 4335 37298 4421 37354
rect 4477 37298 4563 37354
rect 4619 37298 4705 37354
rect 4761 37298 4847 37354
rect 4903 37298 4989 37354
rect 5045 37298 5131 37354
rect 5187 37298 5273 37354
rect 5329 37298 5415 37354
rect 5471 37298 5557 37354
rect 5613 37298 5699 37354
rect 5755 37298 5841 37354
rect 5897 37298 5983 37354
rect 6039 37298 6125 37354
rect 6181 37298 6267 37354
rect 6323 37298 6409 37354
rect 6465 37298 6551 37354
rect 6607 37298 6693 37354
rect 6749 37298 6835 37354
rect 6891 37298 6977 37354
rect 7033 37298 7119 37354
rect 7175 37298 7261 37354
rect 7317 37298 7403 37354
rect 7459 37298 7545 37354
rect 7601 37298 7687 37354
rect 7743 37298 7829 37354
rect 7885 37298 7971 37354
rect 8027 37298 8113 37354
rect 8169 37298 8255 37354
rect 8311 37298 8397 37354
rect 8453 37298 8539 37354
rect 8595 37298 8681 37354
rect 8737 37298 8823 37354
rect 8879 37298 8965 37354
rect 9021 37298 9107 37354
rect 9163 37298 9249 37354
rect 9305 37298 9391 37354
rect 9447 37298 9533 37354
rect 9589 37298 9675 37354
rect 9731 37298 9817 37354
rect 9873 37298 9959 37354
rect 10015 37298 10101 37354
rect 10157 37298 10243 37354
rect 10299 37298 10385 37354
rect 10441 37298 10527 37354
rect 10583 37298 10669 37354
rect 10725 37298 10811 37354
rect 10867 37298 10953 37354
rect 11009 37298 11095 37354
rect 11151 37298 11237 37354
rect 11293 37298 11379 37354
rect 11435 37298 11521 37354
rect 11577 37298 11663 37354
rect 11719 37298 11805 37354
rect 11861 37298 11947 37354
rect 12003 37298 12089 37354
rect 12145 37298 12231 37354
rect 12287 37298 12373 37354
rect 12429 37298 12515 37354
rect 12571 37298 12657 37354
rect 12713 37298 12799 37354
rect 12855 37298 12941 37354
rect 12997 37298 13083 37354
rect 13139 37298 13225 37354
rect 13281 37298 13367 37354
rect 13423 37298 13509 37354
rect 13565 37298 13651 37354
rect 13707 37298 13793 37354
rect 13849 37298 13935 37354
rect 13991 37298 14077 37354
rect 14133 37298 14219 37354
rect 14275 37298 14361 37354
rect 14417 37298 14503 37354
rect 14559 37298 14645 37354
rect 14701 37298 14787 37354
rect 14843 37298 15000 37354
rect 0 37212 15000 37298
rect 0 37156 161 37212
rect 217 37156 303 37212
rect 359 37156 445 37212
rect 501 37156 587 37212
rect 643 37156 729 37212
rect 785 37156 871 37212
rect 927 37156 1013 37212
rect 1069 37156 1155 37212
rect 1211 37156 1297 37212
rect 1353 37156 1439 37212
rect 1495 37156 1581 37212
rect 1637 37156 1723 37212
rect 1779 37156 1865 37212
rect 1921 37156 2007 37212
rect 2063 37156 2149 37212
rect 2205 37156 2291 37212
rect 2347 37156 2433 37212
rect 2489 37156 2575 37212
rect 2631 37156 2717 37212
rect 2773 37156 2859 37212
rect 2915 37156 3001 37212
rect 3057 37156 3143 37212
rect 3199 37156 3285 37212
rect 3341 37156 3427 37212
rect 3483 37156 3569 37212
rect 3625 37156 3711 37212
rect 3767 37156 3853 37212
rect 3909 37156 3995 37212
rect 4051 37156 4137 37212
rect 4193 37156 4279 37212
rect 4335 37156 4421 37212
rect 4477 37156 4563 37212
rect 4619 37156 4705 37212
rect 4761 37156 4847 37212
rect 4903 37156 4989 37212
rect 5045 37156 5131 37212
rect 5187 37156 5273 37212
rect 5329 37156 5415 37212
rect 5471 37156 5557 37212
rect 5613 37156 5699 37212
rect 5755 37156 5841 37212
rect 5897 37156 5983 37212
rect 6039 37156 6125 37212
rect 6181 37156 6267 37212
rect 6323 37156 6409 37212
rect 6465 37156 6551 37212
rect 6607 37156 6693 37212
rect 6749 37156 6835 37212
rect 6891 37156 6977 37212
rect 7033 37156 7119 37212
rect 7175 37156 7261 37212
rect 7317 37156 7403 37212
rect 7459 37156 7545 37212
rect 7601 37156 7687 37212
rect 7743 37156 7829 37212
rect 7885 37156 7971 37212
rect 8027 37156 8113 37212
rect 8169 37156 8255 37212
rect 8311 37156 8397 37212
rect 8453 37156 8539 37212
rect 8595 37156 8681 37212
rect 8737 37156 8823 37212
rect 8879 37156 8965 37212
rect 9021 37156 9107 37212
rect 9163 37156 9249 37212
rect 9305 37156 9391 37212
rect 9447 37156 9533 37212
rect 9589 37156 9675 37212
rect 9731 37156 9817 37212
rect 9873 37156 9959 37212
rect 10015 37156 10101 37212
rect 10157 37156 10243 37212
rect 10299 37156 10385 37212
rect 10441 37156 10527 37212
rect 10583 37156 10669 37212
rect 10725 37156 10811 37212
rect 10867 37156 10953 37212
rect 11009 37156 11095 37212
rect 11151 37156 11237 37212
rect 11293 37156 11379 37212
rect 11435 37156 11521 37212
rect 11577 37156 11663 37212
rect 11719 37156 11805 37212
rect 11861 37156 11947 37212
rect 12003 37156 12089 37212
rect 12145 37156 12231 37212
rect 12287 37156 12373 37212
rect 12429 37156 12515 37212
rect 12571 37156 12657 37212
rect 12713 37156 12799 37212
rect 12855 37156 12941 37212
rect 12997 37156 13083 37212
rect 13139 37156 13225 37212
rect 13281 37156 13367 37212
rect 13423 37156 13509 37212
rect 13565 37156 13651 37212
rect 13707 37156 13793 37212
rect 13849 37156 13935 37212
rect 13991 37156 14077 37212
rect 14133 37156 14219 37212
rect 14275 37156 14361 37212
rect 14417 37156 14503 37212
rect 14559 37156 14645 37212
rect 14701 37156 14787 37212
rect 14843 37156 15000 37212
rect 0 37070 15000 37156
rect 0 37014 161 37070
rect 217 37014 303 37070
rect 359 37014 445 37070
rect 501 37014 587 37070
rect 643 37014 729 37070
rect 785 37014 871 37070
rect 927 37014 1013 37070
rect 1069 37014 1155 37070
rect 1211 37014 1297 37070
rect 1353 37014 1439 37070
rect 1495 37014 1581 37070
rect 1637 37014 1723 37070
rect 1779 37014 1865 37070
rect 1921 37014 2007 37070
rect 2063 37014 2149 37070
rect 2205 37014 2291 37070
rect 2347 37014 2433 37070
rect 2489 37014 2575 37070
rect 2631 37014 2717 37070
rect 2773 37014 2859 37070
rect 2915 37014 3001 37070
rect 3057 37014 3143 37070
rect 3199 37014 3285 37070
rect 3341 37014 3427 37070
rect 3483 37014 3569 37070
rect 3625 37014 3711 37070
rect 3767 37014 3853 37070
rect 3909 37014 3995 37070
rect 4051 37014 4137 37070
rect 4193 37014 4279 37070
rect 4335 37014 4421 37070
rect 4477 37014 4563 37070
rect 4619 37014 4705 37070
rect 4761 37014 4847 37070
rect 4903 37014 4989 37070
rect 5045 37014 5131 37070
rect 5187 37014 5273 37070
rect 5329 37014 5415 37070
rect 5471 37014 5557 37070
rect 5613 37014 5699 37070
rect 5755 37014 5841 37070
rect 5897 37014 5983 37070
rect 6039 37014 6125 37070
rect 6181 37014 6267 37070
rect 6323 37014 6409 37070
rect 6465 37014 6551 37070
rect 6607 37014 6693 37070
rect 6749 37014 6835 37070
rect 6891 37014 6977 37070
rect 7033 37014 7119 37070
rect 7175 37014 7261 37070
rect 7317 37014 7403 37070
rect 7459 37014 7545 37070
rect 7601 37014 7687 37070
rect 7743 37014 7829 37070
rect 7885 37014 7971 37070
rect 8027 37014 8113 37070
rect 8169 37014 8255 37070
rect 8311 37014 8397 37070
rect 8453 37014 8539 37070
rect 8595 37014 8681 37070
rect 8737 37014 8823 37070
rect 8879 37014 8965 37070
rect 9021 37014 9107 37070
rect 9163 37014 9249 37070
rect 9305 37014 9391 37070
rect 9447 37014 9533 37070
rect 9589 37014 9675 37070
rect 9731 37014 9817 37070
rect 9873 37014 9959 37070
rect 10015 37014 10101 37070
rect 10157 37014 10243 37070
rect 10299 37014 10385 37070
rect 10441 37014 10527 37070
rect 10583 37014 10669 37070
rect 10725 37014 10811 37070
rect 10867 37014 10953 37070
rect 11009 37014 11095 37070
rect 11151 37014 11237 37070
rect 11293 37014 11379 37070
rect 11435 37014 11521 37070
rect 11577 37014 11663 37070
rect 11719 37014 11805 37070
rect 11861 37014 11947 37070
rect 12003 37014 12089 37070
rect 12145 37014 12231 37070
rect 12287 37014 12373 37070
rect 12429 37014 12515 37070
rect 12571 37014 12657 37070
rect 12713 37014 12799 37070
rect 12855 37014 12941 37070
rect 12997 37014 13083 37070
rect 13139 37014 13225 37070
rect 13281 37014 13367 37070
rect 13423 37014 13509 37070
rect 13565 37014 13651 37070
rect 13707 37014 13793 37070
rect 13849 37014 13935 37070
rect 13991 37014 14077 37070
rect 14133 37014 14219 37070
rect 14275 37014 14361 37070
rect 14417 37014 14503 37070
rect 14559 37014 14645 37070
rect 14701 37014 14787 37070
rect 14843 37014 15000 37070
rect 0 36928 15000 37014
rect 0 36872 161 36928
rect 217 36872 303 36928
rect 359 36872 445 36928
rect 501 36872 587 36928
rect 643 36872 729 36928
rect 785 36872 871 36928
rect 927 36872 1013 36928
rect 1069 36872 1155 36928
rect 1211 36872 1297 36928
rect 1353 36872 1439 36928
rect 1495 36872 1581 36928
rect 1637 36872 1723 36928
rect 1779 36872 1865 36928
rect 1921 36872 2007 36928
rect 2063 36872 2149 36928
rect 2205 36872 2291 36928
rect 2347 36872 2433 36928
rect 2489 36872 2575 36928
rect 2631 36872 2717 36928
rect 2773 36872 2859 36928
rect 2915 36872 3001 36928
rect 3057 36872 3143 36928
rect 3199 36872 3285 36928
rect 3341 36872 3427 36928
rect 3483 36872 3569 36928
rect 3625 36872 3711 36928
rect 3767 36872 3853 36928
rect 3909 36872 3995 36928
rect 4051 36872 4137 36928
rect 4193 36872 4279 36928
rect 4335 36872 4421 36928
rect 4477 36872 4563 36928
rect 4619 36872 4705 36928
rect 4761 36872 4847 36928
rect 4903 36872 4989 36928
rect 5045 36872 5131 36928
rect 5187 36872 5273 36928
rect 5329 36872 5415 36928
rect 5471 36872 5557 36928
rect 5613 36872 5699 36928
rect 5755 36872 5841 36928
rect 5897 36872 5983 36928
rect 6039 36872 6125 36928
rect 6181 36872 6267 36928
rect 6323 36872 6409 36928
rect 6465 36872 6551 36928
rect 6607 36872 6693 36928
rect 6749 36872 6835 36928
rect 6891 36872 6977 36928
rect 7033 36872 7119 36928
rect 7175 36872 7261 36928
rect 7317 36872 7403 36928
rect 7459 36872 7545 36928
rect 7601 36872 7687 36928
rect 7743 36872 7829 36928
rect 7885 36872 7971 36928
rect 8027 36872 8113 36928
rect 8169 36872 8255 36928
rect 8311 36872 8397 36928
rect 8453 36872 8539 36928
rect 8595 36872 8681 36928
rect 8737 36872 8823 36928
rect 8879 36872 8965 36928
rect 9021 36872 9107 36928
rect 9163 36872 9249 36928
rect 9305 36872 9391 36928
rect 9447 36872 9533 36928
rect 9589 36872 9675 36928
rect 9731 36872 9817 36928
rect 9873 36872 9959 36928
rect 10015 36872 10101 36928
rect 10157 36872 10243 36928
rect 10299 36872 10385 36928
rect 10441 36872 10527 36928
rect 10583 36872 10669 36928
rect 10725 36872 10811 36928
rect 10867 36872 10953 36928
rect 11009 36872 11095 36928
rect 11151 36872 11237 36928
rect 11293 36872 11379 36928
rect 11435 36872 11521 36928
rect 11577 36872 11663 36928
rect 11719 36872 11805 36928
rect 11861 36872 11947 36928
rect 12003 36872 12089 36928
rect 12145 36872 12231 36928
rect 12287 36872 12373 36928
rect 12429 36872 12515 36928
rect 12571 36872 12657 36928
rect 12713 36872 12799 36928
rect 12855 36872 12941 36928
rect 12997 36872 13083 36928
rect 13139 36872 13225 36928
rect 13281 36872 13367 36928
rect 13423 36872 13509 36928
rect 13565 36872 13651 36928
rect 13707 36872 13793 36928
rect 13849 36872 13935 36928
rect 13991 36872 14077 36928
rect 14133 36872 14219 36928
rect 14275 36872 14361 36928
rect 14417 36872 14503 36928
rect 14559 36872 14645 36928
rect 14701 36872 14787 36928
rect 14843 36872 15000 36928
rect 0 36786 15000 36872
rect 0 36730 161 36786
rect 217 36730 303 36786
rect 359 36730 445 36786
rect 501 36730 587 36786
rect 643 36730 729 36786
rect 785 36730 871 36786
rect 927 36730 1013 36786
rect 1069 36730 1155 36786
rect 1211 36730 1297 36786
rect 1353 36730 1439 36786
rect 1495 36730 1581 36786
rect 1637 36730 1723 36786
rect 1779 36730 1865 36786
rect 1921 36730 2007 36786
rect 2063 36730 2149 36786
rect 2205 36730 2291 36786
rect 2347 36730 2433 36786
rect 2489 36730 2575 36786
rect 2631 36730 2717 36786
rect 2773 36730 2859 36786
rect 2915 36730 3001 36786
rect 3057 36730 3143 36786
rect 3199 36730 3285 36786
rect 3341 36730 3427 36786
rect 3483 36730 3569 36786
rect 3625 36730 3711 36786
rect 3767 36730 3853 36786
rect 3909 36730 3995 36786
rect 4051 36730 4137 36786
rect 4193 36730 4279 36786
rect 4335 36730 4421 36786
rect 4477 36730 4563 36786
rect 4619 36730 4705 36786
rect 4761 36730 4847 36786
rect 4903 36730 4989 36786
rect 5045 36730 5131 36786
rect 5187 36730 5273 36786
rect 5329 36730 5415 36786
rect 5471 36730 5557 36786
rect 5613 36730 5699 36786
rect 5755 36730 5841 36786
rect 5897 36730 5983 36786
rect 6039 36730 6125 36786
rect 6181 36730 6267 36786
rect 6323 36730 6409 36786
rect 6465 36730 6551 36786
rect 6607 36730 6693 36786
rect 6749 36730 6835 36786
rect 6891 36730 6977 36786
rect 7033 36730 7119 36786
rect 7175 36730 7261 36786
rect 7317 36730 7403 36786
rect 7459 36730 7545 36786
rect 7601 36730 7687 36786
rect 7743 36730 7829 36786
rect 7885 36730 7971 36786
rect 8027 36730 8113 36786
rect 8169 36730 8255 36786
rect 8311 36730 8397 36786
rect 8453 36730 8539 36786
rect 8595 36730 8681 36786
rect 8737 36730 8823 36786
rect 8879 36730 8965 36786
rect 9021 36730 9107 36786
rect 9163 36730 9249 36786
rect 9305 36730 9391 36786
rect 9447 36730 9533 36786
rect 9589 36730 9675 36786
rect 9731 36730 9817 36786
rect 9873 36730 9959 36786
rect 10015 36730 10101 36786
rect 10157 36730 10243 36786
rect 10299 36730 10385 36786
rect 10441 36730 10527 36786
rect 10583 36730 10669 36786
rect 10725 36730 10811 36786
rect 10867 36730 10953 36786
rect 11009 36730 11095 36786
rect 11151 36730 11237 36786
rect 11293 36730 11379 36786
rect 11435 36730 11521 36786
rect 11577 36730 11663 36786
rect 11719 36730 11805 36786
rect 11861 36730 11947 36786
rect 12003 36730 12089 36786
rect 12145 36730 12231 36786
rect 12287 36730 12373 36786
rect 12429 36730 12515 36786
rect 12571 36730 12657 36786
rect 12713 36730 12799 36786
rect 12855 36730 12941 36786
rect 12997 36730 13083 36786
rect 13139 36730 13225 36786
rect 13281 36730 13367 36786
rect 13423 36730 13509 36786
rect 13565 36730 13651 36786
rect 13707 36730 13793 36786
rect 13849 36730 13935 36786
rect 13991 36730 14077 36786
rect 14133 36730 14219 36786
rect 14275 36730 14361 36786
rect 14417 36730 14503 36786
rect 14559 36730 14645 36786
rect 14701 36730 14787 36786
rect 14843 36730 15000 36786
rect 0 36644 15000 36730
rect 0 36588 161 36644
rect 217 36588 303 36644
rect 359 36588 445 36644
rect 501 36588 587 36644
rect 643 36588 729 36644
rect 785 36588 871 36644
rect 927 36588 1013 36644
rect 1069 36588 1155 36644
rect 1211 36588 1297 36644
rect 1353 36588 1439 36644
rect 1495 36588 1581 36644
rect 1637 36588 1723 36644
rect 1779 36588 1865 36644
rect 1921 36588 2007 36644
rect 2063 36588 2149 36644
rect 2205 36588 2291 36644
rect 2347 36588 2433 36644
rect 2489 36588 2575 36644
rect 2631 36588 2717 36644
rect 2773 36588 2859 36644
rect 2915 36588 3001 36644
rect 3057 36588 3143 36644
rect 3199 36588 3285 36644
rect 3341 36588 3427 36644
rect 3483 36588 3569 36644
rect 3625 36588 3711 36644
rect 3767 36588 3853 36644
rect 3909 36588 3995 36644
rect 4051 36588 4137 36644
rect 4193 36588 4279 36644
rect 4335 36588 4421 36644
rect 4477 36588 4563 36644
rect 4619 36588 4705 36644
rect 4761 36588 4847 36644
rect 4903 36588 4989 36644
rect 5045 36588 5131 36644
rect 5187 36588 5273 36644
rect 5329 36588 5415 36644
rect 5471 36588 5557 36644
rect 5613 36588 5699 36644
rect 5755 36588 5841 36644
rect 5897 36588 5983 36644
rect 6039 36588 6125 36644
rect 6181 36588 6267 36644
rect 6323 36588 6409 36644
rect 6465 36588 6551 36644
rect 6607 36588 6693 36644
rect 6749 36588 6835 36644
rect 6891 36588 6977 36644
rect 7033 36588 7119 36644
rect 7175 36588 7261 36644
rect 7317 36588 7403 36644
rect 7459 36588 7545 36644
rect 7601 36588 7687 36644
rect 7743 36588 7829 36644
rect 7885 36588 7971 36644
rect 8027 36588 8113 36644
rect 8169 36588 8255 36644
rect 8311 36588 8397 36644
rect 8453 36588 8539 36644
rect 8595 36588 8681 36644
rect 8737 36588 8823 36644
rect 8879 36588 8965 36644
rect 9021 36588 9107 36644
rect 9163 36588 9249 36644
rect 9305 36588 9391 36644
rect 9447 36588 9533 36644
rect 9589 36588 9675 36644
rect 9731 36588 9817 36644
rect 9873 36588 9959 36644
rect 10015 36588 10101 36644
rect 10157 36588 10243 36644
rect 10299 36588 10385 36644
rect 10441 36588 10527 36644
rect 10583 36588 10669 36644
rect 10725 36588 10811 36644
rect 10867 36588 10953 36644
rect 11009 36588 11095 36644
rect 11151 36588 11237 36644
rect 11293 36588 11379 36644
rect 11435 36588 11521 36644
rect 11577 36588 11663 36644
rect 11719 36588 11805 36644
rect 11861 36588 11947 36644
rect 12003 36588 12089 36644
rect 12145 36588 12231 36644
rect 12287 36588 12373 36644
rect 12429 36588 12515 36644
rect 12571 36588 12657 36644
rect 12713 36588 12799 36644
rect 12855 36588 12941 36644
rect 12997 36588 13083 36644
rect 13139 36588 13225 36644
rect 13281 36588 13367 36644
rect 13423 36588 13509 36644
rect 13565 36588 13651 36644
rect 13707 36588 13793 36644
rect 13849 36588 13935 36644
rect 13991 36588 14077 36644
rect 14133 36588 14219 36644
rect 14275 36588 14361 36644
rect 14417 36588 14503 36644
rect 14559 36588 14645 36644
rect 14701 36588 14787 36644
rect 14843 36588 15000 36644
rect 0 36502 15000 36588
rect 0 36446 161 36502
rect 217 36446 303 36502
rect 359 36446 445 36502
rect 501 36446 587 36502
rect 643 36446 729 36502
rect 785 36446 871 36502
rect 927 36446 1013 36502
rect 1069 36446 1155 36502
rect 1211 36446 1297 36502
rect 1353 36446 1439 36502
rect 1495 36446 1581 36502
rect 1637 36446 1723 36502
rect 1779 36446 1865 36502
rect 1921 36446 2007 36502
rect 2063 36446 2149 36502
rect 2205 36446 2291 36502
rect 2347 36446 2433 36502
rect 2489 36446 2575 36502
rect 2631 36446 2717 36502
rect 2773 36446 2859 36502
rect 2915 36446 3001 36502
rect 3057 36446 3143 36502
rect 3199 36446 3285 36502
rect 3341 36446 3427 36502
rect 3483 36446 3569 36502
rect 3625 36446 3711 36502
rect 3767 36446 3853 36502
rect 3909 36446 3995 36502
rect 4051 36446 4137 36502
rect 4193 36446 4279 36502
rect 4335 36446 4421 36502
rect 4477 36446 4563 36502
rect 4619 36446 4705 36502
rect 4761 36446 4847 36502
rect 4903 36446 4989 36502
rect 5045 36446 5131 36502
rect 5187 36446 5273 36502
rect 5329 36446 5415 36502
rect 5471 36446 5557 36502
rect 5613 36446 5699 36502
rect 5755 36446 5841 36502
rect 5897 36446 5983 36502
rect 6039 36446 6125 36502
rect 6181 36446 6267 36502
rect 6323 36446 6409 36502
rect 6465 36446 6551 36502
rect 6607 36446 6693 36502
rect 6749 36446 6835 36502
rect 6891 36446 6977 36502
rect 7033 36446 7119 36502
rect 7175 36446 7261 36502
rect 7317 36446 7403 36502
rect 7459 36446 7545 36502
rect 7601 36446 7687 36502
rect 7743 36446 7829 36502
rect 7885 36446 7971 36502
rect 8027 36446 8113 36502
rect 8169 36446 8255 36502
rect 8311 36446 8397 36502
rect 8453 36446 8539 36502
rect 8595 36446 8681 36502
rect 8737 36446 8823 36502
rect 8879 36446 8965 36502
rect 9021 36446 9107 36502
rect 9163 36446 9249 36502
rect 9305 36446 9391 36502
rect 9447 36446 9533 36502
rect 9589 36446 9675 36502
rect 9731 36446 9817 36502
rect 9873 36446 9959 36502
rect 10015 36446 10101 36502
rect 10157 36446 10243 36502
rect 10299 36446 10385 36502
rect 10441 36446 10527 36502
rect 10583 36446 10669 36502
rect 10725 36446 10811 36502
rect 10867 36446 10953 36502
rect 11009 36446 11095 36502
rect 11151 36446 11237 36502
rect 11293 36446 11379 36502
rect 11435 36446 11521 36502
rect 11577 36446 11663 36502
rect 11719 36446 11805 36502
rect 11861 36446 11947 36502
rect 12003 36446 12089 36502
rect 12145 36446 12231 36502
rect 12287 36446 12373 36502
rect 12429 36446 12515 36502
rect 12571 36446 12657 36502
rect 12713 36446 12799 36502
rect 12855 36446 12941 36502
rect 12997 36446 13083 36502
rect 13139 36446 13225 36502
rect 13281 36446 13367 36502
rect 13423 36446 13509 36502
rect 13565 36446 13651 36502
rect 13707 36446 13793 36502
rect 13849 36446 13935 36502
rect 13991 36446 14077 36502
rect 14133 36446 14219 36502
rect 14275 36446 14361 36502
rect 14417 36446 14503 36502
rect 14559 36446 14645 36502
rect 14701 36446 14787 36502
rect 14843 36446 15000 36502
rect 0 36400 15000 36446
rect 937 36200 3937 36400
rect 4337 36200 7337 36400
rect 7737 36200 10737 36400
rect 11137 36200 14137 36400
rect 0 36142 15000 36200
rect 0 36086 161 36142
rect 217 36086 303 36142
rect 359 36086 445 36142
rect 501 36086 587 36142
rect 643 36086 729 36142
rect 785 36086 871 36142
rect 927 36086 1013 36142
rect 1069 36086 1155 36142
rect 1211 36086 1297 36142
rect 1353 36086 1439 36142
rect 1495 36086 1581 36142
rect 1637 36086 1723 36142
rect 1779 36086 1865 36142
rect 1921 36086 2007 36142
rect 2063 36086 2149 36142
rect 2205 36086 2291 36142
rect 2347 36086 2433 36142
rect 2489 36086 2575 36142
rect 2631 36086 2717 36142
rect 2773 36086 2859 36142
rect 2915 36086 3001 36142
rect 3057 36086 3143 36142
rect 3199 36086 3285 36142
rect 3341 36086 3427 36142
rect 3483 36086 3569 36142
rect 3625 36086 3711 36142
rect 3767 36086 3853 36142
rect 3909 36086 3995 36142
rect 4051 36086 4137 36142
rect 4193 36086 4279 36142
rect 4335 36086 4421 36142
rect 4477 36086 4563 36142
rect 4619 36086 4705 36142
rect 4761 36086 4847 36142
rect 4903 36086 4989 36142
rect 5045 36086 5131 36142
rect 5187 36086 5273 36142
rect 5329 36086 5415 36142
rect 5471 36086 5557 36142
rect 5613 36086 5699 36142
rect 5755 36086 5841 36142
rect 5897 36086 5983 36142
rect 6039 36086 6125 36142
rect 6181 36086 6267 36142
rect 6323 36086 6409 36142
rect 6465 36086 6551 36142
rect 6607 36086 6693 36142
rect 6749 36086 6835 36142
rect 6891 36086 6977 36142
rect 7033 36086 7119 36142
rect 7175 36086 7261 36142
rect 7317 36086 7403 36142
rect 7459 36086 7545 36142
rect 7601 36086 7687 36142
rect 7743 36086 7829 36142
rect 7885 36086 7971 36142
rect 8027 36086 8113 36142
rect 8169 36086 8255 36142
rect 8311 36086 8397 36142
rect 8453 36086 8539 36142
rect 8595 36086 8681 36142
rect 8737 36086 8823 36142
rect 8879 36086 8965 36142
rect 9021 36086 9107 36142
rect 9163 36086 9249 36142
rect 9305 36086 9391 36142
rect 9447 36086 9533 36142
rect 9589 36086 9675 36142
rect 9731 36086 9817 36142
rect 9873 36086 9959 36142
rect 10015 36086 10101 36142
rect 10157 36086 10243 36142
rect 10299 36086 10385 36142
rect 10441 36086 10527 36142
rect 10583 36086 10669 36142
rect 10725 36086 10811 36142
rect 10867 36086 10953 36142
rect 11009 36086 11095 36142
rect 11151 36086 11237 36142
rect 11293 36086 11379 36142
rect 11435 36086 11521 36142
rect 11577 36086 11663 36142
rect 11719 36086 11805 36142
rect 11861 36086 11947 36142
rect 12003 36086 12089 36142
rect 12145 36086 12231 36142
rect 12287 36086 12373 36142
rect 12429 36086 12515 36142
rect 12571 36086 12657 36142
rect 12713 36086 12799 36142
rect 12855 36086 12941 36142
rect 12997 36086 13083 36142
rect 13139 36086 13225 36142
rect 13281 36086 13367 36142
rect 13423 36086 13509 36142
rect 13565 36086 13651 36142
rect 13707 36086 13793 36142
rect 13849 36086 13935 36142
rect 13991 36086 14077 36142
rect 14133 36086 14219 36142
rect 14275 36086 14361 36142
rect 14417 36086 14503 36142
rect 14559 36086 14645 36142
rect 14701 36086 14787 36142
rect 14843 36086 15000 36142
rect 0 36000 15000 36086
rect 0 35944 161 36000
rect 217 35944 303 36000
rect 359 35944 445 36000
rect 501 35944 587 36000
rect 643 35944 729 36000
rect 785 35944 871 36000
rect 927 35944 1013 36000
rect 1069 35944 1155 36000
rect 1211 35944 1297 36000
rect 1353 35944 1439 36000
rect 1495 35944 1581 36000
rect 1637 35944 1723 36000
rect 1779 35944 1865 36000
rect 1921 35944 2007 36000
rect 2063 35944 2149 36000
rect 2205 35944 2291 36000
rect 2347 35944 2433 36000
rect 2489 35944 2575 36000
rect 2631 35944 2717 36000
rect 2773 35944 2859 36000
rect 2915 35944 3001 36000
rect 3057 35944 3143 36000
rect 3199 35944 3285 36000
rect 3341 35944 3427 36000
rect 3483 35944 3569 36000
rect 3625 35944 3711 36000
rect 3767 35944 3853 36000
rect 3909 35944 3995 36000
rect 4051 35944 4137 36000
rect 4193 35944 4279 36000
rect 4335 35944 4421 36000
rect 4477 35944 4563 36000
rect 4619 35944 4705 36000
rect 4761 35944 4847 36000
rect 4903 35944 4989 36000
rect 5045 35944 5131 36000
rect 5187 35944 5273 36000
rect 5329 35944 5415 36000
rect 5471 35944 5557 36000
rect 5613 35944 5699 36000
rect 5755 35944 5841 36000
rect 5897 35944 5983 36000
rect 6039 35944 6125 36000
rect 6181 35944 6267 36000
rect 6323 35944 6409 36000
rect 6465 35944 6551 36000
rect 6607 35944 6693 36000
rect 6749 35944 6835 36000
rect 6891 35944 6977 36000
rect 7033 35944 7119 36000
rect 7175 35944 7261 36000
rect 7317 35944 7403 36000
rect 7459 35944 7545 36000
rect 7601 35944 7687 36000
rect 7743 35944 7829 36000
rect 7885 35944 7971 36000
rect 8027 35944 8113 36000
rect 8169 35944 8255 36000
rect 8311 35944 8397 36000
rect 8453 35944 8539 36000
rect 8595 35944 8681 36000
rect 8737 35944 8823 36000
rect 8879 35944 8965 36000
rect 9021 35944 9107 36000
rect 9163 35944 9249 36000
rect 9305 35944 9391 36000
rect 9447 35944 9533 36000
rect 9589 35944 9675 36000
rect 9731 35944 9817 36000
rect 9873 35944 9959 36000
rect 10015 35944 10101 36000
rect 10157 35944 10243 36000
rect 10299 35944 10385 36000
rect 10441 35944 10527 36000
rect 10583 35944 10669 36000
rect 10725 35944 10811 36000
rect 10867 35944 10953 36000
rect 11009 35944 11095 36000
rect 11151 35944 11237 36000
rect 11293 35944 11379 36000
rect 11435 35944 11521 36000
rect 11577 35944 11663 36000
rect 11719 35944 11805 36000
rect 11861 35944 11947 36000
rect 12003 35944 12089 36000
rect 12145 35944 12231 36000
rect 12287 35944 12373 36000
rect 12429 35944 12515 36000
rect 12571 35944 12657 36000
rect 12713 35944 12799 36000
rect 12855 35944 12941 36000
rect 12997 35944 13083 36000
rect 13139 35944 13225 36000
rect 13281 35944 13367 36000
rect 13423 35944 13509 36000
rect 13565 35944 13651 36000
rect 13707 35944 13793 36000
rect 13849 35944 13935 36000
rect 13991 35944 14077 36000
rect 14133 35944 14219 36000
rect 14275 35944 14361 36000
rect 14417 35944 14503 36000
rect 14559 35944 14645 36000
rect 14701 35944 14787 36000
rect 14843 35944 15000 36000
rect 0 35858 15000 35944
rect 0 35802 161 35858
rect 217 35802 303 35858
rect 359 35802 445 35858
rect 501 35802 587 35858
rect 643 35802 729 35858
rect 785 35802 871 35858
rect 927 35802 1013 35858
rect 1069 35802 1155 35858
rect 1211 35802 1297 35858
rect 1353 35802 1439 35858
rect 1495 35802 1581 35858
rect 1637 35802 1723 35858
rect 1779 35802 1865 35858
rect 1921 35802 2007 35858
rect 2063 35802 2149 35858
rect 2205 35802 2291 35858
rect 2347 35802 2433 35858
rect 2489 35802 2575 35858
rect 2631 35802 2717 35858
rect 2773 35802 2859 35858
rect 2915 35802 3001 35858
rect 3057 35802 3143 35858
rect 3199 35802 3285 35858
rect 3341 35802 3427 35858
rect 3483 35802 3569 35858
rect 3625 35802 3711 35858
rect 3767 35802 3853 35858
rect 3909 35802 3995 35858
rect 4051 35802 4137 35858
rect 4193 35802 4279 35858
rect 4335 35802 4421 35858
rect 4477 35802 4563 35858
rect 4619 35802 4705 35858
rect 4761 35802 4847 35858
rect 4903 35802 4989 35858
rect 5045 35802 5131 35858
rect 5187 35802 5273 35858
rect 5329 35802 5415 35858
rect 5471 35802 5557 35858
rect 5613 35802 5699 35858
rect 5755 35802 5841 35858
rect 5897 35802 5983 35858
rect 6039 35802 6125 35858
rect 6181 35802 6267 35858
rect 6323 35802 6409 35858
rect 6465 35802 6551 35858
rect 6607 35802 6693 35858
rect 6749 35802 6835 35858
rect 6891 35802 6977 35858
rect 7033 35802 7119 35858
rect 7175 35802 7261 35858
rect 7317 35802 7403 35858
rect 7459 35802 7545 35858
rect 7601 35802 7687 35858
rect 7743 35802 7829 35858
rect 7885 35802 7971 35858
rect 8027 35802 8113 35858
rect 8169 35802 8255 35858
rect 8311 35802 8397 35858
rect 8453 35802 8539 35858
rect 8595 35802 8681 35858
rect 8737 35802 8823 35858
rect 8879 35802 8965 35858
rect 9021 35802 9107 35858
rect 9163 35802 9249 35858
rect 9305 35802 9391 35858
rect 9447 35802 9533 35858
rect 9589 35802 9675 35858
rect 9731 35802 9817 35858
rect 9873 35802 9959 35858
rect 10015 35802 10101 35858
rect 10157 35802 10243 35858
rect 10299 35802 10385 35858
rect 10441 35802 10527 35858
rect 10583 35802 10669 35858
rect 10725 35802 10811 35858
rect 10867 35802 10953 35858
rect 11009 35802 11095 35858
rect 11151 35802 11237 35858
rect 11293 35802 11379 35858
rect 11435 35802 11521 35858
rect 11577 35802 11663 35858
rect 11719 35802 11805 35858
rect 11861 35802 11947 35858
rect 12003 35802 12089 35858
rect 12145 35802 12231 35858
rect 12287 35802 12373 35858
rect 12429 35802 12515 35858
rect 12571 35802 12657 35858
rect 12713 35802 12799 35858
rect 12855 35802 12941 35858
rect 12997 35802 13083 35858
rect 13139 35802 13225 35858
rect 13281 35802 13367 35858
rect 13423 35802 13509 35858
rect 13565 35802 13651 35858
rect 13707 35802 13793 35858
rect 13849 35802 13935 35858
rect 13991 35802 14077 35858
rect 14133 35802 14219 35858
rect 14275 35802 14361 35858
rect 14417 35802 14503 35858
rect 14559 35802 14645 35858
rect 14701 35802 14787 35858
rect 14843 35802 15000 35858
rect 0 35716 15000 35802
rect 0 35660 161 35716
rect 217 35660 303 35716
rect 359 35660 445 35716
rect 501 35660 587 35716
rect 643 35660 729 35716
rect 785 35660 871 35716
rect 927 35660 1013 35716
rect 1069 35660 1155 35716
rect 1211 35660 1297 35716
rect 1353 35660 1439 35716
rect 1495 35660 1581 35716
rect 1637 35660 1723 35716
rect 1779 35660 1865 35716
rect 1921 35660 2007 35716
rect 2063 35660 2149 35716
rect 2205 35660 2291 35716
rect 2347 35660 2433 35716
rect 2489 35660 2575 35716
rect 2631 35660 2717 35716
rect 2773 35660 2859 35716
rect 2915 35660 3001 35716
rect 3057 35660 3143 35716
rect 3199 35660 3285 35716
rect 3341 35660 3427 35716
rect 3483 35660 3569 35716
rect 3625 35660 3711 35716
rect 3767 35660 3853 35716
rect 3909 35660 3995 35716
rect 4051 35660 4137 35716
rect 4193 35660 4279 35716
rect 4335 35660 4421 35716
rect 4477 35660 4563 35716
rect 4619 35660 4705 35716
rect 4761 35660 4847 35716
rect 4903 35660 4989 35716
rect 5045 35660 5131 35716
rect 5187 35660 5273 35716
rect 5329 35660 5415 35716
rect 5471 35660 5557 35716
rect 5613 35660 5699 35716
rect 5755 35660 5841 35716
rect 5897 35660 5983 35716
rect 6039 35660 6125 35716
rect 6181 35660 6267 35716
rect 6323 35660 6409 35716
rect 6465 35660 6551 35716
rect 6607 35660 6693 35716
rect 6749 35660 6835 35716
rect 6891 35660 6977 35716
rect 7033 35660 7119 35716
rect 7175 35660 7261 35716
rect 7317 35660 7403 35716
rect 7459 35660 7545 35716
rect 7601 35660 7687 35716
rect 7743 35660 7829 35716
rect 7885 35660 7971 35716
rect 8027 35660 8113 35716
rect 8169 35660 8255 35716
rect 8311 35660 8397 35716
rect 8453 35660 8539 35716
rect 8595 35660 8681 35716
rect 8737 35660 8823 35716
rect 8879 35660 8965 35716
rect 9021 35660 9107 35716
rect 9163 35660 9249 35716
rect 9305 35660 9391 35716
rect 9447 35660 9533 35716
rect 9589 35660 9675 35716
rect 9731 35660 9817 35716
rect 9873 35660 9959 35716
rect 10015 35660 10101 35716
rect 10157 35660 10243 35716
rect 10299 35660 10385 35716
rect 10441 35660 10527 35716
rect 10583 35660 10669 35716
rect 10725 35660 10811 35716
rect 10867 35660 10953 35716
rect 11009 35660 11095 35716
rect 11151 35660 11237 35716
rect 11293 35660 11379 35716
rect 11435 35660 11521 35716
rect 11577 35660 11663 35716
rect 11719 35660 11805 35716
rect 11861 35660 11947 35716
rect 12003 35660 12089 35716
rect 12145 35660 12231 35716
rect 12287 35660 12373 35716
rect 12429 35660 12515 35716
rect 12571 35660 12657 35716
rect 12713 35660 12799 35716
rect 12855 35660 12941 35716
rect 12997 35660 13083 35716
rect 13139 35660 13225 35716
rect 13281 35660 13367 35716
rect 13423 35660 13509 35716
rect 13565 35660 13651 35716
rect 13707 35660 13793 35716
rect 13849 35660 13935 35716
rect 13991 35660 14077 35716
rect 14133 35660 14219 35716
rect 14275 35660 14361 35716
rect 14417 35660 14503 35716
rect 14559 35660 14645 35716
rect 14701 35660 14787 35716
rect 14843 35660 15000 35716
rect 0 35574 15000 35660
rect 0 35518 161 35574
rect 217 35518 303 35574
rect 359 35518 445 35574
rect 501 35518 587 35574
rect 643 35518 729 35574
rect 785 35518 871 35574
rect 927 35518 1013 35574
rect 1069 35518 1155 35574
rect 1211 35518 1297 35574
rect 1353 35518 1439 35574
rect 1495 35518 1581 35574
rect 1637 35518 1723 35574
rect 1779 35518 1865 35574
rect 1921 35518 2007 35574
rect 2063 35518 2149 35574
rect 2205 35518 2291 35574
rect 2347 35518 2433 35574
rect 2489 35518 2575 35574
rect 2631 35518 2717 35574
rect 2773 35518 2859 35574
rect 2915 35518 3001 35574
rect 3057 35518 3143 35574
rect 3199 35518 3285 35574
rect 3341 35518 3427 35574
rect 3483 35518 3569 35574
rect 3625 35518 3711 35574
rect 3767 35518 3853 35574
rect 3909 35518 3995 35574
rect 4051 35518 4137 35574
rect 4193 35518 4279 35574
rect 4335 35518 4421 35574
rect 4477 35518 4563 35574
rect 4619 35518 4705 35574
rect 4761 35518 4847 35574
rect 4903 35518 4989 35574
rect 5045 35518 5131 35574
rect 5187 35518 5273 35574
rect 5329 35518 5415 35574
rect 5471 35518 5557 35574
rect 5613 35518 5699 35574
rect 5755 35518 5841 35574
rect 5897 35518 5983 35574
rect 6039 35518 6125 35574
rect 6181 35518 6267 35574
rect 6323 35518 6409 35574
rect 6465 35518 6551 35574
rect 6607 35518 6693 35574
rect 6749 35518 6835 35574
rect 6891 35518 6977 35574
rect 7033 35518 7119 35574
rect 7175 35518 7261 35574
rect 7317 35518 7403 35574
rect 7459 35518 7545 35574
rect 7601 35518 7687 35574
rect 7743 35518 7829 35574
rect 7885 35518 7971 35574
rect 8027 35518 8113 35574
rect 8169 35518 8255 35574
rect 8311 35518 8397 35574
rect 8453 35518 8539 35574
rect 8595 35518 8681 35574
rect 8737 35518 8823 35574
rect 8879 35518 8965 35574
rect 9021 35518 9107 35574
rect 9163 35518 9249 35574
rect 9305 35518 9391 35574
rect 9447 35518 9533 35574
rect 9589 35518 9675 35574
rect 9731 35518 9817 35574
rect 9873 35518 9959 35574
rect 10015 35518 10101 35574
rect 10157 35518 10243 35574
rect 10299 35518 10385 35574
rect 10441 35518 10527 35574
rect 10583 35518 10669 35574
rect 10725 35518 10811 35574
rect 10867 35518 10953 35574
rect 11009 35518 11095 35574
rect 11151 35518 11237 35574
rect 11293 35518 11379 35574
rect 11435 35518 11521 35574
rect 11577 35518 11663 35574
rect 11719 35518 11805 35574
rect 11861 35518 11947 35574
rect 12003 35518 12089 35574
rect 12145 35518 12231 35574
rect 12287 35518 12373 35574
rect 12429 35518 12515 35574
rect 12571 35518 12657 35574
rect 12713 35518 12799 35574
rect 12855 35518 12941 35574
rect 12997 35518 13083 35574
rect 13139 35518 13225 35574
rect 13281 35518 13367 35574
rect 13423 35518 13509 35574
rect 13565 35518 13651 35574
rect 13707 35518 13793 35574
rect 13849 35518 13935 35574
rect 13991 35518 14077 35574
rect 14133 35518 14219 35574
rect 14275 35518 14361 35574
rect 14417 35518 14503 35574
rect 14559 35518 14645 35574
rect 14701 35518 14787 35574
rect 14843 35518 15000 35574
rect 0 35432 15000 35518
rect 0 35376 161 35432
rect 217 35376 303 35432
rect 359 35376 445 35432
rect 501 35376 587 35432
rect 643 35376 729 35432
rect 785 35376 871 35432
rect 927 35376 1013 35432
rect 1069 35376 1155 35432
rect 1211 35376 1297 35432
rect 1353 35376 1439 35432
rect 1495 35376 1581 35432
rect 1637 35376 1723 35432
rect 1779 35376 1865 35432
rect 1921 35376 2007 35432
rect 2063 35376 2149 35432
rect 2205 35376 2291 35432
rect 2347 35376 2433 35432
rect 2489 35376 2575 35432
rect 2631 35376 2717 35432
rect 2773 35376 2859 35432
rect 2915 35376 3001 35432
rect 3057 35376 3143 35432
rect 3199 35376 3285 35432
rect 3341 35376 3427 35432
rect 3483 35376 3569 35432
rect 3625 35376 3711 35432
rect 3767 35376 3853 35432
rect 3909 35376 3995 35432
rect 4051 35376 4137 35432
rect 4193 35376 4279 35432
rect 4335 35376 4421 35432
rect 4477 35376 4563 35432
rect 4619 35376 4705 35432
rect 4761 35376 4847 35432
rect 4903 35376 4989 35432
rect 5045 35376 5131 35432
rect 5187 35376 5273 35432
rect 5329 35376 5415 35432
rect 5471 35376 5557 35432
rect 5613 35376 5699 35432
rect 5755 35376 5841 35432
rect 5897 35376 5983 35432
rect 6039 35376 6125 35432
rect 6181 35376 6267 35432
rect 6323 35376 6409 35432
rect 6465 35376 6551 35432
rect 6607 35376 6693 35432
rect 6749 35376 6835 35432
rect 6891 35376 6977 35432
rect 7033 35376 7119 35432
rect 7175 35376 7261 35432
rect 7317 35376 7403 35432
rect 7459 35376 7545 35432
rect 7601 35376 7687 35432
rect 7743 35376 7829 35432
rect 7885 35376 7971 35432
rect 8027 35376 8113 35432
rect 8169 35376 8255 35432
rect 8311 35376 8397 35432
rect 8453 35376 8539 35432
rect 8595 35376 8681 35432
rect 8737 35376 8823 35432
rect 8879 35376 8965 35432
rect 9021 35376 9107 35432
rect 9163 35376 9249 35432
rect 9305 35376 9391 35432
rect 9447 35376 9533 35432
rect 9589 35376 9675 35432
rect 9731 35376 9817 35432
rect 9873 35376 9959 35432
rect 10015 35376 10101 35432
rect 10157 35376 10243 35432
rect 10299 35376 10385 35432
rect 10441 35376 10527 35432
rect 10583 35376 10669 35432
rect 10725 35376 10811 35432
rect 10867 35376 10953 35432
rect 11009 35376 11095 35432
rect 11151 35376 11237 35432
rect 11293 35376 11379 35432
rect 11435 35376 11521 35432
rect 11577 35376 11663 35432
rect 11719 35376 11805 35432
rect 11861 35376 11947 35432
rect 12003 35376 12089 35432
rect 12145 35376 12231 35432
rect 12287 35376 12373 35432
rect 12429 35376 12515 35432
rect 12571 35376 12657 35432
rect 12713 35376 12799 35432
rect 12855 35376 12941 35432
rect 12997 35376 13083 35432
rect 13139 35376 13225 35432
rect 13281 35376 13367 35432
rect 13423 35376 13509 35432
rect 13565 35376 13651 35432
rect 13707 35376 13793 35432
rect 13849 35376 13935 35432
rect 13991 35376 14077 35432
rect 14133 35376 14219 35432
rect 14275 35376 14361 35432
rect 14417 35376 14503 35432
rect 14559 35376 14645 35432
rect 14701 35376 14787 35432
rect 14843 35376 15000 35432
rect 0 35290 15000 35376
rect 0 35234 161 35290
rect 217 35234 303 35290
rect 359 35234 445 35290
rect 501 35234 587 35290
rect 643 35234 729 35290
rect 785 35234 871 35290
rect 927 35234 1013 35290
rect 1069 35234 1155 35290
rect 1211 35234 1297 35290
rect 1353 35234 1439 35290
rect 1495 35234 1581 35290
rect 1637 35234 1723 35290
rect 1779 35234 1865 35290
rect 1921 35234 2007 35290
rect 2063 35234 2149 35290
rect 2205 35234 2291 35290
rect 2347 35234 2433 35290
rect 2489 35234 2575 35290
rect 2631 35234 2717 35290
rect 2773 35234 2859 35290
rect 2915 35234 3001 35290
rect 3057 35234 3143 35290
rect 3199 35234 3285 35290
rect 3341 35234 3427 35290
rect 3483 35234 3569 35290
rect 3625 35234 3711 35290
rect 3767 35234 3853 35290
rect 3909 35234 3995 35290
rect 4051 35234 4137 35290
rect 4193 35234 4279 35290
rect 4335 35234 4421 35290
rect 4477 35234 4563 35290
rect 4619 35234 4705 35290
rect 4761 35234 4847 35290
rect 4903 35234 4989 35290
rect 5045 35234 5131 35290
rect 5187 35234 5273 35290
rect 5329 35234 5415 35290
rect 5471 35234 5557 35290
rect 5613 35234 5699 35290
rect 5755 35234 5841 35290
rect 5897 35234 5983 35290
rect 6039 35234 6125 35290
rect 6181 35234 6267 35290
rect 6323 35234 6409 35290
rect 6465 35234 6551 35290
rect 6607 35234 6693 35290
rect 6749 35234 6835 35290
rect 6891 35234 6977 35290
rect 7033 35234 7119 35290
rect 7175 35234 7261 35290
rect 7317 35234 7403 35290
rect 7459 35234 7545 35290
rect 7601 35234 7687 35290
rect 7743 35234 7829 35290
rect 7885 35234 7971 35290
rect 8027 35234 8113 35290
rect 8169 35234 8255 35290
rect 8311 35234 8397 35290
rect 8453 35234 8539 35290
rect 8595 35234 8681 35290
rect 8737 35234 8823 35290
rect 8879 35234 8965 35290
rect 9021 35234 9107 35290
rect 9163 35234 9249 35290
rect 9305 35234 9391 35290
rect 9447 35234 9533 35290
rect 9589 35234 9675 35290
rect 9731 35234 9817 35290
rect 9873 35234 9959 35290
rect 10015 35234 10101 35290
rect 10157 35234 10243 35290
rect 10299 35234 10385 35290
rect 10441 35234 10527 35290
rect 10583 35234 10669 35290
rect 10725 35234 10811 35290
rect 10867 35234 10953 35290
rect 11009 35234 11095 35290
rect 11151 35234 11237 35290
rect 11293 35234 11379 35290
rect 11435 35234 11521 35290
rect 11577 35234 11663 35290
rect 11719 35234 11805 35290
rect 11861 35234 11947 35290
rect 12003 35234 12089 35290
rect 12145 35234 12231 35290
rect 12287 35234 12373 35290
rect 12429 35234 12515 35290
rect 12571 35234 12657 35290
rect 12713 35234 12799 35290
rect 12855 35234 12941 35290
rect 12997 35234 13083 35290
rect 13139 35234 13225 35290
rect 13281 35234 13367 35290
rect 13423 35234 13509 35290
rect 13565 35234 13651 35290
rect 13707 35234 13793 35290
rect 13849 35234 13935 35290
rect 13991 35234 14077 35290
rect 14133 35234 14219 35290
rect 14275 35234 14361 35290
rect 14417 35234 14503 35290
rect 14559 35234 14645 35290
rect 14701 35234 14787 35290
rect 14843 35234 15000 35290
rect 0 35148 15000 35234
rect 0 35092 161 35148
rect 217 35092 303 35148
rect 359 35092 445 35148
rect 501 35092 587 35148
rect 643 35092 729 35148
rect 785 35092 871 35148
rect 927 35092 1013 35148
rect 1069 35092 1155 35148
rect 1211 35092 1297 35148
rect 1353 35092 1439 35148
rect 1495 35092 1581 35148
rect 1637 35092 1723 35148
rect 1779 35092 1865 35148
rect 1921 35092 2007 35148
rect 2063 35092 2149 35148
rect 2205 35092 2291 35148
rect 2347 35092 2433 35148
rect 2489 35092 2575 35148
rect 2631 35092 2717 35148
rect 2773 35092 2859 35148
rect 2915 35092 3001 35148
rect 3057 35092 3143 35148
rect 3199 35092 3285 35148
rect 3341 35092 3427 35148
rect 3483 35092 3569 35148
rect 3625 35092 3711 35148
rect 3767 35092 3853 35148
rect 3909 35092 3995 35148
rect 4051 35092 4137 35148
rect 4193 35092 4279 35148
rect 4335 35092 4421 35148
rect 4477 35092 4563 35148
rect 4619 35092 4705 35148
rect 4761 35092 4847 35148
rect 4903 35092 4989 35148
rect 5045 35092 5131 35148
rect 5187 35092 5273 35148
rect 5329 35092 5415 35148
rect 5471 35092 5557 35148
rect 5613 35092 5699 35148
rect 5755 35092 5841 35148
rect 5897 35092 5983 35148
rect 6039 35092 6125 35148
rect 6181 35092 6267 35148
rect 6323 35092 6409 35148
rect 6465 35092 6551 35148
rect 6607 35092 6693 35148
rect 6749 35092 6835 35148
rect 6891 35092 6977 35148
rect 7033 35092 7119 35148
rect 7175 35092 7261 35148
rect 7317 35092 7403 35148
rect 7459 35092 7545 35148
rect 7601 35092 7687 35148
rect 7743 35092 7829 35148
rect 7885 35092 7971 35148
rect 8027 35092 8113 35148
rect 8169 35092 8255 35148
rect 8311 35092 8397 35148
rect 8453 35092 8539 35148
rect 8595 35092 8681 35148
rect 8737 35092 8823 35148
rect 8879 35092 8965 35148
rect 9021 35092 9107 35148
rect 9163 35092 9249 35148
rect 9305 35092 9391 35148
rect 9447 35092 9533 35148
rect 9589 35092 9675 35148
rect 9731 35092 9817 35148
rect 9873 35092 9959 35148
rect 10015 35092 10101 35148
rect 10157 35092 10243 35148
rect 10299 35092 10385 35148
rect 10441 35092 10527 35148
rect 10583 35092 10669 35148
rect 10725 35092 10811 35148
rect 10867 35092 10953 35148
rect 11009 35092 11095 35148
rect 11151 35092 11237 35148
rect 11293 35092 11379 35148
rect 11435 35092 11521 35148
rect 11577 35092 11663 35148
rect 11719 35092 11805 35148
rect 11861 35092 11947 35148
rect 12003 35092 12089 35148
rect 12145 35092 12231 35148
rect 12287 35092 12373 35148
rect 12429 35092 12515 35148
rect 12571 35092 12657 35148
rect 12713 35092 12799 35148
rect 12855 35092 12941 35148
rect 12997 35092 13083 35148
rect 13139 35092 13225 35148
rect 13281 35092 13367 35148
rect 13423 35092 13509 35148
rect 13565 35092 13651 35148
rect 13707 35092 13793 35148
rect 13849 35092 13935 35148
rect 13991 35092 14077 35148
rect 14133 35092 14219 35148
rect 14275 35092 14361 35148
rect 14417 35092 14503 35148
rect 14559 35092 14645 35148
rect 14701 35092 14787 35148
rect 14843 35092 15000 35148
rect 0 35006 15000 35092
rect 0 34950 161 35006
rect 217 34950 303 35006
rect 359 34950 445 35006
rect 501 34950 587 35006
rect 643 34950 729 35006
rect 785 34950 871 35006
rect 927 34950 1013 35006
rect 1069 34950 1155 35006
rect 1211 34950 1297 35006
rect 1353 34950 1439 35006
rect 1495 34950 1581 35006
rect 1637 34950 1723 35006
rect 1779 34950 1865 35006
rect 1921 34950 2007 35006
rect 2063 34950 2149 35006
rect 2205 34950 2291 35006
rect 2347 34950 2433 35006
rect 2489 34950 2575 35006
rect 2631 34950 2717 35006
rect 2773 34950 2859 35006
rect 2915 34950 3001 35006
rect 3057 34950 3143 35006
rect 3199 34950 3285 35006
rect 3341 34950 3427 35006
rect 3483 34950 3569 35006
rect 3625 34950 3711 35006
rect 3767 34950 3853 35006
rect 3909 34950 3995 35006
rect 4051 34950 4137 35006
rect 4193 34950 4279 35006
rect 4335 34950 4421 35006
rect 4477 34950 4563 35006
rect 4619 34950 4705 35006
rect 4761 34950 4847 35006
rect 4903 34950 4989 35006
rect 5045 34950 5131 35006
rect 5187 34950 5273 35006
rect 5329 34950 5415 35006
rect 5471 34950 5557 35006
rect 5613 34950 5699 35006
rect 5755 34950 5841 35006
rect 5897 34950 5983 35006
rect 6039 34950 6125 35006
rect 6181 34950 6267 35006
rect 6323 34950 6409 35006
rect 6465 34950 6551 35006
rect 6607 34950 6693 35006
rect 6749 34950 6835 35006
rect 6891 34950 6977 35006
rect 7033 34950 7119 35006
rect 7175 34950 7261 35006
rect 7317 34950 7403 35006
rect 7459 34950 7545 35006
rect 7601 34950 7687 35006
rect 7743 34950 7829 35006
rect 7885 34950 7971 35006
rect 8027 34950 8113 35006
rect 8169 34950 8255 35006
rect 8311 34950 8397 35006
rect 8453 34950 8539 35006
rect 8595 34950 8681 35006
rect 8737 34950 8823 35006
rect 8879 34950 8965 35006
rect 9021 34950 9107 35006
rect 9163 34950 9249 35006
rect 9305 34950 9391 35006
rect 9447 34950 9533 35006
rect 9589 34950 9675 35006
rect 9731 34950 9817 35006
rect 9873 34950 9959 35006
rect 10015 34950 10101 35006
rect 10157 34950 10243 35006
rect 10299 34950 10385 35006
rect 10441 34950 10527 35006
rect 10583 34950 10669 35006
rect 10725 34950 10811 35006
rect 10867 34950 10953 35006
rect 11009 34950 11095 35006
rect 11151 34950 11237 35006
rect 11293 34950 11379 35006
rect 11435 34950 11521 35006
rect 11577 34950 11663 35006
rect 11719 34950 11805 35006
rect 11861 34950 11947 35006
rect 12003 34950 12089 35006
rect 12145 34950 12231 35006
rect 12287 34950 12373 35006
rect 12429 34950 12515 35006
rect 12571 34950 12657 35006
rect 12713 34950 12799 35006
rect 12855 34950 12941 35006
rect 12997 34950 13083 35006
rect 13139 34950 13225 35006
rect 13281 34950 13367 35006
rect 13423 34950 13509 35006
rect 13565 34950 13651 35006
rect 13707 34950 13793 35006
rect 13849 34950 13935 35006
rect 13991 34950 14077 35006
rect 14133 34950 14219 35006
rect 14275 34950 14361 35006
rect 14417 34950 14503 35006
rect 14559 34950 14645 35006
rect 14701 34950 14787 35006
rect 14843 34950 15000 35006
rect 0 34864 15000 34950
rect 0 34808 161 34864
rect 217 34808 303 34864
rect 359 34808 445 34864
rect 501 34808 587 34864
rect 643 34808 729 34864
rect 785 34808 871 34864
rect 927 34808 1013 34864
rect 1069 34808 1155 34864
rect 1211 34808 1297 34864
rect 1353 34808 1439 34864
rect 1495 34808 1581 34864
rect 1637 34808 1723 34864
rect 1779 34808 1865 34864
rect 1921 34808 2007 34864
rect 2063 34808 2149 34864
rect 2205 34808 2291 34864
rect 2347 34808 2433 34864
rect 2489 34808 2575 34864
rect 2631 34808 2717 34864
rect 2773 34808 2859 34864
rect 2915 34808 3001 34864
rect 3057 34808 3143 34864
rect 3199 34808 3285 34864
rect 3341 34808 3427 34864
rect 3483 34808 3569 34864
rect 3625 34808 3711 34864
rect 3767 34808 3853 34864
rect 3909 34808 3995 34864
rect 4051 34808 4137 34864
rect 4193 34808 4279 34864
rect 4335 34808 4421 34864
rect 4477 34808 4563 34864
rect 4619 34808 4705 34864
rect 4761 34808 4847 34864
rect 4903 34808 4989 34864
rect 5045 34808 5131 34864
rect 5187 34808 5273 34864
rect 5329 34808 5415 34864
rect 5471 34808 5557 34864
rect 5613 34808 5699 34864
rect 5755 34808 5841 34864
rect 5897 34808 5983 34864
rect 6039 34808 6125 34864
rect 6181 34808 6267 34864
rect 6323 34808 6409 34864
rect 6465 34808 6551 34864
rect 6607 34808 6693 34864
rect 6749 34808 6835 34864
rect 6891 34808 6977 34864
rect 7033 34808 7119 34864
rect 7175 34808 7261 34864
rect 7317 34808 7403 34864
rect 7459 34808 7545 34864
rect 7601 34808 7687 34864
rect 7743 34808 7829 34864
rect 7885 34808 7971 34864
rect 8027 34808 8113 34864
rect 8169 34808 8255 34864
rect 8311 34808 8397 34864
rect 8453 34808 8539 34864
rect 8595 34808 8681 34864
rect 8737 34808 8823 34864
rect 8879 34808 8965 34864
rect 9021 34808 9107 34864
rect 9163 34808 9249 34864
rect 9305 34808 9391 34864
rect 9447 34808 9533 34864
rect 9589 34808 9675 34864
rect 9731 34808 9817 34864
rect 9873 34808 9959 34864
rect 10015 34808 10101 34864
rect 10157 34808 10243 34864
rect 10299 34808 10385 34864
rect 10441 34808 10527 34864
rect 10583 34808 10669 34864
rect 10725 34808 10811 34864
rect 10867 34808 10953 34864
rect 11009 34808 11095 34864
rect 11151 34808 11237 34864
rect 11293 34808 11379 34864
rect 11435 34808 11521 34864
rect 11577 34808 11663 34864
rect 11719 34808 11805 34864
rect 11861 34808 11947 34864
rect 12003 34808 12089 34864
rect 12145 34808 12231 34864
rect 12287 34808 12373 34864
rect 12429 34808 12515 34864
rect 12571 34808 12657 34864
rect 12713 34808 12799 34864
rect 12855 34808 12941 34864
rect 12997 34808 13083 34864
rect 13139 34808 13225 34864
rect 13281 34808 13367 34864
rect 13423 34808 13509 34864
rect 13565 34808 13651 34864
rect 13707 34808 13793 34864
rect 13849 34808 13935 34864
rect 13991 34808 14077 34864
rect 14133 34808 14219 34864
rect 14275 34808 14361 34864
rect 14417 34808 14503 34864
rect 14559 34808 14645 34864
rect 14701 34808 14787 34864
rect 14843 34808 15000 34864
rect 0 34722 15000 34808
rect 0 34666 161 34722
rect 217 34666 303 34722
rect 359 34666 445 34722
rect 501 34666 587 34722
rect 643 34666 729 34722
rect 785 34666 871 34722
rect 927 34666 1013 34722
rect 1069 34666 1155 34722
rect 1211 34666 1297 34722
rect 1353 34666 1439 34722
rect 1495 34666 1581 34722
rect 1637 34666 1723 34722
rect 1779 34666 1865 34722
rect 1921 34666 2007 34722
rect 2063 34666 2149 34722
rect 2205 34666 2291 34722
rect 2347 34666 2433 34722
rect 2489 34666 2575 34722
rect 2631 34666 2717 34722
rect 2773 34666 2859 34722
rect 2915 34666 3001 34722
rect 3057 34666 3143 34722
rect 3199 34666 3285 34722
rect 3341 34666 3427 34722
rect 3483 34666 3569 34722
rect 3625 34666 3711 34722
rect 3767 34666 3853 34722
rect 3909 34666 3995 34722
rect 4051 34666 4137 34722
rect 4193 34666 4279 34722
rect 4335 34666 4421 34722
rect 4477 34666 4563 34722
rect 4619 34666 4705 34722
rect 4761 34666 4847 34722
rect 4903 34666 4989 34722
rect 5045 34666 5131 34722
rect 5187 34666 5273 34722
rect 5329 34666 5415 34722
rect 5471 34666 5557 34722
rect 5613 34666 5699 34722
rect 5755 34666 5841 34722
rect 5897 34666 5983 34722
rect 6039 34666 6125 34722
rect 6181 34666 6267 34722
rect 6323 34666 6409 34722
rect 6465 34666 6551 34722
rect 6607 34666 6693 34722
rect 6749 34666 6835 34722
rect 6891 34666 6977 34722
rect 7033 34666 7119 34722
rect 7175 34666 7261 34722
rect 7317 34666 7403 34722
rect 7459 34666 7545 34722
rect 7601 34666 7687 34722
rect 7743 34666 7829 34722
rect 7885 34666 7971 34722
rect 8027 34666 8113 34722
rect 8169 34666 8255 34722
rect 8311 34666 8397 34722
rect 8453 34666 8539 34722
rect 8595 34666 8681 34722
rect 8737 34666 8823 34722
rect 8879 34666 8965 34722
rect 9021 34666 9107 34722
rect 9163 34666 9249 34722
rect 9305 34666 9391 34722
rect 9447 34666 9533 34722
rect 9589 34666 9675 34722
rect 9731 34666 9817 34722
rect 9873 34666 9959 34722
rect 10015 34666 10101 34722
rect 10157 34666 10243 34722
rect 10299 34666 10385 34722
rect 10441 34666 10527 34722
rect 10583 34666 10669 34722
rect 10725 34666 10811 34722
rect 10867 34666 10953 34722
rect 11009 34666 11095 34722
rect 11151 34666 11237 34722
rect 11293 34666 11379 34722
rect 11435 34666 11521 34722
rect 11577 34666 11663 34722
rect 11719 34666 11805 34722
rect 11861 34666 11947 34722
rect 12003 34666 12089 34722
rect 12145 34666 12231 34722
rect 12287 34666 12373 34722
rect 12429 34666 12515 34722
rect 12571 34666 12657 34722
rect 12713 34666 12799 34722
rect 12855 34666 12941 34722
rect 12997 34666 13083 34722
rect 13139 34666 13225 34722
rect 13281 34666 13367 34722
rect 13423 34666 13509 34722
rect 13565 34666 13651 34722
rect 13707 34666 13793 34722
rect 13849 34666 13935 34722
rect 13991 34666 14077 34722
rect 14133 34666 14219 34722
rect 14275 34666 14361 34722
rect 14417 34666 14503 34722
rect 14559 34666 14645 34722
rect 14701 34666 14787 34722
rect 14843 34666 15000 34722
rect 0 34580 15000 34666
rect 0 34524 161 34580
rect 217 34524 303 34580
rect 359 34524 445 34580
rect 501 34524 587 34580
rect 643 34524 729 34580
rect 785 34524 871 34580
rect 927 34524 1013 34580
rect 1069 34524 1155 34580
rect 1211 34524 1297 34580
rect 1353 34524 1439 34580
rect 1495 34524 1581 34580
rect 1637 34524 1723 34580
rect 1779 34524 1865 34580
rect 1921 34524 2007 34580
rect 2063 34524 2149 34580
rect 2205 34524 2291 34580
rect 2347 34524 2433 34580
rect 2489 34524 2575 34580
rect 2631 34524 2717 34580
rect 2773 34524 2859 34580
rect 2915 34524 3001 34580
rect 3057 34524 3143 34580
rect 3199 34524 3285 34580
rect 3341 34524 3427 34580
rect 3483 34524 3569 34580
rect 3625 34524 3711 34580
rect 3767 34524 3853 34580
rect 3909 34524 3995 34580
rect 4051 34524 4137 34580
rect 4193 34524 4279 34580
rect 4335 34524 4421 34580
rect 4477 34524 4563 34580
rect 4619 34524 4705 34580
rect 4761 34524 4847 34580
rect 4903 34524 4989 34580
rect 5045 34524 5131 34580
rect 5187 34524 5273 34580
rect 5329 34524 5415 34580
rect 5471 34524 5557 34580
rect 5613 34524 5699 34580
rect 5755 34524 5841 34580
rect 5897 34524 5983 34580
rect 6039 34524 6125 34580
rect 6181 34524 6267 34580
rect 6323 34524 6409 34580
rect 6465 34524 6551 34580
rect 6607 34524 6693 34580
rect 6749 34524 6835 34580
rect 6891 34524 6977 34580
rect 7033 34524 7119 34580
rect 7175 34524 7261 34580
rect 7317 34524 7403 34580
rect 7459 34524 7545 34580
rect 7601 34524 7687 34580
rect 7743 34524 7829 34580
rect 7885 34524 7971 34580
rect 8027 34524 8113 34580
rect 8169 34524 8255 34580
rect 8311 34524 8397 34580
rect 8453 34524 8539 34580
rect 8595 34524 8681 34580
rect 8737 34524 8823 34580
rect 8879 34524 8965 34580
rect 9021 34524 9107 34580
rect 9163 34524 9249 34580
rect 9305 34524 9391 34580
rect 9447 34524 9533 34580
rect 9589 34524 9675 34580
rect 9731 34524 9817 34580
rect 9873 34524 9959 34580
rect 10015 34524 10101 34580
rect 10157 34524 10243 34580
rect 10299 34524 10385 34580
rect 10441 34524 10527 34580
rect 10583 34524 10669 34580
rect 10725 34524 10811 34580
rect 10867 34524 10953 34580
rect 11009 34524 11095 34580
rect 11151 34524 11237 34580
rect 11293 34524 11379 34580
rect 11435 34524 11521 34580
rect 11577 34524 11663 34580
rect 11719 34524 11805 34580
rect 11861 34524 11947 34580
rect 12003 34524 12089 34580
rect 12145 34524 12231 34580
rect 12287 34524 12373 34580
rect 12429 34524 12515 34580
rect 12571 34524 12657 34580
rect 12713 34524 12799 34580
rect 12855 34524 12941 34580
rect 12997 34524 13083 34580
rect 13139 34524 13225 34580
rect 13281 34524 13367 34580
rect 13423 34524 13509 34580
rect 13565 34524 13651 34580
rect 13707 34524 13793 34580
rect 13849 34524 13935 34580
rect 13991 34524 14077 34580
rect 14133 34524 14219 34580
rect 14275 34524 14361 34580
rect 14417 34524 14503 34580
rect 14559 34524 14645 34580
rect 14701 34524 14787 34580
rect 14843 34524 15000 34580
rect 0 34438 15000 34524
rect 0 34382 161 34438
rect 217 34382 303 34438
rect 359 34382 445 34438
rect 501 34382 587 34438
rect 643 34382 729 34438
rect 785 34382 871 34438
rect 927 34382 1013 34438
rect 1069 34382 1155 34438
rect 1211 34382 1297 34438
rect 1353 34382 1439 34438
rect 1495 34382 1581 34438
rect 1637 34382 1723 34438
rect 1779 34382 1865 34438
rect 1921 34382 2007 34438
rect 2063 34382 2149 34438
rect 2205 34382 2291 34438
rect 2347 34382 2433 34438
rect 2489 34382 2575 34438
rect 2631 34382 2717 34438
rect 2773 34382 2859 34438
rect 2915 34382 3001 34438
rect 3057 34382 3143 34438
rect 3199 34382 3285 34438
rect 3341 34382 3427 34438
rect 3483 34382 3569 34438
rect 3625 34382 3711 34438
rect 3767 34382 3853 34438
rect 3909 34382 3995 34438
rect 4051 34382 4137 34438
rect 4193 34382 4279 34438
rect 4335 34382 4421 34438
rect 4477 34382 4563 34438
rect 4619 34382 4705 34438
rect 4761 34382 4847 34438
rect 4903 34382 4989 34438
rect 5045 34382 5131 34438
rect 5187 34382 5273 34438
rect 5329 34382 5415 34438
rect 5471 34382 5557 34438
rect 5613 34382 5699 34438
rect 5755 34382 5841 34438
rect 5897 34382 5983 34438
rect 6039 34382 6125 34438
rect 6181 34382 6267 34438
rect 6323 34382 6409 34438
rect 6465 34382 6551 34438
rect 6607 34382 6693 34438
rect 6749 34382 6835 34438
rect 6891 34382 6977 34438
rect 7033 34382 7119 34438
rect 7175 34382 7261 34438
rect 7317 34382 7403 34438
rect 7459 34382 7545 34438
rect 7601 34382 7687 34438
rect 7743 34382 7829 34438
rect 7885 34382 7971 34438
rect 8027 34382 8113 34438
rect 8169 34382 8255 34438
rect 8311 34382 8397 34438
rect 8453 34382 8539 34438
rect 8595 34382 8681 34438
rect 8737 34382 8823 34438
rect 8879 34382 8965 34438
rect 9021 34382 9107 34438
rect 9163 34382 9249 34438
rect 9305 34382 9391 34438
rect 9447 34382 9533 34438
rect 9589 34382 9675 34438
rect 9731 34382 9817 34438
rect 9873 34382 9959 34438
rect 10015 34382 10101 34438
rect 10157 34382 10243 34438
rect 10299 34382 10385 34438
rect 10441 34382 10527 34438
rect 10583 34382 10669 34438
rect 10725 34382 10811 34438
rect 10867 34382 10953 34438
rect 11009 34382 11095 34438
rect 11151 34382 11237 34438
rect 11293 34382 11379 34438
rect 11435 34382 11521 34438
rect 11577 34382 11663 34438
rect 11719 34382 11805 34438
rect 11861 34382 11947 34438
rect 12003 34382 12089 34438
rect 12145 34382 12231 34438
rect 12287 34382 12373 34438
rect 12429 34382 12515 34438
rect 12571 34382 12657 34438
rect 12713 34382 12799 34438
rect 12855 34382 12941 34438
rect 12997 34382 13083 34438
rect 13139 34382 13225 34438
rect 13281 34382 13367 34438
rect 13423 34382 13509 34438
rect 13565 34382 13651 34438
rect 13707 34382 13793 34438
rect 13849 34382 13935 34438
rect 13991 34382 14077 34438
rect 14133 34382 14219 34438
rect 14275 34382 14361 34438
rect 14417 34382 14503 34438
rect 14559 34382 14645 34438
rect 14701 34382 14787 34438
rect 14843 34382 15000 34438
rect 0 34296 15000 34382
rect 0 34240 161 34296
rect 217 34240 303 34296
rect 359 34240 445 34296
rect 501 34240 587 34296
rect 643 34240 729 34296
rect 785 34240 871 34296
rect 927 34240 1013 34296
rect 1069 34240 1155 34296
rect 1211 34240 1297 34296
rect 1353 34240 1439 34296
rect 1495 34240 1581 34296
rect 1637 34240 1723 34296
rect 1779 34240 1865 34296
rect 1921 34240 2007 34296
rect 2063 34240 2149 34296
rect 2205 34240 2291 34296
rect 2347 34240 2433 34296
rect 2489 34240 2575 34296
rect 2631 34240 2717 34296
rect 2773 34240 2859 34296
rect 2915 34240 3001 34296
rect 3057 34240 3143 34296
rect 3199 34240 3285 34296
rect 3341 34240 3427 34296
rect 3483 34240 3569 34296
rect 3625 34240 3711 34296
rect 3767 34240 3853 34296
rect 3909 34240 3995 34296
rect 4051 34240 4137 34296
rect 4193 34240 4279 34296
rect 4335 34240 4421 34296
rect 4477 34240 4563 34296
rect 4619 34240 4705 34296
rect 4761 34240 4847 34296
rect 4903 34240 4989 34296
rect 5045 34240 5131 34296
rect 5187 34240 5273 34296
rect 5329 34240 5415 34296
rect 5471 34240 5557 34296
rect 5613 34240 5699 34296
rect 5755 34240 5841 34296
rect 5897 34240 5983 34296
rect 6039 34240 6125 34296
rect 6181 34240 6267 34296
rect 6323 34240 6409 34296
rect 6465 34240 6551 34296
rect 6607 34240 6693 34296
rect 6749 34240 6835 34296
rect 6891 34240 6977 34296
rect 7033 34240 7119 34296
rect 7175 34240 7261 34296
rect 7317 34240 7403 34296
rect 7459 34240 7545 34296
rect 7601 34240 7687 34296
rect 7743 34240 7829 34296
rect 7885 34240 7971 34296
rect 8027 34240 8113 34296
rect 8169 34240 8255 34296
rect 8311 34240 8397 34296
rect 8453 34240 8539 34296
rect 8595 34240 8681 34296
rect 8737 34240 8823 34296
rect 8879 34240 8965 34296
rect 9021 34240 9107 34296
rect 9163 34240 9249 34296
rect 9305 34240 9391 34296
rect 9447 34240 9533 34296
rect 9589 34240 9675 34296
rect 9731 34240 9817 34296
rect 9873 34240 9959 34296
rect 10015 34240 10101 34296
rect 10157 34240 10243 34296
rect 10299 34240 10385 34296
rect 10441 34240 10527 34296
rect 10583 34240 10669 34296
rect 10725 34240 10811 34296
rect 10867 34240 10953 34296
rect 11009 34240 11095 34296
rect 11151 34240 11237 34296
rect 11293 34240 11379 34296
rect 11435 34240 11521 34296
rect 11577 34240 11663 34296
rect 11719 34240 11805 34296
rect 11861 34240 11947 34296
rect 12003 34240 12089 34296
rect 12145 34240 12231 34296
rect 12287 34240 12373 34296
rect 12429 34240 12515 34296
rect 12571 34240 12657 34296
rect 12713 34240 12799 34296
rect 12855 34240 12941 34296
rect 12997 34240 13083 34296
rect 13139 34240 13225 34296
rect 13281 34240 13367 34296
rect 13423 34240 13509 34296
rect 13565 34240 13651 34296
rect 13707 34240 13793 34296
rect 13849 34240 13935 34296
rect 13991 34240 14077 34296
rect 14133 34240 14219 34296
rect 14275 34240 14361 34296
rect 14417 34240 14503 34296
rect 14559 34240 14645 34296
rect 14701 34240 14787 34296
rect 14843 34240 15000 34296
rect 0 34154 15000 34240
rect 0 34098 161 34154
rect 217 34098 303 34154
rect 359 34098 445 34154
rect 501 34098 587 34154
rect 643 34098 729 34154
rect 785 34098 871 34154
rect 927 34098 1013 34154
rect 1069 34098 1155 34154
rect 1211 34098 1297 34154
rect 1353 34098 1439 34154
rect 1495 34098 1581 34154
rect 1637 34098 1723 34154
rect 1779 34098 1865 34154
rect 1921 34098 2007 34154
rect 2063 34098 2149 34154
rect 2205 34098 2291 34154
rect 2347 34098 2433 34154
rect 2489 34098 2575 34154
rect 2631 34098 2717 34154
rect 2773 34098 2859 34154
rect 2915 34098 3001 34154
rect 3057 34098 3143 34154
rect 3199 34098 3285 34154
rect 3341 34098 3427 34154
rect 3483 34098 3569 34154
rect 3625 34098 3711 34154
rect 3767 34098 3853 34154
rect 3909 34098 3995 34154
rect 4051 34098 4137 34154
rect 4193 34098 4279 34154
rect 4335 34098 4421 34154
rect 4477 34098 4563 34154
rect 4619 34098 4705 34154
rect 4761 34098 4847 34154
rect 4903 34098 4989 34154
rect 5045 34098 5131 34154
rect 5187 34098 5273 34154
rect 5329 34098 5415 34154
rect 5471 34098 5557 34154
rect 5613 34098 5699 34154
rect 5755 34098 5841 34154
rect 5897 34098 5983 34154
rect 6039 34098 6125 34154
rect 6181 34098 6267 34154
rect 6323 34098 6409 34154
rect 6465 34098 6551 34154
rect 6607 34098 6693 34154
rect 6749 34098 6835 34154
rect 6891 34098 6977 34154
rect 7033 34098 7119 34154
rect 7175 34098 7261 34154
rect 7317 34098 7403 34154
rect 7459 34098 7545 34154
rect 7601 34098 7687 34154
rect 7743 34098 7829 34154
rect 7885 34098 7971 34154
rect 8027 34098 8113 34154
rect 8169 34098 8255 34154
rect 8311 34098 8397 34154
rect 8453 34098 8539 34154
rect 8595 34098 8681 34154
rect 8737 34098 8823 34154
rect 8879 34098 8965 34154
rect 9021 34098 9107 34154
rect 9163 34098 9249 34154
rect 9305 34098 9391 34154
rect 9447 34098 9533 34154
rect 9589 34098 9675 34154
rect 9731 34098 9817 34154
rect 9873 34098 9959 34154
rect 10015 34098 10101 34154
rect 10157 34098 10243 34154
rect 10299 34098 10385 34154
rect 10441 34098 10527 34154
rect 10583 34098 10669 34154
rect 10725 34098 10811 34154
rect 10867 34098 10953 34154
rect 11009 34098 11095 34154
rect 11151 34098 11237 34154
rect 11293 34098 11379 34154
rect 11435 34098 11521 34154
rect 11577 34098 11663 34154
rect 11719 34098 11805 34154
rect 11861 34098 11947 34154
rect 12003 34098 12089 34154
rect 12145 34098 12231 34154
rect 12287 34098 12373 34154
rect 12429 34098 12515 34154
rect 12571 34098 12657 34154
rect 12713 34098 12799 34154
rect 12855 34098 12941 34154
rect 12997 34098 13083 34154
rect 13139 34098 13225 34154
rect 13281 34098 13367 34154
rect 13423 34098 13509 34154
rect 13565 34098 13651 34154
rect 13707 34098 13793 34154
rect 13849 34098 13935 34154
rect 13991 34098 14077 34154
rect 14133 34098 14219 34154
rect 14275 34098 14361 34154
rect 14417 34098 14503 34154
rect 14559 34098 14645 34154
rect 14701 34098 14787 34154
rect 14843 34098 15000 34154
rect 0 34012 15000 34098
rect 0 33956 161 34012
rect 217 33956 303 34012
rect 359 33956 445 34012
rect 501 33956 587 34012
rect 643 33956 729 34012
rect 785 33956 871 34012
rect 927 33956 1013 34012
rect 1069 33956 1155 34012
rect 1211 33956 1297 34012
rect 1353 33956 1439 34012
rect 1495 33956 1581 34012
rect 1637 33956 1723 34012
rect 1779 33956 1865 34012
rect 1921 33956 2007 34012
rect 2063 33956 2149 34012
rect 2205 33956 2291 34012
rect 2347 33956 2433 34012
rect 2489 33956 2575 34012
rect 2631 33956 2717 34012
rect 2773 33956 2859 34012
rect 2915 33956 3001 34012
rect 3057 33956 3143 34012
rect 3199 33956 3285 34012
rect 3341 33956 3427 34012
rect 3483 33956 3569 34012
rect 3625 33956 3711 34012
rect 3767 33956 3853 34012
rect 3909 33956 3995 34012
rect 4051 33956 4137 34012
rect 4193 33956 4279 34012
rect 4335 33956 4421 34012
rect 4477 33956 4563 34012
rect 4619 33956 4705 34012
rect 4761 33956 4847 34012
rect 4903 33956 4989 34012
rect 5045 33956 5131 34012
rect 5187 33956 5273 34012
rect 5329 33956 5415 34012
rect 5471 33956 5557 34012
rect 5613 33956 5699 34012
rect 5755 33956 5841 34012
rect 5897 33956 5983 34012
rect 6039 33956 6125 34012
rect 6181 33956 6267 34012
rect 6323 33956 6409 34012
rect 6465 33956 6551 34012
rect 6607 33956 6693 34012
rect 6749 33956 6835 34012
rect 6891 33956 6977 34012
rect 7033 33956 7119 34012
rect 7175 33956 7261 34012
rect 7317 33956 7403 34012
rect 7459 33956 7545 34012
rect 7601 33956 7687 34012
rect 7743 33956 7829 34012
rect 7885 33956 7971 34012
rect 8027 33956 8113 34012
rect 8169 33956 8255 34012
rect 8311 33956 8397 34012
rect 8453 33956 8539 34012
rect 8595 33956 8681 34012
rect 8737 33956 8823 34012
rect 8879 33956 8965 34012
rect 9021 33956 9107 34012
rect 9163 33956 9249 34012
rect 9305 33956 9391 34012
rect 9447 33956 9533 34012
rect 9589 33956 9675 34012
rect 9731 33956 9817 34012
rect 9873 33956 9959 34012
rect 10015 33956 10101 34012
rect 10157 33956 10243 34012
rect 10299 33956 10385 34012
rect 10441 33956 10527 34012
rect 10583 33956 10669 34012
rect 10725 33956 10811 34012
rect 10867 33956 10953 34012
rect 11009 33956 11095 34012
rect 11151 33956 11237 34012
rect 11293 33956 11379 34012
rect 11435 33956 11521 34012
rect 11577 33956 11663 34012
rect 11719 33956 11805 34012
rect 11861 33956 11947 34012
rect 12003 33956 12089 34012
rect 12145 33956 12231 34012
rect 12287 33956 12373 34012
rect 12429 33956 12515 34012
rect 12571 33956 12657 34012
rect 12713 33956 12799 34012
rect 12855 33956 12941 34012
rect 12997 33956 13083 34012
rect 13139 33956 13225 34012
rect 13281 33956 13367 34012
rect 13423 33956 13509 34012
rect 13565 33956 13651 34012
rect 13707 33956 13793 34012
rect 13849 33956 13935 34012
rect 13991 33956 14077 34012
rect 14133 33956 14219 34012
rect 14275 33956 14361 34012
rect 14417 33956 14503 34012
rect 14559 33956 14645 34012
rect 14701 33956 14787 34012
rect 14843 33956 15000 34012
rect 0 33870 15000 33956
rect 0 33814 161 33870
rect 217 33814 303 33870
rect 359 33814 445 33870
rect 501 33814 587 33870
rect 643 33814 729 33870
rect 785 33814 871 33870
rect 927 33814 1013 33870
rect 1069 33814 1155 33870
rect 1211 33814 1297 33870
rect 1353 33814 1439 33870
rect 1495 33814 1581 33870
rect 1637 33814 1723 33870
rect 1779 33814 1865 33870
rect 1921 33814 2007 33870
rect 2063 33814 2149 33870
rect 2205 33814 2291 33870
rect 2347 33814 2433 33870
rect 2489 33814 2575 33870
rect 2631 33814 2717 33870
rect 2773 33814 2859 33870
rect 2915 33814 3001 33870
rect 3057 33814 3143 33870
rect 3199 33814 3285 33870
rect 3341 33814 3427 33870
rect 3483 33814 3569 33870
rect 3625 33814 3711 33870
rect 3767 33814 3853 33870
rect 3909 33814 3995 33870
rect 4051 33814 4137 33870
rect 4193 33814 4279 33870
rect 4335 33814 4421 33870
rect 4477 33814 4563 33870
rect 4619 33814 4705 33870
rect 4761 33814 4847 33870
rect 4903 33814 4989 33870
rect 5045 33814 5131 33870
rect 5187 33814 5273 33870
rect 5329 33814 5415 33870
rect 5471 33814 5557 33870
rect 5613 33814 5699 33870
rect 5755 33814 5841 33870
rect 5897 33814 5983 33870
rect 6039 33814 6125 33870
rect 6181 33814 6267 33870
rect 6323 33814 6409 33870
rect 6465 33814 6551 33870
rect 6607 33814 6693 33870
rect 6749 33814 6835 33870
rect 6891 33814 6977 33870
rect 7033 33814 7119 33870
rect 7175 33814 7261 33870
rect 7317 33814 7403 33870
rect 7459 33814 7545 33870
rect 7601 33814 7687 33870
rect 7743 33814 7829 33870
rect 7885 33814 7971 33870
rect 8027 33814 8113 33870
rect 8169 33814 8255 33870
rect 8311 33814 8397 33870
rect 8453 33814 8539 33870
rect 8595 33814 8681 33870
rect 8737 33814 8823 33870
rect 8879 33814 8965 33870
rect 9021 33814 9107 33870
rect 9163 33814 9249 33870
rect 9305 33814 9391 33870
rect 9447 33814 9533 33870
rect 9589 33814 9675 33870
rect 9731 33814 9817 33870
rect 9873 33814 9959 33870
rect 10015 33814 10101 33870
rect 10157 33814 10243 33870
rect 10299 33814 10385 33870
rect 10441 33814 10527 33870
rect 10583 33814 10669 33870
rect 10725 33814 10811 33870
rect 10867 33814 10953 33870
rect 11009 33814 11095 33870
rect 11151 33814 11237 33870
rect 11293 33814 11379 33870
rect 11435 33814 11521 33870
rect 11577 33814 11663 33870
rect 11719 33814 11805 33870
rect 11861 33814 11947 33870
rect 12003 33814 12089 33870
rect 12145 33814 12231 33870
rect 12287 33814 12373 33870
rect 12429 33814 12515 33870
rect 12571 33814 12657 33870
rect 12713 33814 12799 33870
rect 12855 33814 12941 33870
rect 12997 33814 13083 33870
rect 13139 33814 13225 33870
rect 13281 33814 13367 33870
rect 13423 33814 13509 33870
rect 13565 33814 13651 33870
rect 13707 33814 13793 33870
rect 13849 33814 13935 33870
rect 13991 33814 14077 33870
rect 14133 33814 14219 33870
rect 14275 33814 14361 33870
rect 14417 33814 14503 33870
rect 14559 33814 14645 33870
rect 14701 33814 14787 33870
rect 14843 33814 15000 33870
rect 0 33728 15000 33814
rect 0 33672 161 33728
rect 217 33672 303 33728
rect 359 33672 445 33728
rect 501 33672 587 33728
rect 643 33672 729 33728
rect 785 33672 871 33728
rect 927 33672 1013 33728
rect 1069 33672 1155 33728
rect 1211 33672 1297 33728
rect 1353 33672 1439 33728
rect 1495 33672 1581 33728
rect 1637 33672 1723 33728
rect 1779 33672 1865 33728
rect 1921 33672 2007 33728
rect 2063 33672 2149 33728
rect 2205 33672 2291 33728
rect 2347 33672 2433 33728
rect 2489 33672 2575 33728
rect 2631 33672 2717 33728
rect 2773 33672 2859 33728
rect 2915 33672 3001 33728
rect 3057 33672 3143 33728
rect 3199 33672 3285 33728
rect 3341 33672 3427 33728
rect 3483 33672 3569 33728
rect 3625 33672 3711 33728
rect 3767 33672 3853 33728
rect 3909 33672 3995 33728
rect 4051 33672 4137 33728
rect 4193 33672 4279 33728
rect 4335 33672 4421 33728
rect 4477 33672 4563 33728
rect 4619 33672 4705 33728
rect 4761 33672 4847 33728
rect 4903 33672 4989 33728
rect 5045 33672 5131 33728
rect 5187 33672 5273 33728
rect 5329 33672 5415 33728
rect 5471 33672 5557 33728
rect 5613 33672 5699 33728
rect 5755 33672 5841 33728
rect 5897 33672 5983 33728
rect 6039 33672 6125 33728
rect 6181 33672 6267 33728
rect 6323 33672 6409 33728
rect 6465 33672 6551 33728
rect 6607 33672 6693 33728
rect 6749 33672 6835 33728
rect 6891 33672 6977 33728
rect 7033 33672 7119 33728
rect 7175 33672 7261 33728
rect 7317 33672 7403 33728
rect 7459 33672 7545 33728
rect 7601 33672 7687 33728
rect 7743 33672 7829 33728
rect 7885 33672 7971 33728
rect 8027 33672 8113 33728
rect 8169 33672 8255 33728
rect 8311 33672 8397 33728
rect 8453 33672 8539 33728
rect 8595 33672 8681 33728
rect 8737 33672 8823 33728
rect 8879 33672 8965 33728
rect 9021 33672 9107 33728
rect 9163 33672 9249 33728
rect 9305 33672 9391 33728
rect 9447 33672 9533 33728
rect 9589 33672 9675 33728
rect 9731 33672 9817 33728
rect 9873 33672 9959 33728
rect 10015 33672 10101 33728
rect 10157 33672 10243 33728
rect 10299 33672 10385 33728
rect 10441 33672 10527 33728
rect 10583 33672 10669 33728
rect 10725 33672 10811 33728
rect 10867 33672 10953 33728
rect 11009 33672 11095 33728
rect 11151 33672 11237 33728
rect 11293 33672 11379 33728
rect 11435 33672 11521 33728
rect 11577 33672 11663 33728
rect 11719 33672 11805 33728
rect 11861 33672 11947 33728
rect 12003 33672 12089 33728
rect 12145 33672 12231 33728
rect 12287 33672 12373 33728
rect 12429 33672 12515 33728
rect 12571 33672 12657 33728
rect 12713 33672 12799 33728
rect 12855 33672 12941 33728
rect 12997 33672 13083 33728
rect 13139 33672 13225 33728
rect 13281 33672 13367 33728
rect 13423 33672 13509 33728
rect 13565 33672 13651 33728
rect 13707 33672 13793 33728
rect 13849 33672 13935 33728
rect 13991 33672 14077 33728
rect 14133 33672 14219 33728
rect 14275 33672 14361 33728
rect 14417 33672 14503 33728
rect 14559 33672 14645 33728
rect 14701 33672 14787 33728
rect 14843 33672 15000 33728
rect 0 33586 15000 33672
rect 0 33530 161 33586
rect 217 33530 303 33586
rect 359 33530 445 33586
rect 501 33530 587 33586
rect 643 33530 729 33586
rect 785 33530 871 33586
rect 927 33530 1013 33586
rect 1069 33530 1155 33586
rect 1211 33530 1297 33586
rect 1353 33530 1439 33586
rect 1495 33530 1581 33586
rect 1637 33530 1723 33586
rect 1779 33530 1865 33586
rect 1921 33530 2007 33586
rect 2063 33530 2149 33586
rect 2205 33530 2291 33586
rect 2347 33530 2433 33586
rect 2489 33530 2575 33586
rect 2631 33530 2717 33586
rect 2773 33530 2859 33586
rect 2915 33530 3001 33586
rect 3057 33530 3143 33586
rect 3199 33530 3285 33586
rect 3341 33530 3427 33586
rect 3483 33530 3569 33586
rect 3625 33530 3711 33586
rect 3767 33530 3853 33586
rect 3909 33530 3995 33586
rect 4051 33530 4137 33586
rect 4193 33530 4279 33586
rect 4335 33530 4421 33586
rect 4477 33530 4563 33586
rect 4619 33530 4705 33586
rect 4761 33530 4847 33586
rect 4903 33530 4989 33586
rect 5045 33530 5131 33586
rect 5187 33530 5273 33586
rect 5329 33530 5415 33586
rect 5471 33530 5557 33586
rect 5613 33530 5699 33586
rect 5755 33530 5841 33586
rect 5897 33530 5983 33586
rect 6039 33530 6125 33586
rect 6181 33530 6267 33586
rect 6323 33530 6409 33586
rect 6465 33530 6551 33586
rect 6607 33530 6693 33586
rect 6749 33530 6835 33586
rect 6891 33530 6977 33586
rect 7033 33530 7119 33586
rect 7175 33530 7261 33586
rect 7317 33530 7403 33586
rect 7459 33530 7545 33586
rect 7601 33530 7687 33586
rect 7743 33530 7829 33586
rect 7885 33530 7971 33586
rect 8027 33530 8113 33586
rect 8169 33530 8255 33586
rect 8311 33530 8397 33586
rect 8453 33530 8539 33586
rect 8595 33530 8681 33586
rect 8737 33530 8823 33586
rect 8879 33530 8965 33586
rect 9021 33530 9107 33586
rect 9163 33530 9249 33586
rect 9305 33530 9391 33586
rect 9447 33530 9533 33586
rect 9589 33530 9675 33586
rect 9731 33530 9817 33586
rect 9873 33530 9959 33586
rect 10015 33530 10101 33586
rect 10157 33530 10243 33586
rect 10299 33530 10385 33586
rect 10441 33530 10527 33586
rect 10583 33530 10669 33586
rect 10725 33530 10811 33586
rect 10867 33530 10953 33586
rect 11009 33530 11095 33586
rect 11151 33530 11237 33586
rect 11293 33530 11379 33586
rect 11435 33530 11521 33586
rect 11577 33530 11663 33586
rect 11719 33530 11805 33586
rect 11861 33530 11947 33586
rect 12003 33530 12089 33586
rect 12145 33530 12231 33586
rect 12287 33530 12373 33586
rect 12429 33530 12515 33586
rect 12571 33530 12657 33586
rect 12713 33530 12799 33586
rect 12855 33530 12941 33586
rect 12997 33530 13083 33586
rect 13139 33530 13225 33586
rect 13281 33530 13367 33586
rect 13423 33530 13509 33586
rect 13565 33530 13651 33586
rect 13707 33530 13793 33586
rect 13849 33530 13935 33586
rect 13991 33530 14077 33586
rect 14133 33530 14219 33586
rect 14275 33530 14361 33586
rect 14417 33530 14503 33586
rect 14559 33530 14645 33586
rect 14701 33530 14787 33586
rect 14843 33530 15000 33586
rect 0 33444 15000 33530
rect 0 33388 161 33444
rect 217 33388 303 33444
rect 359 33388 445 33444
rect 501 33388 587 33444
rect 643 33388 729 33444
rect 785 33388 871 33444
rect 927 33388 1013 33444
rect 1069 33388 1155 33444
rect 1211 33388 1297 33444
rect 1353 33388 1439 33444
rect 1495 33388 1581 33444
rect 1637 33388 1723 33444
rect 1779 33388 1865 33444
rect 1921 33388 2007 33444
rect 2063 33388 2149 33444
rect 2205 33388 2291 33444
rect 2347 33388 2433 33444
rect 2489 33388 2575 33444
rect 2631 33388 2717 33444
rect 2773 33388 2859 33444
rect 2915 33388 3001 33444
rect 3057 33388 3143 33444
rect 3199 33388 3285 33444
rect 3341 33388 3427 33444
rect 3483 33388 3569 33444
rect 3625 33388 3711 33444
rect 3767 33388 3853 33444
rect 3909 33388 3995 33444
rect 4051 33388 4137 33444
rect 4193 33388 4279 33444
rect 4335 33388 4421 33444
rect 4477 33388 4563 33444
rect 4619 33388 4705 33444
rect 4761 33388 4847 33444
rect 4903 33388 4989 33444
rect 5045 33388 5131 33444
rect 5187 33388 5273 33444
rect 5329 33388 5415 33444
rect 5471 33388 5557 33444
rect 5613 33388 5699 33444
rect 5755 33388 5841 33444
rect 5897 33388 5983 33444
rect 6039 33388 6125 33444
rect 6181 33388 6267 33444
rect 6323 33388 6409 33444
rect 6465 33388 6551 33444
rect 6607 33388 6693 33444
rect 6749 33388 6835 33444
rect 6891 33388 6977 33444
rect 7033 33388 7119 33444
rect 7175 33388 7261 33444
rect 7317 33388 7403 33444
rect 7459 33388 7545 33444
rect 7601 33388 7687 33444
rect 7743 33388 7829 33444
rect 7885 33388 7971 33444
rect 8027 33388 8113 33444
rect 8169 33388 8255 33444
rect 8311 33388 8397 33444
rect 8453 33388 8539 33444
rect 8595 33388 8681 33444
rect 8737 33388 8823 33444
rect 8879 33388 8965 33444
rect 9021 33388 9107 33444
rect 9163 33388 9249 33444
rect 9305 33388 9391 33444
rect 9447 33388 9533 33444
rect 9589 33388 9675 33444
rect 9731 33388 9817 33444
rect 9873 33388 9959 33444
rect 10015 33388 10101 33444
rect 10157 33388 10243 33444
rect 10299 33388 10385 33444
rect 10441 33388 10527 33444
rect 10583 33388 10669 33444
rect 10725 33388 10811 33444
rect 10867 33388 10953 33444
rect 11009 33388 11095 33444
rect 11151 33388 11237 33444
rect 11293 33388 11379 33444
rect 11435 33388 11521 33444
rect 11577 33388 11663 33444
rect 11719 33388 11805 33444
rect 11861 33388 11947 33444
rect 12003 33388 12089 33444
rect 12145 33388 12231 33444
rect 12287 33388 12373 33444
rect 12429 33388 12515 33444
rect 12571 33388 12657 33444
rect 12713 33388 12799 33444
rect 12855 33388 12941 33444
rect 12997 33388 13083 33444
rect 13139 33388 13225 33444
rect 13281 33388 13367 33444
rect 13423 33388 13509 33444
rect 13565 33388 13651 33444
rect 13707 33388 13793 33444
rect 13849 33388 13935 33444
rect 13991 33388 14077 33444
rect 14133 33388 14219 33444
rect 14275 33388 14361 33444
rect 14417 33388 14503 33444
rect 14559 33388 14645 33444
rect 14701 33388 14787 33444
rect 14843 33388 15000 33444
rect 0 33302 15000 33388
rect 0 33246 161 33302
rect 217 33246 303 33302
rect 359 33246 445 33302
rect 501 33246 587 33302
rect 643 33246 729 33302
rect 785 33246 871 33302
rect 927 33246 1013 33302
rect 1069 33246 1155 33302
rect 1211 33246 1297 33302
rect 1353 33246 1439 33302
rect 1495 33246 1581 33302
rect 1637 33246 1723 33302
rect 1779 33246 1865 33302
rect 1921 33246 2007 33302
rect 2063 33246 2149 33302
rect 2205 33246 2291 33302
rect 2347 33246 2433 33302
rect 2489 33246 2575 33302
rect 2631 33246 2717 33302
rect 2773 33246 2859 33302
rect 2915 33246 3001 33302
rect 3057 33246 3143 33302
rect 3199 33246 3285 33302
rect 3341 33246 3427 33302
rect 3483 33246 3569 33302
rect 3625 33246 3711 33302
rect 3767 33246 3853 33302
rect 3909 33246 3995 33302
rect 4051 33246 4137 33302
rect 4193 33246 4279 33302
rect 4335 33246 4421 33302
rect 4477 33246 4563 33302
rect 4619 33246 4705 33302
rect 4761 33246 4847 33302
rect 4903 33246 4989 33302
rect 5045 33246 5131 33302
rect 5187 33246 5273 33302
rect 5329 33246 5415 33302
rect 5471 33246 5557 33302
rect 5613 33246 5699 33302
rect 5755 33246 5841 33302
rect 5897 33246 5983 33302
rect 6039 33246 6125 33302
rect 6181 33246 6267 33302
rect 6323 33246 6409 33302
rect 6465 33246 6551 33302
rect 6607 33246 6693 33302
rect 6749 33246 6835 33302
rect 6891 33246 6977 33302
rect 7033 33246 7119 33302
rect 7175 33246 7261 33302
rect 7317 33246 7403 33302
rect 7459 33246 7545 33302
rect 7601 33246 7687 33302
rect 7743 33246 7829 33302
rect 7885 33246 7971 33302
rect 8027 33246 8113 33302
rect 8169 33246 8255 33302
rect 8311 33246 8397 33302
rect 8453 33246 8539 33302
rect 8595 33246 8681 33302
rect 8737 33246 8823 33302
rect 8879 33246 8965 33302
rect 9021 33246 9107 33302
rect 9163 33246 9249 33302
rect 9305 33246 9391 33302
rect 9447 33246 9533 33302
rect 9589 33246 9675 33302
rect 9731 33246 9817 33302
rect 9873 33246 9959 33302
rect 10015 33246 10101 33302
rect 10157 33246 10243 33302
rect 10299 33246 10385 33302
rect 10441 33246 10527 33302
rect 10583 33246 10669 33302
rect 10725 33246 10811 33302
rect 10867 33246 10953 33302
rect 11009 33246 11095 33302
rect 11151 33246 11237 33302
rect 11293 33246 11379 33302
rect 11435 33246 11521 33302
rect 11577 33246 11663 33302
rect 11719 33246 11805 33302
rect 11861 33246 11947 33302
rect 12003 33246 12089 33302
rect 12145 33246 12231 33302
rect 12287 33246 12373 33302
rect 12429 33246 12515 33302
rect 12571 33246 12657 33302
rect 12713 33246 12799 33302
rect 12855 33246 12941 33302
rect 12997 33246 13083 33302
rect 13139 33246 13225 33302
rect 13281 33246 13367 33302
rect 13423 33246 13509 33302
rect 13565 33246 13651 33302
rect 13707 33246 13793 33302
rect 13849 33246 13935 33302
rect 13991 33246 14077 33302
rect 14133 33246 14219 33302
rect 14275 33246 14361 33302
rect 14417 33246 14503 33302
rect 14559 33246 14645 33302
rect 14701 33246 14787 33302
rect 14843 33246 15000 33302
rect 0 33200 15000 33246
rect 937 33000 3937 33200
rect 4337 33000 7337 33200
rect 7737 33000 10737 33200
rect 11137 33000 14137 33200
rect 0 32941 15000 33000
rect 0 32885 161 32941
rect 217 32885 303 32941
rect 359 32885 445 32941
rect 501 32885 587 32941
rect 643 32885 729 32941
rect 785 32885 871 32941
rect 927 32885 1013 32941
rect 1069 32885 1155 32941
rect 1211 32885 1297 32941
rect 1353 32885 1439 32941
rect 1495 32885 1581 32941
rect 1637 32885 1723 32941
rect 1779 32885 1865 32941
rect 1921 32885 2007 32941
rect 2063 32885 2149 32941
rect 2205 32885 2291 32941
rect 2347 32885 2433 32941
rect 2489 32885 2575 32941
rect 2631 32885 2717 32941
rect 2773 32885 2859 32941
rect 2915 32885 3001 32941
rect 3057 32885 3143 32941
rect 3199 32885 3285 32941
rect 3341 32885 3427 32941
rect 3483 32885 3569 32941
rect 3625 32885 3711 32941
rect 3767 32885 3853 32941
rect 3909 32885 3995 32941
rect 4051 32885 4137 32941
rect 4193 32885 4279 32941
rect 4335 32885 4421 32941
rect 4477 32885 4563 32941
rect 4619 32885 4705 32941
rect 4761 32885 4847 32941
rect 4903 32885 4989 32941
rect 5045 32885 5131 32941
rect 5187 32885 5273 32941
rect 5329 32885 5415 32941
rect 5471 32885 5557 32941
rect 5613 32885 5699 32941
rect 5755 32885 5841 32941
rect 5897 32885 5983 32941
rect 6039 32885 6125 32941
rect 6181 32885 6267 32941
rect 6323 32885 6409 32941
rect 6465 32885 6551 32941
rect 6607 32885 6693 32941
rect 6749 32885 6835 32941
rect 6891 32885 6977 32941
rect 7033 32885 7119 32941
rect 7175 32885 7261 32941
rect 7317 32885 7403 32941
rect 7459 32885 7545 32941
rect 7601 32885 7687 32941
rect 7743 32885 7829 32941
rect 7885 32885 7971 32941
rect 8027 32885 8113 32941
rect 8169 32885 8255 32941
rect 8311 32885 8397 32941
rect 8453 32885 8539 32941
rect 8595 32885 8681 32941
rect 8737 32885 8823 32941
rect 8879 32885 8965 32941
rect 9021 32885 9107 32941
rect 9163 32885 9249 32941
rect 9305 32885 9391 32941
rect 9447 32885 9533 32941
rect 9589 32885 9675 32941
rect 9731 32885 9817 32941
rect 9873 32885 9959 32941
rect 10015 32885 10101 32941
rect 10157 32885 10243 32941
rect 10299 32885 10385 32941
rect 10441 32885 10527 32941
rect 10583 32885 10669 32941
rect 10725 32885 10811 32941
rect 10867 32885 10953 32941
rect 11009 32885 11095 32941
rect 11151 32885 11237 32941
rect 11293 32885 11379 32941
rect 11435 32885 11521 32941
rect 11577 32885 11663 32941
rect 11719 32885 11805 32941
rect 11861 32885 11947 32941
rect 12003 32885 12089 32941
rect 12145 32885 12231 32941
rect 12287 32885 12373 32941
rect 12429 32885 12515 32941
rect 12571 32885 12657 32941
rect 12713 32885 12799 32941
rect 12855 32885 12941 32941
rect 12997 32885 13083 32941
rect 13139 32885 13225 32941
rect 13281 32885 13367 32941
rect 13423 32885 13509 32941
rect 13565 32885 13651 32941
rect 13707 32885 13793 32941
rect 13849 32885 13935 32941
rect 13991 32885 14077 32941
rect 14133 32885 14219 32941
rect 14275 32885 14361 32941
rect 14417 32885 14503 32941
rect 14559 32885 14645 32941
rect 14701 32885 14787 32941
rect 14843 32885 15000 32941
rect 0 32799 15000 32885
rect 0 32743 161 32799
rect 217 32743 303 32799
rect 359 32743 445 32799
rect 501 32743 587 32799
rect 643 32743 729 32799
rect 785 32743 871 32799
rect 927 32743 1013 32799
rect 1069 32743 1155 32799
rect 1211 32743 1297 32799
rect 1353 32743 1439 32799
rect 1495 32743 1581 32799
rect 1637 32743 1723 32799
rect 1779 32743 1865 32799
rect 1921 32743 2007 32799
rect 2063 32743 2149 32799
rect 2205 32743 2291 32799
rect 2347 32743 2433 32799
rect 2489 32743 2575 32799
rect 2631 32743 2717 32799
rect 2773 32743 2859 32799
rect 2915 32743 3001 32799
rect 3057 32743 3143 32799
rect 3199 32743 3285 32799
rect 3341 32743 3427 32799
rect 3483 32743 3569 32799
rect 3625 32743 3711 32799
rect 3767 32743 3853 32799
rect 3909 32743 3995 32799
rect 4051 32743 4137 32799
rect 4193 32743 4279 32799
rect 4335 32743 4421 32799
rect 4477 32743 4563 32799
rect 4619 32743 4705 32799
rect 4761 32743 4847 32799
rect 4903 32743 4989 32799
rect 5045 32743 5131 32799
rect 5187 32743 5273 32799
rect 5329 32743 5415 32799
rect 5471 32743 5557 32799
rect 5613 32743 5699 32799
rect 5755 32743 5841 32799
rect 5897 32743 5983 32799
rect 6039 32743 6125 32799
rect 6181 32743 6267 32799
rect 6323 32743 6409 32799
rect 6465 32743 6551 32799
rect 6607 32743 6693 32799
rect 6749 32743 6835 32799
rect 6891 32743 6977 32799
rect 7033 32743 7119 32799
rect 7175 32743 7261 32799
rect 7317 32743 7403 32799
rect 7459 32743 7545 32799
rect 7601 32743 7687 32799
rect 7743 32743 7829 32799
rect 7885 32743 7971 32799
rect 8027 32743 8113 32799
rect 8169 32743 8255 32799
rect 8311 32743 8397 32799
rect 8453 32743 8539 32799
rect 8595 32743 8681 32799
rect 8737 32743 8823 32799
rect 8879 32743 8965 32799
rect 9021 32743 9107 32799
rect 9163 32743 9249 32799
rect 9305 32743 9391 32799
rect 9447 32743 9533 32799
rect 9589 32743 9675 32799
rect 9731 32743 9817 32799
rect 9873 32743 9959 32799
rect 10015 32743 10101 32799
rect 10157 32743 10243 32799
rect 10299 32743 10385 32799
rect 10441 32743 10527 32799
rect 10583 32743 10669 32799
rect 10725 32743 10811 32799
rect 10867 32743 10953 32799
rect 11009 32743 11095 32799
rect 11151 32743 11237 32799
rect 11293 32743 11379 32799
rect 11435 32743 11521 32799
rect 11577 32743 11663 32799
rect 11719 32743 11805 32799
rect 11861 32743 11947 32799
rect 12003 32743 12089 32799
rect 12145 32743 12231 32799
rect 12287 32743 12373 32799
rect 12429 32743 12515 32799
rect 12571 32743 12657 32799
rect 12713 32743 12799 32799
rect 12855 32743 12941 32799
rect 12997 32743 13083 32799
rect 13139 32743 13225 32799
rect 13281 32743 13367 32799
rect 13423 32743 13509 32799
rect 13565 32743 13651 32799
rect 13707 32743 13793 32799
rect 13849 32743 13935 32799
rect 13991 32743 14077 32799
rect 14133 32743 14219 32799
rect 14275 32743 14361 32799
rect 14417 32743 14503 32799
rect 14559 32743 14645 32799
rect 14701 32743 14787 32799
rect 14843 32743 15000 32799
rect 0 32657 15000 32743
rect 0 32601 161 32657
rect 217 32601 303 32657
rect 359 32601 445 32657
rect 501 32601 587 32657
rect 643 32601 729 32657
rect 785 32601 871 32657
rect 927 32601 1013 32657
rect 1069 32601 1155 32657
rect 1211 32601 1297 32657
rect 1353 32601 1439 32657
rect 1495 32601 1581 32657
rect 1637 32601 1723 32657
rect 1779 32601 1865 32657
rect 1921 32601 2007 32657
rect 2063 32601 2149 32657
rect 2205 32601 2291 32657
rect 2347 32601 2433 32657
rect 2489 32601 2575 32657
rect 2631 32601 2717 32657
rect 2773 32601 2859 32657
rect 2915 32601 3001 32657
rect 3057 32601 3143 32657
rect 3199 32601 3285 32657
rect 3341 32601 3427 32657
rect 3483 32601 3569 32657
rect 3625 32601 3711 32657
rect 3767 32601 3853 32657
rect 3909 32601 3995 32657
rect 4051 32601 4137 32657
rect 4193 32601 4279 32657
rect 4335 32601 4421 32657
rect 4477 32601 4563 32657
rect 4619 32601 4705 32657
rect 4761 32601 4847 32657
rect 4903 32601 4989 32657
rect 5045 32601 5131 32657
rect 5187 32601 5273 32657
rect 5329 32601 5415 32657
rect 5471 32601 5557 32657
rect 5613 32601 5699 32657
rect 5755 32601 5841 32657
rect 5897 32601 5983 32657
rect 6039 32601 6125 32657
rect 6181 32601 6267 32657
rect 6323 32601 6409 32657
rect 6465 32601 6551 32657
rect 6607 32601 6693 32657
rect 6749 32601 6835 32657
rect 6891 32601 6977 32657
rect 7033 32601 7119 32657
rect 7175 32601 7261 32657
rect 7317 32601 7403 32657
rect 7459 32601 7545 32657
rect 7601 32601 7687 32657
rect 7743 32601 7829 32657
rect 7885 32601 7971 32657
rect 8027 32601 8113 32657
rect 8169 32601 8255 32657
rect 8311 32601 8397 32657
rect 8453 32601 8539 32657
rect 8595 32601 8681 32657
rect 8737 32601 8823 32657
rect 8879 32601 8965 32657
rect 9021 32601 9107 32657
rect 9163 32601 9249 32657
rect 9305 32601 9391 32657
rect 9447 32601 9533 32657
rect 9589 32601 9675 32657
rect 9731 32601 9817 32657
rect 9873 32601 9959 32657
rect 10015 32601 10101 32657
rect 10157 32601 10243 32657
rect 10299 32601 10385 32657
rect 10441 32601 10527 32657
rect 10583 32601 10669 32657
rect 10725 32601 10811 32657
rect 10867 32601 10953 32657
rect 11009 32601 11095 32657
rect 11151 32601 11237 32657
rect 11293 32601 11379 32657
rect 11435 32601 11521 32657
rect 11577 32601 11663 32657
rect 11719 32601 11805 32657
rect 11861 32601 11947 32657
rect 12003 32601 12089 32657
rect 12145 32601 12231 32657
rect 12287 32601 12373 32657
rect 12429 32601 12515 32657
rect 12571 32601 12657 32657
rect 12713 32601 12799 32657
rect 12855 32601 12941 32657
rect 12997 32601 13083 32657
rect 13139 32601 13225 32657
rect 13281 32601 13367 32657
rect 13423 32601 13509 32657
rect 13565 32601 13651 32657
rect 13707 32601 13793 32657
rect 13849 32601 13935 32657
rect 13991 32601 14077 32657
rect 14133 32601 14219 32657
rect 14275 32601 14361 32657
rect 14417 32601 14503 32657
rect 14559 32601 14645 32657
rect 14701 32601 14787 32657
rect 14843 32601 15000 32657
rect 0 32515 15000 32601
rect 0 32459 161 32515
rect 217 32459 303 32515
rect 359 32459 445 32515
rect 501 32459 587 32515
rect 643 32459 729 32515
rect 785 32459 871 32515
rect 927 32459 1013 32515
rect 1069 32459 1155 32515
rect 1211 32459 1297 32515
rect 1353 32459 1439 32515
rect 1495 32459 1581 32515
rect 1637 32459 1723 32515
rect 1779 32459 1865 32515
rect 1921 32459 2007 32515
rect 2063 32459 2149 32515
rect 2205 32459 2291 32515
rect 2347 32459 2433 32515
rect 2489 32459 2575 32515
rect 2631 32459 2717 32515
rect 2773 32459 2859 32515
rect 2915 32459 3001 32515
rect 3057 32459 3143 32515
rect 3199 32459 3285 32515
rect 3341 32459 3427 32515
rect 3483 32459 3569 32515
rect 3625 32459 3711 32515
rect 3767 32459 3853 32515
rect 3909 32459 3995 32515
rect 4051 32459 4137 32515
rect 4193 32459 4279 32515
rect 4335 32459 4421 32515
rect 4477 32459 4563 32515
rect 4619 32459 4705 32515
rect 4761 32459 4847 32515
rect 4903 32459 4989 32515
rect 5045 32459 5131 32515
rect 5187 32459 5273 32515
rect 5329 32459 5415 32515
rect 5471 32459 5557 32515
rect 5613 32459 5699 32515
rect 5755 32459 5841 32515
rect 5897 32459 5983 32515
rect 6039 32459 6125 32515
rect 6181 32459 6267 32515
rect 6323 32459 6409 32515
rect 6465 32459 6551 32515
rect 6607 32459 6693 32515
rect 6749 32459 6835 32515
rect 6891 32459 6977 32515
rect 7033 32459 7119 32515
rect 7175 32459 7261 32515
rect 7317 32459 7403 32515
rect 7459 32459 7545 32515
rect 7601 32459 7687 32515
rect 7743 32459 7829 32515
rect 7885 32459 7971 32515
rect 8027 32459 8113 32515
rect 8169 32459 8255 32515
rect 8311 32459 8397 32515
rect 8453 32459 8539 32515
rect 8595 32459 8681 32515
rect 8737 32459 8823 32515
rect 8879 32459 8965 32515
rect 9021 32459 9107 32515
rect 9163 32459 9249 32515
rect 9305 32459 9391 32515
rect 9447 32459 9533 32515
rect 9589 32459 9675 32515
rect 9731 32459 9817 32515
rect 9873 32459 9959 32515
rect 10015 32459 10101 32515
rect 10157 32459 10243 32515
rect 10299 32459 10385 32515
rect 10441 32459 10527 32515
rect 10583 32459 10669 32515
rect 10725 32459 10811 32515
rect 10867 32459 10953 32515
rect 11009 32459 11095 32515
rect 11151 32459 11237 32515
rect 11293 32459 11379 32515
rect 11435 32459 11521 32515
rect 11577 32459 11663 32515
rect 11719 32459 11805 32515
rect 11861 32459 11947 32515
rect 12003 32459 12089 32515
rect 12145 32459 12231 32515
rect 12287 32459 12373 32515
rect 12429 32459 12515 32515
rect 12571 32459 12657 32515
rect 12713 32459 12799 32515
rect 12855 32459 12941 32515
rect 12997 32459 13083 32515
rect 13139 32459 13225 32515
rect 13281 32459 13367 32515
rect 13423 32459 13509 32515
rect 13565 32459 13651 32515
rect 13707 32459 13793 32515
rect 13849 32459 13935 32515
rect 13991 32459 14077 32515
rect 14133 32459 14219 32515
rect 14275 32459 14361 32515
rect 14417 32459 14503 32515
rect 14559 32459 14645 32515
rect 14701 32459 14787 32515
rect 14843 32459 15000 32515
rect 0 32373 15000 32459
rect 0 32317 161 32373
rect 217 32317 303 32373
rect 359 32317 445 32373
rect 501 32317 587 32373
rect 643 32317 729 32373
rect 785 32317 871 32373
rect 927 32317 1013 32373
rect 1069 32317 1155 32373
rect 1211 32317 1297 32373
rect 1353 32317 1439 32373
rect 1495 32317 1581 32373
rect 1637 32317 1723 32373
rect 1779 32317 1865 32373
rect 1921 32317 2007 32373
rect 2063 32317 2149 32373
rect 2205 32317 2291 32373
rect 2347 32317 2433 32373
rect 2489 32317 2575 32373
rect 2631 32317 2717 32373
rect 2773 32317 2859 32373
rect 2915 32317 3001 32373
rect 3057 32317 3143 32373
rect 3199 32317 3285 32373
rect 3341 32317 3427 32373
rect 3483 32317 3569 32373
rect 3625 32317 3711 32373
rect 3767 32317 3853 32373
rect 3909 32317 3995 32373
rect 4051 32317 4137 32373
rect 4193 32317 4279 32373
rect 4335 32317 4421 32373
rect 4477 32317 4563 32373
rect 4619 32317 4705 32373
rect 4761 32317 4847 32373
rect 4903 32317 4989 32373
rect 5045 32317 5131 32373
rect 5187 32317 5273 32373
rect 5329 32317 5415 32373
rect 5471 32317 5557 32373
rect 5613 32317 5699 32373
rect 5755 32317 5841 32373
rect 5897 32317 5983 32373
rect 6039 32317 6125 32373
rect 6181 32317 6267 32373
rect 6323 32317 6409 32373
rect 6465 32317 6551 32373
rect 6607 32317 6693 32373
rect 6749 32317 6835 32373
rect 6891 32317 6977 32373
rect 7033 32317 7119 32373
rect 7175 32317 7261 32373
rect 7317 32317 7403 32373
rect 7459 32317 7545 32373
rect 7601 32317 7687 32373
rect 7743 32317 7829 32373
rect 7885 32317 7971 32373
rect 8027 32317 8113 32373
rect 8169 32317 8255 32373
rect 8311 32317 8397 32373
rect 8453 32317 8539 32373
rect 8595 32317 8681 32373
rect 8737 32317 8823 32373
rect 8879 32317 8965 32373
rect 9021 32317 9107 32373
rect 9163 32317 9249 32373
rect 9305 32317 9391 32373
rect 9447 32317 9533 32373
rect 9589 32317 9675 32373
rect 9731 32317 9817 32373
rect 9873 32317 9959 32373
rect 10015 32317 10101 32373
rect 10157 32317 10243 32373
rect 10299 32317 10385 32373
rect 10441 32317 10527 32373
rect 10583 32317 10669 32373
rect 10725 32317 10811 32373
rect 10867 32317 10953 32373
rect 11009 32317 11095 32373
rect 11151 32317 11237 32373
rect 11293 32317 11379 32373
rect 11435 32317 11521 32373
rect 11577 32317 11663 32373
rect 11719 32317 11805 32373
rect 11861 32317 11947 32373
rect 12003 32317 12089 32373
rect 12145 32317 12231 32373
rect 12287 32317 12373 32373
rect 12429 32317 12515 32373
rect 12571 32317 12657 32373
rect 12713 32317 12799 32373
rect 12855 32317 12941 32373
rect 12997 32317 13083 32373
rect 13139 32317 13225 32373
rect 13281 32317 13367 32373
rect 13423 32317 13509 32373
rect 13565 32317 13651 32373
rect 13707 32317 13793 32373
rect 13849 32317 13935 32373
rect 13991 32317 14077 32373
rect 14133 32317 14219 32373
rect 14275 32317 14361 32373
rect 14417 32317 14503 32373
rect 14559 32317 14645 32373
rect 14701 32317 14787 32373
rect 14843 32317 15000 32373
rect 0 32231 15000 32317
rect 0 32175 161 32231
rect 217 32175 303 32231
rect 359 32175 445 32231
rect 501 32175 587 32231
rect 643 32175 729 32231
rect 785 32175 871 32231
rect 927 32175 1013 32231
rect 1069 32175 1155 32231
rect 1211 32175 1297 32231
rect 1353 32175 1439 32231
rect 1495 32175 1581 32231
rect 1637 32175 1723 32231
rect 1779 32175 1865 32231
rect 1921 32175 2007 32231
rect 2063 32175 2149 32231
rect 2205 32175 2291 32231
rect 2347 32175 2433 32231
rect 2489 32175 2575 32231
rect 2631 32175 2717 32231
rect 2773 32175 2859 32231
rect 2915 32175 3001 32231
rect 3057 32175 3143 32231
rect 3199 32175 3285 32231
rect 3341 32175 3427 32231
rect 3483 32175 3569 32231
rect 3625 32175 3711 32231
rect 3767 32175 3853 32231
rect 3909 32175 3995 32231
rect 4051 32175 4137 32231
rect 4193 32175 4279 32231
rect 4335 32175 4421 32231
rect 4477 32175 4563 32231
rect 4619 32175 4705 32231
rect 4761 32175 4847 32231
rect 4903 32175 4989 32231
rect 5045 32175 5131 32231
rect 5187 32175 5273 32231
rect 5329 32175 5415 32231
rect 5471 32175 5557 32231
rect 5613 32175 5699 32231
rect 5755 32175 5841 32231
rect 5897 32175 5983 32231
rect 6039 32175 6125 32231
rect 6181 32175 6267 32231
rect 6323 32175 6409 32231
rect 6465 32175 6551 32231
rect 6607 32175 6693 32231
rect 6749 32175 6835 32231
rect 6891 32175 6977 32231
rect 7033 32175 7119 32231
rect 7175 32175 7261 32231
rect 7317 32175 7403 32231
rect 7459 32175 7545 32231
rect 7601 32175 7687 32231
rect 7743 32175 7829 32231
rect 7885 32175 7971 32231
rect 8027 32175 8113 32231
rect 8169 32175 8255 32231
rect 8311 32175 8397 32231
rect 8453 32175 8539 32231
rect 8595 32175 8681 32231
rect 8737 32175 8823 32231
rect 8879 32175 8965 32231
rect 9021 32175 9107 32231
rect 9163 32175 9249 32231
rect 9305 32175 9391 32231
rect 9447 32175 9533 32231
rect 9589 32175 9675 32231
rect 9731 32175 9817 32231
rect 9873 32175 9959 32231
rect 10015 32175 10101 32231
rect 10157 32175 10243 32231
rect 10299 32175 10385 32231
rect 10441 32175 10527 32231
rect 10583 32175 10669 32231
rect 10725 32175 10811 32231
rect 10867 32175 10953 32231
rect 11009 32175 11095 32231
rect 11151 32175 11237 32231
rect 11293 32175 11379 32231
rect 11435 32175 11521 32231
rect 11577 32175 11663 32231
rect 11719 32175 11805 32231
rect 11861 32175 11947 32231
rect 12003 32175 12089 32231
rect 12145 32175 12231 32231
rect 12287 32175 12373 32231
rect 12429 32175 12515 32231
rect 12571 32175 12657 32231
rect 12713 32175 12799 32231
rect 12855 32175 12941 32231
rect 12997 32175 13083 32231
rect 13139 32175 13225 32231
rect 13281 32175 13367 32231
rect 13423 32175 13509 32231
rect 13565 32175 13651 32231
rect 13707 32175 13793 32231
rect 13849 32175 13935 32231
rect 13991 32175 14077 32231
rect 14133 32175 14219 32231
rect 14275 32175 14361 32231
rect 14417 32175 14503 32231
rect 14559 32175 14645 32231
rect 14701 32175 14787 32231
rect 14843 32175 15000 32231
rect 0 32089 15000 32175
rect 0 32033 161 32089
rect 217 32033 303 32089
rect 359 32033 445 32089
rect 501 32033 587 32089
rect 643 32033 729 32089
rect 785 32033 871 32089
rect 927 32033 1013 32089
rect 1069 32033 1155 32089
rect 1211 32033 1297 32089
rect 1353 32033 1439 32089
rect 1495 32033 1581 32089
rect 1637 32033 1723 32089
rect 1779 32033 1865 32089
rect 1921 32033 2007 32089
rect 2063 32033 2149 32089
rect 2205 32033 2291 32089
rect 2347 32033 2433 32089
rect 2489 32033 2575 32089
rect 2631 32033 2717 32089
rect 2773 32033 2859 32089
rect 2915 32033 3001 32089
rect 3057 32033 3143 32089
rect 3199 32033 3285 32089
rect 3341 32033 3427 32089
rect 3483 32033 3569 32089
rect 3625 32033 3711 32089
rect 3767 32033 3853 32089
rect 3909 32033 3995 32089
rect 4051 32033 4137 32089
rect 4193 32033 4279 32089
rect 4335 32033 4421 32089
rect 4477 32033 4563 32089
rect 4619 32033 4705 32089
rect 4761 32033 4847 32089
rect 4903 32033 4989 32089
rect 5045 32033 5131 32089
rect 5187 32033 5273 32089
rect 5329 32033 5415 32089
rect 5471 32033 5557 32089
rect 5613 32033 5699 32089
rect 5755 32033 5841 32089
rect 5897 32033 5983 32089
rect 6039 32033 6125 32089
rect 6181 32033 6267 32089
rect 6323 32033 6409 32089
rect 6465 32033 6551 32089
rect 6607 32033 6693 32089
rect 6749 32033 6835 32089
rect 6891 32033 6977 32089
rect 7033 32033 7119 32089
rect 7175 32033 7261 32089
rect 7317 32033 7403 32089
rect 7459 32033 7545 32089
rect 7601 32033 7687 32089
rect 7743 32033 7829 32089
rect 7885 32033 7971 32089
rect 8027 32033 8113 32089
rect 8169 32033 8255 32089
rect 8311 32033 8397 32089
rect 8453 32033 8539 32089
rect 8595 32033 8681 32089
rect 8737 32033 8823 32089
rect 8879 32033 8965 32089
rect 9021 32033 9107 32089
rect 9163 32033 9249 32089
rect 9305 32033 9391 32089
rect 9447 32033 9533 32089
rect 9589 32033 9675 32089
rect 9731 32033 9817 32089
rect 9873 32033 9959 32089
rect 10015 32033 10101 32089
rect 10157 32033 10243 32089
rect 10299 32033 10385 32089
rect 10441 32033 10527 32089
rect 10583 32033 10669 32089
rect 10725 32033 10811 32089
rect 10867 32033 10953 32089
rect 11009 32033 11095 32089
rect 11151 32033 11237 32089
rect 11293 32033 11379 32089
rect 11435 32033 11521 32089
rect 11577 32033 11663 32089
rect 11719 32033 11805 32089
rect 11861 32033 11947 32089
rect 12003 32033 12089 32089
rect 12145 32033 12231 32089
rect 12287 32033 12373 32089
rect 12429 32033 12515 32089
rect 12571 32033 12657 32089
rect 12713 32033 12799 32089
rect 12855 32033 12941 32089
rect 12997 32033 13083 32089
rect 13139 32033 13225 32089
rect 13281 32033 13367 32089
rect 13423 32033 13509 32089
rect 13565 32033 13651 32089
rect 13707 32033 13793 32089
rect 13849 32033 13935 32089
rect 13991 32033 14077 32089
rect 14133 32033 14219 32089
rect 14275 32033 14361 32089
rect 14417 32033 14503 32089
rect 14559 32033 14645 32089
rect 14701 32033 14787 32089
rect 14843 32033 15000 32089
rect 0 31947 15000 32033
rect 0 31891 161 31947
rect 217 31891 303 31947
rect 359 31891 445 31947
rect 501 31891 587 31947
rect 643 31891 729 31947
rect 785 31891 871 31947
rect 927 31891 1013 31947
rect 1069 31891 1155 31947
rect 1211 31891 1297 31947
rect 1353 31891 1439 31947
rect 1495 31891 1581 31947
rect 1637 31891 1723 31947
rect 1779 31891 1865 31947
rect 1921 31891 2007 31947
rect 2063 31891 2149 31947
rect 2205 31891 2291 31947
rect 2347 31891 2433 31947
rect 2489 31891 2575 31947
rect 2631 31891 2717 31947
rect 2773 31891 2859 31947
rect 2915 31891 3001 31947
rect 3057 31891 3143 31947
rect 3199 31891 3285 31947
rect 3341 31891 3427 31947
rect 3483 31891 3569 31947
rect 3625 31891 3711 31947
rect 3767 31891 3853 31947
rect 3909 31891 3995 31947
rect 4051 31891 4137 31947
rect 4193 31891 4279 31947
rect 4335 31891 4421 31947
rect 4477 31891 4563 31947
rect 4619 31891 4705 31947
rect 4761 31891 4847 31947
rect 4903 31891 4989 31947
rect 5045 31891 5131 31947
rect 5187 31891 5273 31947
rect 5329 31891 5415 31947
rect 5471 31891 5557 31947
rect 5613 31891 5699 31947
rect 5755 31891 5841 31947
rect 5897 31891 5983 31947
rect 6039 31891 6125 31947
rect 6181 31891 6267 31947
rect 6323 31891 6409 31947
rect 6465 31891 6551 31947
rect 6607 31891 6693 31947
rect 6749 31891 6835 31947
rect 6891 31891 6977 31947
rect 7033 31891 7119 31947
rect 7175 31891 7261 31947
rect 7317 31891 7403 31947
rect 7459 31891 7545 31947
rect 7601 31891 7687 31947
rect 7743 31891 7829 31947
rect 7885 31891 7971 31947
rect 8027 31891 8113 31947
rect 8169 31891 8255 31947
rect 8311 31891 8397 31947
rect 8453 31891 8539 31947
rect 8595 31891 8681 31947
rect 8737 31891 8823 31947
rect 8879 31891 8965 31947
rect 9021 31891 9107 31947
rect 9163 31891 9249 31947
rect 9305 31891 9391 31947
rect 9447 31891 9533 31947
rect 9589 31891 9675 31947
rect 9731 31891 9817 31947
rect 9873 31891 9959 31947
rect 10015 31891 10101 31947
rect 10157 31891 10243 31947
rect 10299 31891 10385 31947
rect 10441 31891 10527 31947
rect 10583 31891 10669 31947
rect 10725 31891 10811 31947
rect 10867 31891 10953 31947
rect 11009 31891 11095 31947
rect 11151 31891 11237 31947
rect 11293 31891 11379 31947
rect 11435 31891 11521 31947
rect 11577 31891 11663 31947
rect 11719 31891 11805 31947
rect 11861 31891 11947 31947
rect 12003 31891 12089 31947
rect 12145 31891 12231 31947
rect 12287 31891 12373 31947
rect 12429 31891 12515 31947
rect 12571 31891 12657 31947
rect 12713 31891 12799 31947
rect 12855 31891 12941 31947
rect 12997 31891 13083 31947
rect 13139 31891 13225 31947
rect 13281 31891 13367 31947
rect 13423 31891 13509 31947
rect 13565 31891 13651 31947
rect 13707 31891 13793 31947
rect 13849 31891 13935 31947
rect 13991 31891 14077 31947
rect 14133 31891 14219 31947
rect 14275 31891 14361 31947
rect 14417 31891 14503 31947
rect 14559 31891 14645 31947
rect 14701 31891 14787 31947
rect 14843 31891 15000 31947
rect 0 31805 15000 31891
rect 0 31749 161 31805
rect 217 31749 303 31805
rect 359 31749 445 31805
rect 501 31749 587 31805
rect 643 31749 729 31805
rect 785 31749 871 31805
rect 927 31749 1013 31805
rect 1069 31749 1155 31805
rect 1211 31749 1297 31805
rect 1353 31749 1439 31805
rect 1495 31749 1581 31805
rect 1637 31749 1723 31805
rect 1779 31749 1865 31805
rect 1921 31749 2007 31805
rect 2063 31749 2149 31805
rect 2205 31749 2291 31805
rect 2347 31749 2433 31805
rect 2489 31749 2575 31805
rect 2631 31749 2717 31805
rect 2773 31749 2859 31805
rect 2915 31749 3001 31805
rect 3057 31749 3143 31805
rect 3199 31749 3285 31805
rect 3341 31749 3427 31805
rect 3483 31749 3569 31805
rect 3625 31749 3711 31805
rect 3767 31749 3853 31805
rect 3909 31749 3995 31805
rect 4051 31749 4137 31805
rect 4193 31749 4279 31805
rect 4335 31749 4421 31805
rect 4477 31749 4563 31805
rect 4619 31749 4705 31805
rect 4761 31749 4847 31805
rect 4903 31749 4989 31805
rect 5045 31749 5131 31805
rect 5187 31749 5273 31805
rect 5329 31749 5415 31805
rect 5471 31749 5557 31805
rect 5613 31749 5699 31805
rect 5755 31749 5841 31805
rect 5897 31749 5983 31805
rect 6039 31749 6125 31805
rect 6181 31749 6267 31805
rect 6323 31749 6409 31805
rect 6465 31749 6551 31805
rect 6607 31749 6693 31805
rect 6749 31749 6835 31805
rect 6891 31749 6977 31805
rect 7033 31749 7119 31805
rect 7175 31749 7261 31805
rect 7317 31749 7403 31805
rect 7459 31749 7545 31805
rect 7601 31749 7687 31805
rect 7743 31749 7829 31805
rect 7885 31749 7971 31805
rect 8027 31749 8113 31805
rect 8169 31749 8255 31805
rect 8311 31749 8397 31805
rect 8453 31749 8539 31805
rect 8595 31749 8681 31805
rect 8737 31749 8823 31805
rect 8879 31749 8965 31805
rect 9021 31749 9107 31805
rect 9163 31749 9249 31805
rect 9305 31749 9391 31805
rect 9447 31749 9533 31805
rect 9589 31749 9675 31805
rect 9731 31749 9817 31805
rect 9873 31749 9959 31805
rect 10015 31749 10101 31805
rect 10157 31749 10243 31805
rect 10299 31749 10385 31805
rect 10441 31749 10527 31805
rect 10583 31749 10669 31805
rect 10725 31749 10811 31805
rect 10867 31749 10953 31805
rect 11009 31749 11095 31805
rect 11151 31749 11237 31805
rect 11293 31749 11379 31805
rect 11435 31749 11521 31805
rect 11577 31749 11663 31805
rect 11719 31749 11805 31805
rect 11861 31749 11947 31805
rect 12003 31749 12089 31805
rect 12145 31749 12231 31805
rect 12287 31749 12373 31805
rect 12429 31749 12515 31805
rect 12571 31749 12657 31805
rect 12713 31749 12799 31805
rect 12855 31749 12941 31805
rect 12997 31749 13083 31805
rect 13139 31749 13225 31805
rect 13281 31749 13367 31805
rect 13423 31749 13509 31805
rect 13565 31749 13651 31805
rect 13707 31749 13793 31805
rect 13849 31749 13935 31805
rect 13991 31749 14077 31805
rect 14133 31749 14219 31805
rect 14275 31749 14361 31805
rect 14417 31749 14503 31805
rect 14559 31749 14645 31805
rect 14701 31749 14787 31805
rect 14843 31749 15000 31805
rect 0 31663 15000 31749
rect 0 31607 161 31663
rect 217 31607 303 31663
rect 359 31607 445 31663
rect 501 31607 587 31663
rect 643 31607 729 31663
rect 785 31607 871 31663
rect 927 31607 1013 31663
rect 1069 31607 1155 31663
rect 1211 31607 1297 31663
rect 1353 31607 1439 31663
rect 1495 31607 1581 31663
rect 1637 31607 1723 31663
rect 1779 31607 1865 31663
rect 1921 31607 2007 31663
rect 2063 31607 2149 31663
rect 2205 31607 2291 31663
rect 2347 31607 2433 31663
rect 2489 31607 2575 31663
rect 2631 31607 2717 31663
rect 2773 31607 2859 31663
rect 2915 31607 3001 31663
rect 3057 31607 3143 31663
rect 3199 31607 3285 31663
rect 3341 31607 3427 31663
rect 3483 31607 3569 31663
rect 3625 31607 3711 31663
rect 3767 31607 3853 31663
rect 3909 31607 3995 31663
rect 4051 31607 4137 31663
rect 4193 31607 4279 31663
rect 4335 31607 4421 31663
rect 4477 31607 4563 31663
rect 4619 31607 4705 31663
rect 4761 31607 4847 31663
rect 4903 31607 4989 31663
rect 5045 31607 5131 31663
rect 5187 31607 5273 31663
rect 5329 31607 5415 31663
rect 5471 31607 5557 31663
rect 5613 31607 5699 31663
rect 5755 31607 5841 31663
rect 5897 31607 5983 31663
rect 6039 31607 6125 31663
rect 6181 31607 6267 31663
rect 6323 31607 6409 31663
rect 6465 31607 6551 31663
rect 6607 31607 6693 31663
rect 6749 31607 6835 31663
rect 6891 31607 6977 31663
rect 7033 31607 7119 31663
rect 7175 31607 7261 31663
rect 7317 31607 7403 31663
rect 7459 31607 7545 31663
rect 7601 31607 7687 31663
rect 7743 31607 7829 31663
rect 7885 31607 7971 31663
rect 8027 31607 8113 31663
rect 8169 31607 8255 31663
rect 8311 31607 8397 31663
rect 8453 31607 8539 31663
rect 8595 31607 8681 31663
rect 8737 31607 8823 31663
rect 8879 31607 8965 31663
rect 9021 31607 9107 31663
rect 9163 31607 9249 31663
rect 9305 31607 9391 31663
rect 9447 31607 9533 31663
rect 9589 31607 9675 31663
rect 9731 31607 9817 31663
rect 9873 31607 9959 31663
rect 10015 31607 10101 31663
rect 10157 31607 10243 31663
rect 10299 31607 10385 31663
rect 10441 31607 10527 31663
rect 10583 31607 10669 31663
rect 10725 31607 10811 31663
rect 10867 31607 10953 31663
rect 11009 31607 11095 31663
rect 11151 31607 11237 31663
rect 11293 31607 11379 31663
rect 11435 31607 11521 31663
rect 11577 31607 11663 31663
rect 11719 31607 11805 31663
rect 11861 31607 11947 31663
rect 12003 31607 12089 31663
rect 12145 31607 12231 31663
rect 12287 31607 12373 31663
rect 12429 31607 12515 31663
rect 12571 31607 12657 31663
rect 12713 31607 12799 31663
rect 12855 31607 12941 31663
rect 12997 31607 13083 31663
rect 13139 31607 13225 31663
rect 13281 31607 13367 31663
rect 13423 31607 13509 31663
rect 13565 31607 13651 31663
rect 13707 31607 13793 31663
rect 13849 31607 13935 31663
rect 13991 31607 14077 31663
rect 14133 31607 14219 31663
rect 14275 31607 14361 31663
rect 14417 31607 14503 31663
rect 14559 31607 14645 31663
rect 14701 31607 14787 31663
rect 14843 31607 15000 31663
rect 0 31521 15000 31607
rect 0 31465 161 31521
rect 217 31465 303 31521
rect 359 31465 445 31521
rect 501 31465 587 31521
rect 643 31465 729 31521
rect 785 31465 871 31521
rect 927 31465 1013 31521
rect 1069 31465 1155 31521
rect 1211 31465 1297 31521
rect 1353 31465 1439 31521
rect 1495 31465 1581 31521
rect 1637 31465 1723 31521
rect 1779 31465 1865 31521
rect 1921 31465 2007 31521
rect 2063 31465 2149 31521
rect 2205 31465 2291 31521
rect 2347 31465 2433 31521
rect 2489 31465 2575 31521
rect 2631 31465 2717 31521
rect 2773 31465 2859 31521
rect 2915 31465 3001 31521
rect 3057 31465 3143 31521
rect 3199 31465 3285 31521
rect 3341 31465 3427 31521
rect 3483 31465 3569 31521
rect 3625 31465 3711 31521
rect 3767 31465 3853 31521
rect 3909 31465 3995 31521
rect 4051 31465 4137 31521
rect 4193 31465 4279 31521
rect 4335 31465 4421 31521
rect 4477 31465 4563 31521
rect 4619 31465 4705 31521
rect 4761 31465 4847 31521
rect 4903 31465 4989 31521
rect 5045 31465 5131 31521
rect 5187 31465 5273 31521
rect 5329 31465 5415 31521
rect 5471 31465 5557 31521
rect 5613 31465 5699 31521
rect 5755 31465 5841 31521
rect 5897 31465 5983 31521
rect 6039 31465 6125 31521
rect 6181 31465 6267 31521
rect 6323 31465 6409 31521
rect 6465 31465 6551 31521
rect 6607 31465 6693 31521
rect 6749 31465 6835 31521
rect 6891 31465 6977 31521
rect 7033 31465 7119 31521
rect 7175 31465 7261 31521
rect 7317 31465 7403 31521
rect 7459 31465 7545 31521
rect 7601 31465 7687 31521
rect 7743 31465 7829 31521
rect 7885 31465 7971 31521
rect 8027 31465 8113 31521
rect 8169 31465 8255 31521
rect 8311 31465 8397 31521
rect 8453 31465 8539 31521
rect 8595 31465 8681 31521
rect 8737 31465 8823 31521
rect 8879 31465 8965 31521
rect 9021 31465 9107 31521
rect 9163 31465 9249 31521
rect 9305 31465 9391 31521
rect 9447 31465 9533 31521
rect 9589 31465 9675 31521
rect 9731 31465 9817 31521
rect 9873 31465 9959 31521
rect 10015 31465 10101 31521
rect 10157 31465 10243 31521
rect 10299 31465 10385 31521
rect 10441 31465 10527 31521
rect 10583 31465 10669 31521
rect 10725 31465 10811 31521
rect 10867 31465 10953 31521
rect 11009 31465 11095 31521
rect 11151 31465 11237 31521
rect 11293 31465 11379 31521
rect 11435 31465 11521 31521
rect 11577 31465 11663 31521
rect 11719 31465 11805 31521
rect 11861 31465 11947 31521
rect 12003 31465 12089 31521
rect 12145 31465 12231 31521
rect 12287 31465 12373 31521
rect 12429 31465 12515 31521
rect 12571 31465 12657 31521
rect 12713 31465 12799 31521
rect 12855 31465 12941 31521
rect 12997 31465 13083 31521
rect 13139 31465 13225 31521
rect 13281 31465 13367 31521
rect 13423 31465 13509 31521
rect 13565 31465 13651 31521
rect 13707 31465 13793 31521
rect 13849 31465 13935 31521
rect 13991 31465 14077 31521
rect 14133 31465 14219 31521
rect 14275 31465 14361 31521
rect 14417 31465 14503 31521
rect 14559 31465 14645 31521
rect 14701 31465 14787 31521
rect 14843 31465 15000 31521
rect 0 31379 15000 31465
rect 0 31323 161 31379
rect 217 31323 303 31379
rect 359 31323 445 31379
rect 501 31323 587 31379
rect 643 31323 729 31379
rect 785 31323 871 31379
rect 927 31323 1013 31379
rect 1069 31323 1155 31379
rect 1211 31323 1297 31379
rect 1353 31323 1439 31379
rect 1495 31323 1581 31379
rect 1637 31323 1723 31379
rect 1779 31323 1865 31379
rect 1921 31323 2007 31379
rect 2063 31323 2149 31379
rect 2205 31323 2291 31379
rect 2347 31323 2433 31379
rect 2489 31323 2575 31379
rect 2631 31323 2717 31379
rect 2773 31323 2859 31379
rect 2915 31323 3001 31379
rect 3057 31323 3143 31379
rect 3199 31323 3285 31379
rect 3341 31323 3427 31379
rect 3483 31323 3569 31379
rect 3625 31323 3711 31379
rect 3767 31323 3853 31379
rect 3909 31323 3995 31379
rect 4051 31323 4137 31379
rect 4193 31323 4279 31379
rect 4335 31323 4421 31379
rect 4477 31323 4563 31379
rect 4619 31323 4705 31379
rect 4761 31323 4847 31379
rect 4903 31323 4989 31379
rect 5045 31323 5131 31379
rect 5187 31323 5273 31379
rect 5329 31323 5415 31379
rect 5471 31323 5557 31379
rect 5613 31323 5699 31379
rect 5755 31323 5841 31379
rect 5897 31323 5983 31379
rect 6039 31323 6125 31379
rect 6181 31323 6267 31379
rect 6323 31323 6409 31379
rect 6465 31323 6551 31379
rect 6607 31323 6693 31379
rect 6749 31323 6835 31379
rect 6891 31323 6977 31379
rect 7033 31323 7119 31379
rect 7175 31323 7261 31379
rect 7317 31323 7403 31379
rect 7459 31323 7545 31379
rect 7601 31323 7687 31379
rect 7743 31323 7829 31379
rect 7885 31323 7971 31379
rect 8027 31323 8113 31379
rect 8169 31323 8255 31379
rect 8311 31323 8397 31379
rect 8453 31323 8539 31379
rect 8595 31323 8681 31379
rect 8737 31323 8823 31379
rect 8879 31323 8965 31379
rect 9021 31323 9107 31379
rect 9163 31323 9249 31379
rect 9305 31323 9391 31379
rect 9447 31323 9533 31379
rect 9589 31323 9675 31379
rect 9731 31323 9817 31379
rect 9873 31323 9959 31379
rect 10015 31323 10101 31379
rect 10157 31323 10243 31379
rect 10299 31323 10385 31379
rect 10441 31323 10527 31379
rect 10583 31323 10669 31379
rect 10725 31323 10811 31379
rect 10867 31323 10953 31379
rect 11009 31323 11095 31379
rect 11151 31323 11237 31379
rect 11293 31323 11379 31379
rect 11435 31323 11521 31379
rect 11577 31323 11663 31379
rect 11719 31323 11805 31379
rect 11861 31323 11947 31379
rect 12003 31323 12089 31379
rect 12145 31323 12231 31379
rect 12287 31323 12373 31379
rect 12429 31323 12515 31379
rect 12571 31323 12657 31379
rect 12713 31323 12799 31379
rect 12855 31323 12941 31379
rect 12997 31323 13083 31379
rect 13139 31323 13225 31379
rect 13281 31323 13367 31379
rect 13423 31323 13509 31379
rect 13565 31323 13651 31379
rect 13707 31323 13793 31379
rect 13849 31323 13935 31379
rect 13991 31323 14077 31379
rect 14133 31323 14219 31379
rect 14275 31323 14361 31379
rect 14417 31323 14503 31379
rect 14559 31323 14645 31379
rect 14701 31323 14787 31379
rect 14843 31323 15000 31379
rect 0 31237 15000 31323
rect 0 31181 161 31237
rect 217 31181 303 31237
rect 359 31181 445 31237
rect 501 31181 587 31237
rect 643 31181 729 31237
rect 785 31181 871 31237
rect 927 31181 1013 31237
rect 1069 31181 1155 31237
rect 1211 31181 1297 31237
rect 1353 31181 1439 31237
rect 1495 31181 1581 31237
rect 1637 31181 1723 31237
rect 1779 31181 1865 31237
rect 1921 31181 2007 31237
rect 2063 31181 2149 31237
rect 2205 31181 2291 31237
rect 2347 31181 2433 31237
rect 2489 31181 2575 31237
rect 2631 31181 2717 31237
rect 2773 31181 2859 31237
rect 2915 31181 3001 31237
rect 3057 31181 3143 31237
rect 3199 31181 3285 31237
rect 3341 31181 3427 31237
rect 3483 31181 3569 31237
rect 3625 31181 3711 31237
rect 3767 31181 3853 31237
rect 3909 31181 3995 31237
rect 4051 31181 4137 31237
rect 4193 31181 4279 31237
rect 4335 31181 4421 31237
rect 4477 31181 4563 31237
rect 4619 31181 4705 31237
rect 4761 31181 4847 31237
rect 4903 31181 4989 31237
rect 5045 31181 5131 31237
rect 5187 31181 5273 31237
rect 5329 31181 5415 31237
rect 5471 31181 5557 31237
rect 5613 31181 5699 31237
rect 5755 31181 5841 31237
rect 5897 31181 5983 31237
rect 6039 31181 6125 31237
rect 6181 31181 6267 31237
rect 6323 31181 6409 31237
rect 6465 31181 6551 31237
rect 6607 31181 6693 31237
rect 6749 31181 6835 31237
rect 6891 31181 6977 31237
rect 7033 31181 7119 31237
rect 7175 31181 7261 31237
rect 7317 31181 7403 31237
rect 7459 31181 7545 31237
rect 7601 31181 7687 31237
rect 7743 31181 7829 31237
rect 7885 31181 7971 31237
rect 8027 31181 8113 31237
rect 8169 31181 8255 31237
rect 8311 31181 8397 31237
rect 8453 31181 8539 31237
rect 8595 31181 8681 31237
rect 8737 31181 8823 31237
rect 8879 31181 8965 31237
rect 9021 31181 9107 31237
rect 9163 31181 9249 31237
rect 9305 31181 9391 31237
rect 9447 31181 9533 31237
rect 9589 31181 9675 31237
rect 9731 31181 9817 31237
rect 9873 31181 9959 31237
rect 10015 31181 10101 31237
rect 10157 31181 10243 31237
rect 10299 31181 10385 31237
rect 10441 31181 10527 31237
rect 10583 31181 10669 31237
rect 10725 31181 10811 31237
rect 10867 31181 10953 31237
rect 11009 31181 11095 31237
rect 11151 31181 11237 31237
rect 11293 31181 11379 31237
rect 11435 31181 11521 31237
rect 11577 31181 11663 31237
rect 11719 31181 11805 31237
rect 11861 31181 11947 31237
rect 12003 31181 12089 31237
rect 12145 31181 12231 31237
rect 12287 31181 12373 31237
rect 12429 31181 12515 31237
rect 12571 31181 12657 31237
rect 12713 31181 12799 31237
rect 12855 31181 12941 31237
rect 12997 31181 13083 31237
rect 13139 31181 13225 31237
rect 13281 31181 13367 31237
rect 13423 31181 13509 31237
rect 13565 31181 13651 31237
rect 13707 31181 13793 31237
rect 13849 31181 13935 31237
rect 13991 31181 14077 31237
rect 14133 31181 14219 31237
rect 14275 31181 14361 31237
rect 14417 31181 14503 31237
rect 14559 31181 14645 31237
rect 14701 31181 14787 31237
rect 14843 31181 15000 31237
rect 0 31095 15000 31181
rect 0 31039 161 31095
rect 217 31039 303 31095
rect 359 31039 445 31095
rect 501 31039 587 31095
rect 643 31039 729 31095
rect 785 31039 871 31095
rect 927 31039 1013 31095
rect 1069 31039 1155 31095
rect 1211 31039 1297 31095
rect 1353 31039 1439 31095
rect 1495 31039 1581 31095
rect 1637 31039 1723 31095
rect 1779 31039 1865 31095
rect 1921 31039 2007 31095
rect 2063 31039 2149 31095
rect 2205 31039 2291 31095
rect 2347 31039 2433 31095
rect 2489 31039 2575 31095
rect 2631 31039 2717 31095
rect 2773 31039 2859 31095
rect 2915 31039 3001 31095
rect 3057 31039 3143 31095
rect 3199 31039 3285 31095
rect 3341 31039 3427 31095
rect 3483 31039 3569 31095
rect 3625 31039 3711 31095
rect 3767 31039 3853 31095
rect 3909 31039 3995 31095
rect 4051 31039 4137 31095
rect 4193 31039 4279 31095
rect 4335 31039 4421 31095
rect 4477 31039 4563 31095
rect 4619 31039 4705 31095
rect 4761 31039 4847 31095
rect 4903 31039 4989 31095
rect 5045 31039 5131 31095
rect 5187 31039 5273 31095
rect 5329 31039 5415 31095
rect 5471 31039 5557 31095
rect 5613 31039 5699 31095
rect 5755 31039 5841 31095
rect 5897 31039 5983 31095
rect 6039 31039 6125 31095
rect 6181 31039 6267 31095
rect 6323 31039 6409 31095
rect 6465 31039 6551 31095
rect 6607 31039 6693 31095
rect 6749 31039 6835 31095
rect 6891 31039 6977 31095
rect 7033 31039 7119 31095
rect 7175 31039 7261 31095
rect 7317 31039 7403 31095
rect 7459 31039 7545 31095
rect 7601 31039 7687 31095
rect 7743 31039 7829 31095
rect 7885 31039 7971 31095
rect 8027 31039 8113 31095
rect 8169 31039 8255 31095
rect 8311 31039 8397 31095
rect 8453 31039 8539 31095
rect 8595 31039 8681 31095
rect 8737 31039 8823 31095
rect 8879 31039 8965 31095
rect 9021 31039 9107 31095
rect 9163 31039 9249 31095
rect 9305 31039 9391 31095
rect 9447 31039 9533 31095
rect 9589 31039 9675 31095
rect 9731 31039 9817 31095
rect 9873 31039 9959 31095
rect 10015 31039 10101 31095
rect 10157 31039 10243 31095
rect 10299 31039 10385 31095
rect 10441 31039 10527 31095
rect 10583 31039 10669 31095
rect 10725 31039 10811 31095
rect 10867 31039 10953 31095
rect 11009 31039 11095 31095
rect 11151 31039 11237 31095
rect 11293 31039 11379 31095
rect 11435 31039 11521 31095
rect 11577 31039 11663 31095
rect 11719 31039 11805 31095
rect 11861 31039 11947 31095
rect 12003 31039 12089 31095
rect 12145 31039 12231 31095
rect 12287 31039 12373 31095
rect 12429 31039 12515 31095
rect 12571 31039 12657 31095
rect 12713 31039 12799 31095
rect 12855 31039 12941 31095
rect 12997 31039 13083 31095
rect 13139 31039 13225 31095
rect 13281 31039 13367 31095
rect 13423 31039 13509 31095
rect 13565 31039 13651 31095
rect 13707 31039 13793 31095
rect 13849 31039 13935 31095
rect 13991 31039 14077 31095
rect 14133 31039 14219 31095
rect 14275 31039 14361 31095
rect 14417 31039 14503 31095
rect 14559 31039 14645 31095
rect 14701 31039 14787 31095
rect 14843 31039 15000 31095
rect 0 30953 15000 31039
rect 0 30897 161 30953
rect 217 30897 303 30953
rect 359 30897 445 30953
rect 501 30897 587 30953
rect 643 30897 729 30953
rect 785 30897 871 30953
rect 927 30897 1013 30953
rect 1069 30897 1155 30953
rect 1211 30897 1297 30953
rect 1353 30897 1439 30953
rect 1495 30897 1581 30953
rect 1637 30897 1723 30953
rect 1779 30897 1865 30953
rect 1921 30897 2007 30953
rect 2063 30897 2149 30953
rect 2205 30897 2291 30953
rect 2347 30897 2433 30953
rect 2489 30897 2575 30953
rect 2631 30897 2717 30953
rect 2773 30897 2859 30953
rect 2915 30897 3001 30953
rect 3057 30897 3143 30953
rect 3199 30897 3285 30953
rect 3341 30897 3427 30953
rect 3483 30897 3569 30953
rect 3625 30897 3711 30953
rect 3767 30897 3853 30953
rect 3909 30897 3995 30953
rect 4051 30897 4137 30953
rect 4193 30897 4279 30953
rect 4335 30897 4421 30953
rect 4477 30897 4563 30953
rect 4619 30897 4705 30953
rect 4761 30897 4847 30953
rect 4903 30897 4989 30953
rect 5045 30897 5131 30953
rect 5187 30897 5273 30953
rect 5329 30897 5415 30953
rect 5471 30897 5557 30953
rect 5613 30897 5699 30953
rect 5755 30897 5841 30953
rect 5897 30897 5983 30953
rect 6039 30897 6125 30953
rect 6181 30897 6267 30953
rect 6323 30897 6409 30953
rect 6465 30897 6551 30953
rect 6607 30897 6693 30953
rect 6749 30897 6835 30953
rect 6891 30897 6977 30953
rect 7033 30897 7119 30953
rect 7175 30897 7261 30953
rect 7317 30897 7403 30953
rect 7459 30897 7545 30953
rect 7601 30897 7687 30953
rect 7743 30897 7829 30953
rect 7885 30897 7971 30953
rect 8027 30897 8113 30953
rect 8169 30897 8255 30953
rect 8311 30897 8397 30953
rect 8453 30897 8539 30953
rect 8595 30897 8681 30953
rect 8737 30897 8823 30953
rect 8879 30897 8965 30953
rect 9021 30897 9107 30953
rect 9163 30897 9249 30953
rect 9305 30897 9391 30953
rect 9447 30897 9533 30953
rect 9589 30897 9675 30953
rect 9731 30897 9817 30953
rect 9873 30897 9959 30953
rect 10015 30897 10101 30953
rect 10157 30897 10243 30953
rect 10299 30897 10385 30953
rect 10441 30897 10527 30953
rect 10583 30897 10669 30953
rect 10725 30897 10811 30953
rect 10867 30897 10953 30953
rect 11009 30897 11095 30953
rect 11151 30897 11237 30953
rect 11293 30897 11379 30953
rect 11435 30897 11521 30953
rect 11577 30897 11663 30953
rect 11719 30897 11805 30953
rect 11861 30897 11947 30953
rect 12003 30897 12089 30953
rect 12145 30897 12231 30953
rect 12287 30897 12373 30953
rect 12429 30897 12515 30953
rect 12571 30897 12657 30953
rect 12713 30897 12799 30953
rect 12855 30897 12941 30953
rect 12997 30897 13083 30953
rect 13139 30897 13225 30953
rect 13281 30897 13367 30953
rect 13423 30897 13509 30953
rect 13565 30897 13651 30953
rect 13707 30897 13793 30953
rect 13849 30897 13935 30953
rect 13991 30897 14077 30953
rect 14133 30897 14219 30953
rect 14275 30897 14361 30953
rect 14417 30897 14503 30953
rect 14559 30897 14645 30953
rect 14701 30897 14787 30953
rect 14843 30897 15000 30953
rect 0 30811 15000 30897
rect 0 30755 161 30811
rect 217 30755 303 30811
rect 359 30755 445 30811
rect 501 30755 587 30811
rect 643 30755 729 30811
rect 785 30755 871 30811
rect 927 30755 1013 30811
rect 1069 30755 1155 30811
rect 1211 30755 1297 30811
rect 1353 30755 1439 30811
rect 1495 30755 1581 30811
rect 1637 30755 1723 30811
rect 1779 30755 1865 30811
rect 1921 30755 2007 30811
rect 2063 30755 2149 30811
rect 2205 30755 2291 30811
rect 2347 30755 2433 30811
rect 2489 30755 2575 30811
rect 2631 30755 2717 30811
rect 2773 30755 2859 30811
rect 2915 30755 3001 30811
rect 3057 30755 3143 30811
rect 3199 30755 3285 30811
rect 3341 30755 3427 30811
rect 3483 30755 3569 30811
rect 3625 30755 3711 30811
rect 3767 30755 3853 30811
rect 3909 30755 3995 30811
rect 4051 30755 4137 30811
rect 4193 30755 4279 30811
rect 4335 30755 4421 30811
rect 4477 30755 4563 30811
rect 4619 30755 4705 30811
rect 4761 30755 4847 30811
rect 4903 30755 4989 30811
rect 5045 30755 5131 30811
rect 5187 30755 5273 30811
rect 5329 30755 5415 30811
rect 5471 30755 5557 30811
rect 5613 30755 5699 30811
rect 5755 30755 5841 30811
rect 5897 30755 5983 30811
rect 6039 30755 6125 30811
rect 6181 30755 6267 30811
rect 6323 30755 6409 30811
rect 6465 30755 6551 30811
rect 6607 30755 6693 30811
rect 6749 30755 6835 30811
rect 6891 30755 6977 30811
rect 7033 30755 7119 30811
rect 7175 30755 7261 30811
rect 7317 30755 7403 30811
rect 7459 30755 7545 30811
rect 7601 30755 7687 30811
rect 7743 30755 7829 30811
rect 7885 30755 7971 30811
rect 8027 30755 8113 30811
rect 8169 30755 8255 30811
rect 8311 30755 8397 30811
rect 8453 30755 8539 30811
rect 8595 30755 8681 30811
rect 8737 30755 8823 30811
rect 8879 30755 8965 30811
rect 9021 30755 9107 30811
rect 9163 30755 9249 30811
rect 9305 30755 9391 30811
rect 9447 30755 9533 30811
rect 9589 30755 9675 30811
rect 9731 30755 9817 30811
rect 9873 30755 9959 30811
rect 10015 30755 10101 30811
rect 10157 30755 10243 30811
rect 10299 30755 10385 30811
rect 10441 30755 10527 30811
rect 10583 30755 10669 30811
rect 10725 30755 10811 30811
rect 10867 30755 10953 30811
rect 11009 30755 11095 30811
rect 11151 30755 11237 30811
rect 11293 30755 11379 30811
rect 11435 30755 11521 30811
rect 11577 30755 11663 30811
rect 11719 30755 11805 30811
rect 11861 30755 11947 30811
rect 12003 30755 12089 30811
rect 12145 30755 12231 30811
rect 12287 30755 12373 30811
rect 12429 30755 12515 30811
rect 12571 30755 12657 30811
rect 12713 30755 12799 30811
rect 12855 30755 12941 30811
rect 12997 30755 13083 30811
rect 13139 30755 13225 30811
rect 13281 30755 13367 30811
rect 13423 30755 13509 30811
rect 13565 30755 13651 30811
rect 13707 30755 13793 30811
rect 13849 30755 13935 30811
rect 13991 30755 14077 30811
rect 14133 30755 14219 30811
rect 14275 30755 14361 30811
rect 14417 30755 14503 30811
rect 14559 30755 14645 30811
rect 14701 30755 14787 30811
rect 14843 30755 15000 30811
rect 0 30669 15000 30755
rect 0 30613 161 30669
rect 217 30613 303 30669
rect 359 30613 445 30669
rect 501 30613 587 30669
rect 643 30613 729 30669
rect 785 30613 871 30669
rect 927 30613 1013 30669
rect 1069 30613 1155 30669
rect 1211 30613 1297 30669
rect 1353 30613 1439 30669
rect 1495 30613 1581 30669
rect 1637 30613 1723 30669
rect 1779 30613 1865 30669
rect 1921 30613 2007 30669
rect 2063 30613 2149 30669
rect 2205 30613 2291 30669
rect 2347 30613 2433 30669
rect 2489 30613 2575 30669
rect 2631 30613 2717 30669
rect 2773 30613 2859 30669
rect 2915 30613 3001 30669
rect 3057 30613 3143 30669
rect 3199 30613 3285 30669
rect 3341 30613 3427 30669
rect 3483 30613 3569 30669
rect 3625 30613 3711 30669
rect 3767 30613 3853 30669
rect 3909 30613 3995 30669
rect 4051 30613 4137 30669
rect 4193 30613 4279 30669
rect 4335 30613 4421 30669
rect 4477 30613 4563 30669
rect 4619 30613 4705 30669
rect 4761 30613 4847 30669
rect 4903 30613 4989 30669
rect 5045 30613 5131 30669
rect 5187 30613 5273 30669
rect 5329 30613 5415 30669
rect 5471 30613 5557 30669
rect 5613 30613 5699 30669
rect 5755 30613 5841 30669
rect 5897 30613 5983 30669
rect 6039 30613 6125 30669
rect 6181 30613 6267 30669
rect 6323 30613 6409 30669
rect 6465 30613 6551 30669
rect 6607 30613 6693 30669
rect 6749 30613 6835 30669
rect 6891 30613 6977 30669
rect 7033 30613 7119 30669
rect 7175 30613 7261 30669
rect 7317 30613 7403 30669
rect 7459 30613 7545 30669
rect 7601 30613 7687 30669
rect 7743 30613 7829 30669
rect 7885 30613 7971 30669
rect 8027 30613 8113 30669
rect 8169 30613 8255 30669
rect 8311 30613 8397 30669
rect 8453 30613 8539 30669
rect 8595 30613 8681 30669
rect 8737 30613 8823 30669
rect 8879 30613 8965 30669
rect 9021 30613 9107 30669
rect 9163 30613 9249 30669
rect 9305 30613 9391 30669
rect 9447 30613 9533 30669
rect 9589 30613 9675 30669
rect 9731 30613 9817 30669
rect 9873 30613 9959 30669
rect 10015 30613 10101 30669
rect 10157 30613 10243 30669
rect 10299 30613 10385 30669
rect 10441 30613 10527 30669
rect 10583 30613 10669 30669
rect 10725 30613 10811 30669
rect 10867 30613 10953 30669
rect 11009 30613 11095 30669
rect 11151 30613 11237 30669
rect 11293 30613 11379 30669
rect 11435 30613 11521 30669
rect 11577 30613 11663 30669
rect 11719 30613 11805 30669
rect 11861 30613 11947 30669
rect 12003 30613 12089 30669
rect 12145 30613 12231 30669
rect 12287 30613 12373 30669
rect 12429 30613 12515 30669
rect 12571 30613 12657 30669
rect 12713 30613 12799 30669
rect 12855 30613 12941 30669
rect 12997 30613 13083 30669
rect 13139 30613 13225 30669
rect 13281 30613 13367 30669
rect 13423 30613 13509 30669
rect 13565 30613 13651 30669
rect 13707 30613 13793 30669
rect 13849 30613 13935 30669
rect 13991 30613 14077 30669
rect 14133 30613 14219 30669
rect 14275 30613 14361 30669
rect 14417 30613 14503 30669
rect 14559 30613 14645 30669
rect 14701 30613 14787 30669
rect 14843 30613 15000 30669
rect 0 30527 15000 30613
rect 0 30471 161 30527
rect 217 30471 303 30527
rect 359 30471 445 30527
rect 501 30471 587 30527
rect 643 30471 729 30527
rect 785 30471 871 30527
rect 927 30471 1013 30527
rect 1069 30471 1155 30527
rect 1211 30471 1297 30527
rect 1353 30471 1439 30527
rect 1495 30471 1581 30527
rect 1637 30471 1723 30527
rect 1779 30471 1865 30527
rect 1921 30471 2007 30527
rect 2063 30471 2149 30527
rect 2205 30471 2291 30527
rect 2347 30471 2433 30527
rect 2489 30471 2575 30527
rect 2631 30471 2717 30527
rect 2773 30471 2859 30527
rect 2915 30471 3001 30527
rect 3057 30471 3143 30527
rect 3199 30471 3285 30527
rect 3341 30471 3427 30527
rect 3483 30471 3569 30527
rect 3625 30471 3711 30527
rect 3767 30471 3853 30527
rect 3909 30471 3995 30527
rect 4051 30471 4137 30527
rect 4193 30471 4279 30527
rect 4335 30471 4421 30527
rect 4477 30471 4563 30527
rect 4619 30471 4705 30527
rect 4761 30471 4847 30527
rect 4903 30471 4989 30527
rect 5045 30471 5131 30527
rect 5187 30471 5273 30527
rect 5329 30471 5415 30527
rect 5471 30471 5557 30527
rect 5613 30471 5699 30527
rect 5755 30471 5841 30527
rect 5897 30471 5983 30527
rect 6039 30471 6125 30527
rect 6181 30471 6267 30527
rect 6323 30471 6409 30527
rect 6465 30471 6551 30527
rect 6607 30471 6693 30527
rect 6749 30471 6835 30527
rect 6891 30471 6977 30527
rect 7033 30471 7119 30527
rect 7175 30471 7261 30527
rect 7317 30471 7403 30527
rect 7459 30471 7545 30527
rect 7601 30471 7687 30527
rect 7743 30471 7829 30527
rect 7885 30471 7971 30527
rect 8027 30471 8113 30527
rect 8169 30471 8255 30527
rect 8311 30471 8397 30527
rect 8453 30471 8539 30527
rect 8595 30471 8681 30527
rect 8737 30471 8823 30527
rect 8879 30471 8965 30527
rect 9021 30471 9107 30527
rect 9163 30471 9249 30527
rect 9305 30471 9391 30527
rect 9447 30471 9533 30527
rect 9589 30471 9675 30527
rect 9731 30471 9817 30527
rect 9873 30471 9959 30527
rect 10015 30471 10101 30527
rect 10157 30471 10243 30527
rect 10299 30471 10385 30527
rect 10441 30471 10527 30527
rect 10583 30471 10669 30527
rect 10725 30471 10811 30527
rect 10867 30471 10953 30527
rect 11009 30471 11095 30527
rect 11151 30471 11237 30527
rect 11293 30471 11379 30527
rect 11435 30471 11521 30527
rect 11577 30471 11663 30527
rect 11719 30471 11805 30527
rect 11861 30471 11947 30527
rect 12003 30471 12089 30527
rect 12145 30471 12231 30527
rect 12287 30471 12373 30527
rect 12429 30471 12515 30527
rect 12571 30471 12657 30527
rect 12713 30471 12799 30527
rect 12855 30471 12941 30527
rect 12997 30471 13083 30527
rect 13139 30471 13225 30527
rect 13281 30471 13367 30527
rect 13423 30471 13509 30527
rect 13565 30471 13651 30527
rect 13707 30471 13793 30527
rect 13849 30471 13935 30527
rect 13991 30471 14077 30527
rect 14133 30471 14219 30527
rect 14275 30471 14361 30527
rect 14417 30471 14503 30527
rect 14559 30471 14645 30527
rect 14701 30471 14787 30527
rect 14843 30471 15000 30527
rect 0 30385 15000 30471
rect 0 30329 161 30385
rect 217 30329 303 30385
rect 359 30329 445 30385
rect 501 30329 587 30385
rect 643 30329 729 30385
rect 785 30329 871 30385
rect 927 30329 1013 30385
rect 1069 30329 1155 30385
rect 1211 30329 1297 30385
rect 1353 30329 1439 30385
rect 1495 30329 1581 30385
rect 1637 30329 1723 30385
rect 1779 30329 1865 30385
rect 1921 30329 2007 30385
rect 2063 30329 2149 30385
rect 2205 30329 2291 30385
rect 2347 30329 2433 30385
rect 2489 30329 2575 30385
rect 2631 30329 2717 30385
rect 2773 30329 2859 30385
rect 2915 30329 3001 30385
rect 3057 30329 3143 30385
rect 3199 30329 3285 30385
rect 3341 30329 3427 30385
rect 3483 30329 3569 30385
rect 3625 30329 3711 30385
rect 3767 30329 3853 30385
rect 3909 30329 3995 30385
rect 4051 30329 4137 30385
rect 4193 30329 4279 30385
rect 4335 30329 4421 30385
rect 4477 30329 4563 30385
rect 4619 30329 4705 30385
rect 4761 30329 4847 30385
rect 4903 30329 4989 30385
rect 5045 30329 5131 30385
rect 5187 30329 5273 30385
rect 5329 30329 5415 30385
rect 5471 30329 5557 30385
rect 5613 30329 5699 30385
rect 5755 30329 5841 30385
rect 5897 30329 5983 30385
rect 6039 30329 6125 30385
rect 6181 30329 6267 30385
rect 6323 30329 6409 30385
rect 6465 30329 6551 30385
rect 6607 30329 6693 30385
rect 6749 30329 6835 30385
rect 6891 30329 6977 30385
rect 7033 30329 7119 30385
rect 7175 30329 7261 30385
rect 7317 30329 7403 30385
rect 7459 30329 7545 30385
rect 7601 30329 7687 30385
rect 7743 30329 7829 30385
rect 7885 30329 7971 30385
rect 8027 30329 8113 30385
rect 8169 30329 8255 30385
rect 8311 30329 8397 30385
rect 8453 30329 8539 30385
rect 8595 30329 8681 30385
rect 8737 30329 8823 30385
rect 8879 30329 8965 30385
rect 9021 30329 9107 30385
rect 9163 30329 9249 30385
rect 9305 30329 9391 30385
rect 9447 30329 9533 30385
rect 9589 30329 9675 30385
rect 9731 30329 9817 30385
rect 9873 30329 9959 30385
rect 10015 30329 10101 30385
rect 10157 30329 10243 30385
rect 10299 30329 10385 30385
rect 10441 30329 10527 30385
rect 10583 30329 10669 30385
rect 10725 30329 10811 30385
rect 10867 30329 10953 30385
rect 11009 30329 11095 30385
rect 11151 30329 11237 30385
rect 11293 30329 11379 30385
rect 11435 30329 11521 30385
rect 11577 30329 11663 30385
rect 11719 30329 11805 30385
rect 11861 30329 11947 30385
rect 12003 30329 12089 30385
rect 12145 30329 12231 30385
rect 12287 30329 12373 30385
rect 12429 30329 12515 30385
rect 12571 30329 12657 30385
rect 12713 30329 12799 30385
rect 12855 30329 12941 30385
rect 12997 30329 13083 30385
rect 13139 30329 13225 30385
rect 13281 30329 13367 30385
rect 13423 30329 13509 30385
rect 13565 30329 13651 30385
rect 13707 30329 13793 30385
rect 13849 30329 13935 30385
rect 13991 30329 14077 30385
rect 14133 30329 14219 30385
rect 14275 30329 14361 30385
rect 14417 30329 14503 30385
rect 14559 30329 14645 30385
rect 14701 30329 14787 30385
rect 14843 30329 15000 30385
rect 0 30243 15000 30329
rect 0 30187 161 30243
rect 217 30187 303 30243
rect 359 30187 445 30243
rect 501 30187 587 30243
rect 643 30187 729 30243
rect 785 30187 871 30243
rect 927 30187 1013 30243
rect 1069 30187 1155 30243
rect 1211 30187 1297 30243
rect 1353 30187 1439 30243
rect 1495 30187 1581 30243
rect 1637 30187 1723 30243
rect 1779 30187 1865 30243
rect 1921 30187 2007 30243
rect 2063 30187 2149 30243
rect 2205 30187 2291 30243
rect 2347 30187 2433 30243
rect 2489 30187 2575 30243
rect 2631 30187 2717 30243
rect 2773 30187 2859 30243
rect 2915 30187 3001 30243
rect 3057 30187 3143 30243
rect 3199 30187 3285 30243
rect 3341 30187 3427 30243
rect 3483 30187 3569 30243
rect 3625 30187 3711 30243
rect 3767 30187 3853 30243
rect 3909 30187 3995 30243
rect 4051 30187 4137 30243
rect 4193 30187 4279 30243
rect 4335 30187 4421 30243
rect 4477 30187 4563 30243
rect 4619 30187 4705 30243
rect 4761 30187 4847 30243
rect 4903 30187 4989 30243
rect 5045 30187 5131 30243
rect 5187 30187 5273 30243
rect 5329 30187 5415 30243
rect 5471 30187 5557 30243
rect 5613 30187 5699 30243
rect 5755 30187 5841 30243
rect 5897 30187 5983 30243
rect 6039 30187 6125 30243
rect 6181 30187 6267 30243
rect 6323 30187 6409 30243
rect 6465 30187 6551 30243
rect 6607 30187 6693 30243
rect 6749 30187 6835 30243
rect 6891 30187 6977 30243
rect 7033 30187 7119 30243
rect 7175 30187 7261 30243
rect 7317 30187 7403 30243
rect 7459 30187 7545 30243
rect 7601 30187 7687 30243
rect 7743 30187 7829 30243
rect 7885 30187 7971 30243
rect 8027 30187 8113 30243
rect 8169 30187 8255 30243
rect 8311 30187 8397 30243
rect 8453 30187 8539 30243
rect 8595 30187 8681 30243
rect 8737 30187 8823 30243
rect 8879 30187 8965 30243
rect 9021 30187 9107 30243
rect 9163 30187 9249 30243
rect 9305 30187 9391 30243
rect 9447 30187 9533 30243
rect 9589 30187 9675 30243
rect 9731 30187 9817 30243
rect 9873 30187 9959 30243
rect 10015 30187 10101 30243
rect 10157 30187 10243 30243
rect 10299 30187 10385 30243
rect 10441 30187 10527 30243
rect 10583 30187 10669 30243
rect 10725 30187 10811 30243
rect 10867 30187 10953 30243
rect 11009 30187 11095 30243
rect 11151 30187 11237 30243
rect 11293 30187 11379 30243
rect 11435 30187 11521 30243
rect 11577 30187 11663 30243
rect 11719 30187 11805 30243
rect 11861 30187 11947 30243
rect 12003 30187 12089 30243
rect 12145 30187 12231 30243
rect 12287 30187 12373 30243
rect 12429 30187 12515 30243
rect 12571 30187 12657 30243
rect 12713 30187 12799 30243
rect 12855 30187 12941 30243
rect 12997 30187 13083 30243
rect 13139 30187 13225 30243
rect 13281 30187 13367 30243
rect 13423 30187 13509 30243
rect 13565 30187 13651 30243
rect 13707 30187 13793 30243
rect 13849 30187 13935 30243
rect 13991 30187 14077 30243
rect 14133 30187 14219 30243
rect 14275 30187 14361 30243
rect 14417 30187 14503 30243
rect 14559 30187 14645 30243
rect 14701 30187 14787 30243
rect 14843 30187 15000 30243
rect 0 30101 15000 30187
rect 0 30045 161 30101
rect 217 30045 303 30101
rect 359 30045 445 30101
rect 501 30045 587 30101
rect 643 30045 729 30101
rect 785 30045 871 30101
rect 927 30045 1013 30101
rect 1069 30045 1155 30101
rect 1211 30045 1297 30101
rect 1353 30045 1439 30101
rect 1495 30045 1581 30101
rect 1637 30045 1723 30101
rect 1779 30045 1865 30101
rect 1921 30045 2007 30101
rect 2063 30045 2149 30101
rect 2205 30045 2291 30101
rect 2347 30045 2433 30101
rect 2489 30045 2575 30101
rect 2631 30045 2717 30101
rect 2773 30045 2859 30101
rect 2915 30045 3001 30101
rect 3057 30045 3143 30101
rect 3199 30045 3285 30101
rect 3341 30045 3427 30101
rect 3483 30045 3569 30101
rect 3625 30045 3711 30101
rect 3767 30045 3853 30101
rect 3909 30045 3995 30101
rect 4051 30045 4137 30101
rect 4193 30045 4279 30101
rect 4335 30045 4421 30101
rect 4477 30045 4563 30101
rect 4619 30045 4705 30101
rect 4761 30045 4847 30101
rect 4903 30045 4989 30101
rect 5045 30045 5131 30101
rect 5187 30045 5273 30101
rect 5329 30045 5415 30101
rect 5471 30045 5557 30101
rect 5613 30045 5699 30101
rect 5755 30045 5841 30101
rect 5897 30045 5983 30101
rect 6039 30045 6125 30101
rect 6181 30045 6267 30101
rect 6323 30045 6409 30101
rect 6465 30045 6551 30101
rect 6607 30045 6693 30101
rect 6749 30045 6835 30101
rect 6891 30045 6977 30101
rect 7033 30045 7119 30101
rect 7175 30045 7261 30101
rect 7317 30045 7403 30101
rect 7459 30045 7545 30101
rect 7601 30045 7687 30101
rect 7743 30045 7829 30101
rect 7885 30045 7971 30101
rect 8027 30045 8113 30101
rect 8169 30045 8255 30101
rect 8311 30045 8397 30101
rect 8453 30045 8539 30101
rect 8595 30045 8681 30101
rect 8737 30045 8823 30101
rect 8879 30045 8965 30101
rect 9021 30045 9107 30101
rect 9163 30045 9249 30101
rect 9305 30045 9391 30101
rect 9447 30045 9533 30101
rect 9589 30045 9675 30101
rect 9731 30045 9817 30101
rect 9873 30045 9959 30101
rect 10015 30045 10101 30101
rect 10157 30045 10243 30101
rect 10299 30045 10385 30101
rect 10441 30045 10527 30101
rect 10583 30045 10669 30101
rect 10725 30045 10811 30101
rect 10867 30045 10953 30101
rect 11009 30045 11095 30101
rect 11151 30045 11237 30101
rect 11293 30045 11379 30101
rect 11435 30045 11521 30101
rect 11577 30045 11663 30101
rect 11719 30045 11805 30101
rect 11861 30045 11947 30101
rect 12003 30045 12089 30101
rect 12145 30045 12231 30101
rect 12287 30045 12373 30101
rect 12429 30045 12515 30101
rect 12571 30045 12657 30101
rect 12713 30045 12799 30101
rect 12855 30045 12941 30101
rect 12997 30045 13083 30101
rect 13139 30045 13225 30101
rect 13281 30045 13367 30101
rect 13423 30045 13509 30101
rect 13565 30045 13651 30101
rect 13707 30045 13793 30101
rect 13849 30045 13935 30101
rect 13991 30045 14077 30101
rect 14133 30045 14219 30101
rect 14275 30045 14361 30101
rect 14417 30045 14503 30101
rect 14559 30045 14645 30101
rect 14701 30045 14787 30101
rect 14843 30045 15000 30101
rect 0 30000 15000 30045
rect 937 29800 3937 30000
rect 4337 29800 7337 30000
rect 7737 29800 10737 30000
rect 11137 29800 14137 30000
rect 0 29741 15000 29800
rect 0 29685 161 29741
rect 217 29685 303 29741
rect 359 29685 445 29741
rect 501 29685 587 29741
rect 643 29685 729 29741
rect 785 29685 871 29741
rect 927 29685 1013 29741
rect 1069 29685 1155 29741
rect 1211 29685 1297 29741
rect 1353 29685 1439 29741
rect 1495 29685 1581 29741
rect 1637 29685 1723 29741
rect 1779 29685 1865 29741
rect 1921 29685 2007 29741
rect 2063 29685 2149 29741
rect 2205 29685 2291 29741
rect 2347 29685 2433 29741
rect 2489 29685 2575 29741
rect 2631 29685 2717 29741
rect 2773 29685 2859 29741
rect 2915 29685 3001 29741
rect 3057 29685 3143 29741
rect 3199 29685 3285 29741
rect 3341 29685 3427 29741
rect 3483 29685 3569 29741
rect 3625 29685 3711 29741
rect 3767 29685 3853 29741
rect 3909 29685 3995 29741
rect 4051 29685 4137 29741
rect 4193 29685 4279 29741
rect 4335 29685 4421 29741
rect 4477 29685 4563 29741
rect 4619 29685 4705 29741
rect 4761 29685 4847 29741
rect 4903 29685 4989 29741
rect 5045 29685 5131 29741
rect 5187 29685 5273 29741
rect 5329 29685 5415 29741
rect 5471 29685 5557 29741
rect 5613 29685 5699 29741
rect 5755 29685 5841 29741
rect 5897 29685 5983 29741
rect 6039 29685 6125 29741
rect 6181 29685 6267 29741
rect 6323 29685 6409 29741
rect 6465 29685 6551 29741
rect 6607 29685 6693 29741
rect 6749 29685 6835 29741
rect 6891 29685 6977 29741
rect 7033 29685 7119 29741
rect 7175 29685 7261 29741
rect 7317 29685 7403 29741
rect 7459 29685 7545 29741
rect 7601 29685 7687 29741
rect 7743 29685 7829 29741
rect 7885 29685 7971 29741
rect 8027 29685 8113 29741
rect 8169 29685 8255 29741
rect 8311 29685 8397 29741
rect 8453 29685 8539 29741
rect 8595 29685 8681 29741
rect 8737 29685 8823 29741
rect 8879 29685 8965 29741
rect 9021 29685 9107 29741
rect 9163 29685 9249 29741
rect 9305 29685 9391 29741
rect 9447 29685 9533 29741
rect 9589 29685 9675 29741
rect 9731 29685 9817 29741
rect 9873 29685 9959 29741
rect 10015 29685 10101 29741
rect 10157 29685 10243 29741
rect 10299 29685 10385 29741
rect 10441 29685 10527 29741
rect 10583 29685 10669 29741
rect 10725 29685 10811 29741
rect 10867 29685 10953 29741
rect 11009 29685 11095 29741
rect 11151 29685 11237 29741
rect 11293 29685 11379 29741
rect 11435 29685 11521 29741
rect 11577 29685 11663 29741
rect 11719 29685 11805 29741
rect 11861 29685 11947 29741
rect 12003 29685 12089 29741
rect 12145 29685 12231 29741
rect 12287 29685 12373 29741
rect 12429 29685 12515 29741
rect 12571 29685 12657 29741
rect 12713 29685 12799 29741
rect 12855 29685 12941 29741
rect 12997 29685 13083 29741
rect 13139 29685 13225 29741
rect 13281 29685 13367 29741
rect 13423 29685 13509 29741
rect 13565 29685 13651 29741
rect 13707 29685 13793 29741
rect 13849 29685 13935 29741
rect 13991 29685 14077 29741
rect 14133 29685 14219 29741
rect 14275 29685 14361 29741
rect 14417 29685 14503 29741
rect 14559 29685 14645 29741
rect 14701 29685 14787 29741
rect 14843 29685 15000 29741
rect 0 29599 15000 29685
rect 0 29543 161 29599
rect 217 29543 303 29599
rect 359 29543 445 29599
rect 501 29543 587 29599
rect 643 29543 729 29599
rect 785 29543 871 29599
rect 927 29543 1013 29599
rect 1069 29543 1155 29599
rect 1211 29543 1297 29599
rect 1353 29543 1439 29599
rect 1495 29543 1581 29599
rect 1637 29543 1723 29599
rect 1779 29543 1865 29599
rect 1921 29543 2007 29599
rect 2063 29543 2149 29599
rect 2205 29543 2291 29599
rect 2347 29543 2433 29599
rect 2489 29543 2575 29599
rect 2631 29543 2717 29599
rect 2773 29543 2859 29599
rect 2915 29543 3001 29599
rect 3057 29543 3143 29599
rect 3199 29543 3285 29599
rect 3341 29543 3427 29599
rect 3483 29543 3569 29599
rect 3625 29543 3711 29599
rect 3767 29543 3853 29599
rect 3909 29543 3995 29599
rect 4051 29543 4137 29599
rect 4193 29543 4279 29599
rect 4335 29543 4421 29599
rect 4477 29543 4563 29599
rect 4619 29543 4705 29599
rect 4761 29543 4847 29599
rect 4903 29543 4989 29599
rect 5045 29543 5131 29599
rect 5187 29543 5273 29599
rect 5329 29543 5415 29599
rect 5471 29543 5557 29599
rect 5613 29543 5699 29599
rect 5755 29543 5841 29599
rect 5897 29543 5983 29599
rect 6039 29543 6125 29599
rect 6181 29543 6267 29599
rect 6323 29543 6409 29599
rect 6465 29543 6551 29599
rect 6607 29543 6693 29599
rect 6749 29543 6835 29599
rect 6891 29543 6977 29599
rect 7033 29543 7119 29599
rect 7175 29543 7261 29599
rect 7317 29543 7403 29599
rect 7459 29543 7545 29599
rect 7601 29543 7687 29599
rect 7743 29543 7829 29599
rect 7885 29543 7971 29599
rect 8027 29543 8113 29599
rect 8169 29543 8255 29599
rect 8311 29543 8397 29599
rect 8453 29543 8539 29599
rect 8595 29543 8681 29599
rect 8737 29543 8823 29599
rect 8879 29543 8965 29599
rect 9021 29543 9107 29599
rect 9163 29543 9249 29599
rect 9305 29543 9391 29599
rect 9447 29543 9533 29599
rect 9589 29543 9675 29599
rect 9731 29543 9817 29599
rect 9873 29543 9959 29599
rect 10015 29543 10101 29599
rect 10157 29543 10243 29599
rect 10299 29543 10385 29599
rect 10441 29543 10527 29599
rect 10583 29543 10669 29599
rect 10725 29543 10811 29599
rect 10867 29543 10953 29599
rect 11009 29543 11095 29599
rect 11151 29543 11237 29599
rect 11293 29543 11379 29599
rect 11435 29543 11521 29599
rect 11577 29543 11663 29599
rect 11719 29543 11805 29599
rect 11861 29543 11947 29599
rect 12003 29543 12089 29599
rect 12145 29543 12231 29599
rect 12287 29543 12373 29599
rect 12429 29543 12515 29599
rect 12571 29543 12657 29599
rect 12713 29543 12799 29599
rect 12855 29543 12941 29599
rect 12997 29543 13083 29599
rect 13139 29543 13225 29599
rect 13281 29543 13367 29599
rect 13423 29543 13509 29599
rect 13565 29543 13651 29599
rect 13707 29543 13793 29599
rect 13849 29543 13935 29599
rect 13991 29543 14077 29599
rect 14133 29543 14219 29599
rect 14275 29543 14361 29599
rect 14417 29543 14503 29599
rect 14559 29543 14645 29599
rect 14701 29543 14787 29599
rect 14843 29543 15000 29599
rect 0 29457 15000 29543
rect 0 29401 161 29457
rect 217 29401 303 29457
rect 359 29401 445 29457
rect 501 29401 587 29457
rect 643 29401 729 29457
rect 785 29401 871 29457
rect 927 29401 1013 29457
rect 1069 29401 1155 29457
rect 1211 29401 1297 29457
rect 1353 29401 1439 29457
rect 1495 29401 1581 29457
rect 1637 29401 1723 29457
rect 1779 29401 1865 29457
rect 1921 29401 2007 29457
rect 2063 29401 2149 29457
rect 2205 29401 2291 29457
rect 2347 29401 2433 29457
rect 2489 29401 2575 29457
rect 2631 29401 2717 29457
rect 2773 29401 2859 29457
rect 2915 29401 3001 29457
rect 3057 29401 3143 29457
rect 3199 29401 3285 29457
rect 3341 29401 3427 29457
rect 3483 29401 3569 29457
rect 3625 29401 3711 29457
rect 3767 29401 3853 29457
rect 3909 29401 3995 29457
rect 4051 29401 4137 29457
rect 4193 29401 4279 29457
rect 4335 29401 4421 29457
rect 4477 29401 4563 29457
rect 4619 29401 4705 29457
rect 4761 29401 4847 29457
rect 4903 29401 4989 29457
rect 5045 29401 5131 29457
rect 5187 29401 5273 29457
rect 5329 29401 5415 29457
rect 5471 29401 5557 29457
rect 5613 29401 5699 29457
rect 5755 29401 5841 29457
rect 5897 29401 5983 29457
rect 6039 29401 6125 29457
rect 6181 29401 6267 29457
rect 6323 29401 6409 29457
rect 6465 29401 6551 29457
rect 6607 29401 6693 29457
rect 6749 29401 6835 29457
rect 6891 29401 6977 29457
rect 7033 29401 7119 29457
rect 7175 29401 7261 29457
rect 7317 29401 7403 29457
rect 7459 29401 7545 29457
rect 7601 29401 7687 29457
rect 7743 29401 7829 29457
rect 7885 29401 7971 29457
rect 8027 29401 8113 29457
rect 8169 29401 8255 29457
rect 8311 29401 8397 29457
rect 8453 29401 8539 29457
rect 8595 29401 8681 29457
rect 8737 29401 8823 29457
rect 8879 29401 8965 29457
rect 9021 29401 9107 29457
rect 9163 29401 9249 29457
rect 9305 29401 9391 29457
rect 9447 29401 9533 29457
rect 9589 29401 9675 29457
rect 9731 29401 9817 29457
rect 9873 29401 9959 29457
rect 10015 29401 10101 29457
rect 10157 29401 10243 29457
rect 10299 29401 10385 29457
rect 10441 29401 10527 29457
rect 10583 29401 10669 29457
rect 10725 29401 10811 29457
rect 10867 29401 10953 29457
rect 11009 29401 11095 29457
rect 11151 29401 11237 29457
rect 11293 29401 11379 29457
rect 11435 29401 11521 29457
rect 11577 29401 11663 29457
rect 11719 29401 11805 29457
rect 11861 29401 11947 29457
rect 12003 29401 12089 29457
rect 12145 29401 12231 29457
rect 12287 29401 12373 29457
rect 12429 29401 12515 29457
rect 12571 29401 12657 29457
rect 12713 29401 12799 29457
rect 12855 29401 12941 29457
rect 12997 29401 13083 29457
rect 13139 29401 13225 29457
rect 13281 29401 13367 29457
rect 13423 29401 13509 29457
rect 13565 29401 13651 29457
rect 13707 29401 13793 29457
rect 13849 29401 13935 29457
rect 13991 29401 14077 29457
rect 14133 29401 14219 29457
rect 14275 29401 14361 29457
rect 14417 29401 14503 29457
rect 14559 29401 14645 29457
rect 14701 29401 14787 29457
rect 14843 29401 15000 29457
rect 0 29315 15000 29401
rect 0 29259 161 29315
rect 217 29259 303 29315
rect 359 29259 445 29315
rect 501 29259 587 29315
rect 643 29259 729 29315
rect 785 29259 871 29315
rect 927 29259 1013 29315
rect 1069 29259 1155 29315
rect 1211 29259 1297 29315
rect 1353 29259 1439 29315
rect 1495 29259 1581 29315
rect 1637 29259 1723 29315
rect 1779 29259 1865 29315
rect 1921 29259 2007 29315
rect 2063 29259 2149 29315
rect 2205 29259 2291 29315
rect 2347 29259 2433 29315
rect 2489 29259 2575 29315
rect 2631 29259 2717 29315
rect 2773 29259 2859 29315
rect 2915 29259 3001 29315
rect 3057 29259 3143 29315
rect 3199 29259 3285 29315
rect 3341 29259 3427 29315
rect 3483 29259 3569 29315
rect 3625 29259 3711 29315
rect 3767 29259 3853 29315
rect 3909 29259 3995 29315
rect 4051 29259 4137 29315
rect 4193 29259 4279 29315
rect 4335 29259 4421 29315
rect 4477 29259 4563 29315
rect 4619 29259 4705 29315
rect 4761 29259 4847 29315
rect 4903 29259 4989 29315
rect 5045 29259 5131 29315
rect 5187 29259 5273 29315
rect 5329 29259 5415 29315
rect 5471 29259 5557 29315
rect 5613 29259 5699 29315
rect 5755 29259 5841 29315
rect 5897 29259 5983 29315
rect 6039 29259 6125 29315
rect 6181 29259 6267 29315
rect 6323 29259 6409 29315
rect 6465 29259 6551 29315
rect 6607 29259 6693 29315
rect 6749 29259 6835 29315
rect 6891 29259 6977 29315
rect 7033 29259 7119 29315
rect 7175 29259 7261 29315
rect 7317 29259 7403 29315
rect 7459 29259 7545 29315
rect 7601 29259 7687 29315
rect 7743 29259 7829 29315
rect 7885 29259 7971 29315
rect 8027 29259 8113 29315
rect 8169 29259 8255 29315
rect 8311 29259 8397 29315
rect 8453 29259 8539 29315
rect 8595 29259 8681 29315
rect 8737 29259 8823 29315
rect 8879 29259 8965 29315
rect 9021 29259 9107 29315
rect 9163 29259 9249 29315
rect 9305 29259 9391 29315
rect 9447 29259 9533 29315
rect 9589 29259 9675 29315
rect 9731 29259 9817 29315
rect 9873 29259 9959 29315
rect 10015 29259 10101 29315
rect 10157 29259 10243 29315
rect 10299 29259 10385 29315
rect 10441 29259 10527 29315
rect 10583 29259 10669 29315
rect 10725 29259 10811 29315
rect 10867 29259 10953 29315
rect 11009 29259 11095 29315
rect 11151 29259 11237 29315
rect 11293 29259 11379 29315
rect 11435 29259 11521 29315
rect 11577 29259 11663 29315
rect 11719 29259 11805 29315
rect 11861 29259 11947 29315
rect 12003 29259 12089 29315
rect 12145 29259 12231 29315
rect 12287 29259 12373 29315
rect 12429 29259 12515 29315
rect 12571 29259 12657 29315
rect 12713 29259 12799 29315
rect 12855 29259 12941 29315
rect 12997 29259 13083 29315
rect 13139 29259 13225 29315
rect 13281 29259 13367 29315
rect 13423 29259 13509 29315
rect 13565 29259 13651 29315
rect 13707 29259 13793 29315
rect 13849 29259 13935 29315
rect 13991 29259 14077 29315
rect 14133 29259 14219 29315
rect 14275 29259 14361 29315
rect 14417 29259 14503 29315
rect 14559 29259 14645 29315
rect 14701 29259 14787 29315
rect 14843 29259 15000 29315
rect 0 29173 15000 29259
rect 0 29117 161 29173
rect 217 29117 303 29173
rect 359 29117 445 29173
rect 501 29117 587 29173
rect 643 29117 729 29173
rect 785 29117 871 29173
rect 927 29117 1013 29173
rect 1069 29117 1155 29173
rect 1211 29117 1297 29173
rect 1353 29117 1439 29173
rect 1495 29117 1581 29173
rect 1637 29117 1723 29173
rect 1779 29117 1865 29173
rect 1921 29117 2007 29173
rect 2063 29117 2149 29173
rect 2205 29117 2291 29173
rect 2347 29117 2433 29173
rect 2489 29117 2575 29173
rect 2631 29117 2717 29173
rect 2773 29117 2859 29173
rect 2915 29117 3001 29173
rect 3057 29117 3143 29173
rect 3199 29117 3285 29173
rect 3341 29117 3427 29173
rect 3483 29117 3569 29173
rect 3625 29117 3711 29173
rect 3767 29117 3853 29173
rect 3909 29117 3995 29173
rect 4051 29117 4137 29173
rect 4193 29117 4279 29173
rect 4335 29117 4421 29173
rect 4477 29117 4563 29173
rect 4619 29117 4705 29173
rect 4761 29117 4847 29173
rect 4903 29117 4989 29173
rect 5045 29117 5131 29173
rect 5187 29117 5273 29173
rect 5329 29117 5415 29173
rect 5471 29117 5557 29173
rect 5613 29117 5699 29173
rect 5755 29117 5841 29173
rect 5897 29117 5983 29173
rect 6039 29117 6125 29173
rect 6181 29117 6267 29173
rect 6323 29117 6409 29173
rect 6465 29117 6551 29173
rect 6607 29117 6693 29173
rect 6749 29117 6835 29173
rect 6891 29117 6977 29173
rect 7033 29117 7119 29173
rect 7175 29117 7261 29173
rect 7317 29117 7403 29173
rect 7459 29117 7545 29173
rect 7601 29117 7687 29173
rect 7743 29117 7829 29173
rect 7885 29117 7971 29173
rect 8027 29117 8113 29173
rect 8169 29117 8255 29173
rect 8311 29117 8397 29173
rect 8453 29117 8539 29173
rect 8595 29117 8681 29173
rect 8737 29117 8823 29173
rect 8879 29117 8965 29173
rect 9021 29117 9107 29173
rect 9163 29117 9249 29173
rect 9305 29117 9391 29173
rect 9447 29117 9533 29173
rect 9589 29117 9675 29173
rect 9731 29117 9817 29173
rect 9873 29117 9959 29173
rect 10015 29117 10101 29173
rect 10157 29117 10243 29173
rect 10299 29117 10385 29173
rect 10441 29117 10527 29173
rect 10583 29117 10669 29173
rect 10725 29117 10811 29173
rect 10867 29117 10953 29173
rect 11009 29117 11095 29173
rect 11151 29117 11237 29173
rect 11293 29117 11379 29173
rect 11435 29117 11521 29173
rect 11577 29117 11663 29173
rect 11719 29117 11805 29173
rect 11861 29117 11947 29173
rect 12003 29117 12089 29173
rect 12145 29117 12231 29173
rect 12287 29117 12373 29173
rect 12429 29117 12515 29173
rect 12571 29117 12657 29173
rect 12713 29117 12799 29173
rect 12855 29117 12941 29173
rect 12997 29117 13083 29173
rect 13139 29117 13225 29173
rect 13281 29117 13367 29173
rect 13423 29117 13509 29173
rect 13565 29117 13651 29173
rect 13707 29117 13793 29173
rect 13849 29117 13935 29173
rect 13991 29117 14077 29173
rect 14133 29117 14219 29173
rect 14275 29117 14361 29173
rect 14417 29117 14503 29173
rect 14559 29117 14645 29173
rect 14701 29117 14787 29173
rect 14843 29117 15000 29173
rect 0 29031 15000 29117
rect 0 28975 161 29031
rect 217 28975 303 29031
rect 359 28975 445 29031
rect 501 28975 587 29031
rect 643 28975 729 29031
rect 785 28975 871 29031
rect 927 28975 1013 29031
rect 1069 28975 1155 29031
rect 1211 28975 1297 29031
rect 1353 28975 1439 29031
rect 1495 28975 1581 29031
rect 1637 28975 1723 29031
rect 1779 28975 1865 29031
rect 1921 28975 2007 29031
rect 2063 28975 2149 29031
rect 2205 28975 2291 29031
rect 2347 28975 2433 29031
rect 2489 28975 2575 29031
rect 2631 28975 2717 29031
rect 2773 28975 2859 29031
rect 2915 28975 3001 29031
rect 3057 28975 3143 29031
rect 3199 28975 3285 29031
rect 3341 28975 3427 29031
rect 3483 28975 3569 29031
rect 3625 28975 3711 29031
rect 3767 28975 3853 29031
rect 3909 28975 3995 29031
rect 4051 28975 4137 29031
rect 4193 28975 4279 29031
rect 4335 28975 4421 29031
rect 4477 28975 4563 29031
rect 4619 28975 4705 29031
rect 4761 28975 4847 29031
rect 4903 28975 4989 29031
rect 5045 28975 5131 29031
rect 5187 28975 5273 29031
rect 5329 28975 5415 29031
rect 5471 28975 5557 29031
rect 5613 28975 5699 29031
rect 5755 28975 5841 29031
rect 5897 28975 5983 29031
rect 6039 28975 6125 29031
rect 6181 28975 6267 29031
rect 6323 28975 6409 29031
rect 6465 28975 6551 29031
rect 6607 28975 6693 29031
rect 6749 28975 6835 29031
rect 6891 28975 6977 29031
rect 7033 28975 7119 29031
rect 7175 28975 7261 29031
rect 7317 28975 7403 29031
rect 7459 28975 7545 29031
rect 7601 28975 7687 29031
rect 7743 28975 7829 29031
rect 7885 28975 7971 29031
rect 8027 28975 8113 29031
rect 8169 28975 8255 29031
rect 8311 28975 8397 29031
rect 8453 28975 8539 29031
rect 8595 28975 8681 29031
rect 8737 28975 8823 29031
rect 8879 28975 8965 29031
rect 9021 28975 9107 29031
rect 9163 28975 9249 29031
rect 9305 28975 9391 29031
rect 9447 28975 9533 29031
rect 9589 28975 9675 29031
rect 9731 28975 9817 29031
rect 9873 28975 9959 29031
rect 10015 28975 10101 29031
rect 10157 28975 10243 29031
rect 10299 28975 10385 29031
rect 10441 28975 10527 29031
rect 10583 28975 10669 29031
rect 10725 28975 10811 29031
rect 10867 28975 10953 29031
rect 11009 28975 11095 29031
rect 11151 28975 11237 29031
rect 11293 28975 11379 29031
rect 11435 28975 11521 29031
rect 11577 28975 11663 29031
rect 11719 28975 11805 29031
rect 11861 28975 11947 29031
rect 12003 28975 12089 29031
rect 12145 28975 12231 29031
rect 12287 28975 12373 29031
rect 12429 28975 12515 29031
rect 12571 28975 12657 29031
rect 12713 28975 12799 29031
rect 12855 28975 12941 29031
rect 12997 28975 13083 29031
rect 13139 28975 13225 29031
rect 13281 28975 13367 29031
rect 13423 28975 13509 29031
rect 13565 28975 13651 29031
rect 13707 28975 13793 29031
rect 13849 28975 13935 29031
rect 13991 28975 14077 29031
rect 14133 28975 14219 29031
rect 14275 28975 14361 29031
rect 14417 28975 14503 29031
rect 14559 28975 14645 29031
rect 14701 28975 14787 29031
rect 14843 28975 15000 29031
rect 0 28889 15000 28975
rect 0 28833 161 28889
rect 217 28833 303 28889
rect 359 28833 445 28889
rect 501 28833 587 28889
rect 643 28833 729 28889
rect 785 28833 871 28889
rect 927 28833 1013 28889
rect 1069 28833 1155 28889
rect 1211 28833 1297 28889
rect 1353 28833 1439 28889
rect 1495 28833 1581 28889
rect 1637 28833 1723 28889
rect 1779 28833 1865 28889
rect 1921 28833 2007 28889
rect 2063 28833 2149 28889
rect 2205 28833 2291 28889
rect 2347 28833 2433 28889
rect 2489 28833 2575 28889
rect 2631 28833 2717 28889
rect 2773 28833 2859 28889
rect 2915 28833 3001 28889
rect 3057 28833 3143 28889
rect 3199 28833 3285 28889
rect 3341 28833 3427 28889
rect 3483 28833 3569 28889
rect 3625 28833 3711 28889
rect 3767 28833 3853 28889
rect 3909 28833 3995 28889
rect 4051 28833 4137 28889
rect 4193 28833 4279 28889
rect 4335 28833 4421 28889
rect 4477 28833 4563 28889
rect 4619 28833 4705 28889
rect 4761 28833 4847 28889
rect 4903 28833 4989 28889
rect 5045 28833 5131 28889
rect 5187 28833 5273 28889
rect 5329 28833 5415 28889
rect 5471 28833 5557 28889
rect 5613 28833 5699 28889
rect 5755 28833 5841 28889
rect 5897 28833 5983 28889
rect 6039 28833 6125 28889
rect 6181 28833 6267 28889
rect 6323 28833 6409 28889
rect 6465 28833 6551 28889
rect 6607 28833 6693 28889
rect 6749 28833 6835 28889
rect 6891 28833 6977 28889
rect 7033 28833 7119 28889
rect 7175 28833 7261 28889
rect 7317 28833 7403 28889
rect 7459 28833 7545 28889
rect 7601 28833 7687 28889
rect 7743 28833 7829 28889
rect 7885 28833 7971 28889
rect 8027 28833 8113 28889
rect 8169 28833 8255 28889
rect 8311 28833 8397 28889
rect 8453 28833 8539 28889
rect 8595 28833 8681 28889
rect 8737 28833 8823 28889
rect 8879 28833 8965 28889
rect 9021 28833 9107 28889
rect 9163 28833 9249 28889
rect 9305 28833 9391 28889
rect 9447 28833 9533 28889
rect 9589 28833 9675 28889
rect 9731 28833 9817 28889
rect 9873 28833 9959 28889
rect 10015 28833 10101 28889
rect 10157 28833 10243 28889
rect 10299 28833 10385 28889
rect 10441 28833 10527 28889
rect 10583 28833 10669 28889
rect 10725 28833 10811 28889
rect 10867 28833 10953 28889
rect 11009 28833 11095 28889
rect 11151 28833 11237 28889
rect 11293 28833 11379 28889
rect 11435 28833 11521 28889
rect 11577 28833 11663 28889
rect 11719 28833 11805 28889
rect 11861 28833 11947 28889
rect 12003 28833 12089 28889
rect 12145 28833 12231 28889
rect 12287 28833 12373 28889
rect 12429 28833 12515 28889
rect 12571 28833 12657 28889
rect 12713 28833 12799 28889
rect 12855 28833 12941 28889
rect 12997 28833 13083 28889
rect 13139 28833 13225 28889
rect 13281 28833 13367 28889
rect 13423 28833 13509 28889
rect 13565 28833 13651 28889
rect 13707 28833 13793 28889
rect 13849 28833 13935 28889
rect 13991 28833 14077 28889
rect 14133 28833 14219 28889
rect 14275 28833 14361 28889
rect 14417 28833 14503 28889
rect 14559 28833 14645 28889
rect 14701 28833 14787 28889
rect 14843 28833 15000 28889
rect 0 28747 15000 28833
rect 0 28691 161 28747
rect 217 28691 303 28747
rect 359 28691 445 28747
rect 501 28691 587 28747
rect 643 28691 729 28747
rect 785 28691 871 28747
rect 927 28691 1013 28747
rect 1069 28691 1155 28747
rect 1211 28691 1297 28747
rect 1353 28691 1439 28747
rect 1495 28691 1581 28747
rect 1637 28691 1723 28747
rect 1779 28691 1865 28747
rect 1921 28691 2007 28747
rect 2063 28691 2149 28747
rect 2205 28691 2291 28747
rect 2347 28691 2433 28747
rect 2489 28691 2575 28747
rect 2631 28691 2717 28747
rect 2773 28691 2859 28747
rect 2915 28691 3001 28747
rect 3057 28691 3143 28747
rect 3199 28691 3285 28747
rect 3341 28691 3427 28747
rect 3483 28691 3569 28747
rect 3625 28691 3711 28747
rect 3767 28691 3853 28747
rect 3909 28691 3995 28747
rect 4051 28691 4137 28747
rect 4193 28691 4279 28747
rect 4335 28691 4421 28747
rect 4477 28691 4563 28747
rect 4619 28691 4705 28747
rect 4761 28691 4847 28747
rect 4903 28691 4989 28747
rect 5045 28691 5131 28747
rect 5187 28691 5273 28747
rect 5329 28691 5415 28747
rect 5471 28691 5557 28747
rect 5613 28691 5699 28747
rect 5755 28691 5841 28747
rect 5897 28691 5983 28747
rect 6039 28691 6125 28747
rect 6181 28691 6267 28747
rect 6323 28691 6409 28747
rect 6465 28691 6551 28747
rect 6607 28691 6693 28747
rect 6749 28691 6835 28747
rect 6891 28691 6977 28747
rect 7033 28691 7119 28747
rect 7175 28691 7261 28747
rect 7317 28691 7403 28747
rect 7459 28691 7545 28747
rect 7601 28691 7687 28747
rect 7743 28691 7829 28747
rect 7885 28691 7971 28747
rect 8027 28691 8113 28747
rect 8169 28691 8255 28747
rect 8311 28691 8397 28747
rect 8453 28691 8539 28747
rect 8595 28691 8681 28747
rect 8737 28691 8823 28747
rect 8879 28691 8965 28747
rect 9021 28691 9107 28747
rect 9163 28691 9249 28747
rect 9305 28691 9391 28747
rect 9447 28691 9533 28747
rect 9589 28691 9675 28747
rect 9731 28691 9817 28747
rect 9873 28691 9959 28747
rect 10015 28691 10101 28747
rect 10157 28691 10243 28747
rect 10299 28691 10385 28747
rect 10441 28691 10527 28747
rect 10583 28691 10669 28747
rect 10725 28691 10811 28747
rect 10867 28691 10953 28747
rect 11009 28691 11095 28747
rect 11151 28691 11237 28747
rect 11293 28691 11379 28747
rect 11435 28691 11521 28747
rect 11577 28691 11663 28747
rect 11719 28691 11805 28747
rect 11861 28691 11947 28747
rect 12003 28691 12089 28747
rect 12145 28691 12231 28747
rect 12287 28691 12373 28747
rect 12429 28691 12515 28747
rect 12571 28691 12657 28747
rect 12713 28691 12799 28747
rect 12855 28691 12941 28747
rect 12997 28691 13083 28747
rect 13139 28691 13225 28747
rect 13281 28691 13367 28747
rect 13423 28691 13509 28747
rect 13565 28691 13651 28747
rect 13707 28691 13793 28747
rect 13849 28691 13935 28747
rect 13991 28691 14077 28747
rect 14133 28691 14219 28747
rect 14275 28691 14361 28747
rect 14417 28691 14503 28747
rect 14559 28691 14645 28747
rect 14701 28691 14787 28747
rect 14843 28691 15000 28747
rect 0 28605 15000 28691
rect 0 28549 161 28605
rect 217 28549 303 28605
rect 359 28549 445 28605
rect 501 28549 587 28605
rect 643 28549 729 28605
rect 785 28549 871 28605
rect 927 28549 1013 28605
rect 1069 28549 1155 28605
rect 1211 28549 1297 28605
rect 1353 28549 1439 28605
rect 1495 28549 1581 28605
rect 1637 28549 1723 28605
rect 1779 28549 1865 28605
rect 1921 28549 2007 28605
rect 2063 28549 2149 28605
rect 2205 28549 2291 28605
rect 2347 28549 2433 28605
rect 2489 28549 2575 28605
rect 2631 28549 2717 28605
rect 2773 28549 2859 28605
rect 2915 28549 3001 28605
rect 3057 28549 3143 28605
rect 3199 28549 3285 28605
rect 3341 28549 3427 28605
rect 3483 28549 3569 28605
rect 3625 28549 3711 28605
rect 3767 28549 3853 28605
rect 3909 28549 3995 28605
rect 4051 28549 4137 28605
rect 4193 28549 4279 28605
rect 4335 28549 4421 28605
rect 4477 28549 4563 28605
rect 4619 28549 4705 28605
rect 4761 28549 4847 28605
rect 4903 28549 4989 28605
rect 5045 28549 5131 28605
rect 5187 28549 5273 28605
rect 5329 28549 5415 28605
rect 5471 28549 5557 28605
rect 5613 28549 5699 28605
rect 5755 28549 5841 28605
rect 5897 28549 5983 28605
rect 6039 28549 6125 28605
rect 6181 28549 6267 28605
rect 6323 28549 6409 28605
rect 6465 28549 6551 28605
rect 6607 28549 6693 28605
rect 6749 28549 6835 28605
rect 6891 28549 6977 28605
rect 7033 28549 7119 28605
rect 7175 28549 7261 28605
rect 7317 28549 7403 28605
rect 7459 28549 7545 28605
rect 7601 28549 7687 28605
rect 7743 28549 7829 28605
rect 7885 28549 7971 28605
rect 8027 28549 8113 28605
rect 8169 28549 8255 28605
rect 8311 28549 8397 28605
rect 8453 28549 8539 28605
rect 8595 28549 8681 28605
rect 8737 28549 8823 28605
rect 8879 28549 8965 28605
rect 9021 28549 9107 28605
rect 9163 28549 9249 28605
rect 9305 28549 9391 28605
rect 9447 28549 9533 28605
rect 9589 28549 9675 28605
rect 9731 28549 9817 28605
rect 9873 28549 9959 28605
rect 10015 28549 10101 28605
rect 10157 28549 10243 28605
rect 10299 28549 10385 28605
rect 10441 28549 10527 28605
rect 10583 28549 10669 28605
rect 10725 28549 10811 28605
rect 10867 28549 10953 28605
rect 11009 28549 11095 28605
rect 11151 28549 11237 28605
rect 11293 28549 11379 28605
rect 11435 28549 11521 28605
rect 11577 28549 11663 28605
rect 11719 28549 11805 28605
rect 11861 28549 11947 28605
rect 12003 28549 12089 28605
rect 12145 28549 12231 28605
rect 12287 28549 12373 28605
rect 12429 28549 12515 28605
rect 12571 28549 12657 28605
rect 12713 28549 12799 28605
rect 12855 28549 12941 28605
rect 12997 28549 13083 28605
rect 13139 28549 13225 28605
rect 13281 28549 13367 28605
rect 13423 28549 13509 28605
rect 13565 28549 13651 28605
rect 13707 28549 13793 28605
rect 13849 28549 13935 28605
rect 13991 28549 14077 28605
rect 14133 28549 14219 28605
rect 14275 28549 14361 28605
rect 14417 28549 14503 28605
rect 14559 28549 14645 28605
rect 14701 28549 14787 28605
rect 14843 28549 15000 28605
rect 0 28463 15000 28549
rect 0 28407 161 28463
rect 217 28407 303 28463
rect 359 28407 445 28463
rect 501 28407 587 28463
rect 643 28407 729 28463
rect 785 28407 871 28463
rect 927 28407 1013 28463
rect 1069 28407 1155 28463
rect 1211 28407 1297 28463
rect 1353 28407 1439 28463
rect 1495 28407 1581 28463
rect 1637 28407 1723 28463
rect 1779 28407 1865 28463
rect 1921 28407 2007 28463
rect 2063 28407 2149 28463
rect 2205 28407 2291 28463
rect 2347 28407 2433 28463
rect 2489 28407 2575 28463
rect 2631 28407 2717 28463
rect 2773 28407 2859 28463
rect 2915 28407 3001 28463
rect 3057 28407 3143 28463
rect 3199 28407 3285 28463
rect 3341 28407 3427 28463
rect 3483 28407 3569 28463
rect 3625 28407 3711 28463
rect 3767 28407 3853 28463
rect 3909 28407 3995 28463
rect 4051 28407 4137 28463
rect 4193 28407 4279 28463
rect 4335 28407 4421 28463
rect 4477 28407 4563 28463
rect 4619 28407 4705 28463
rect 4761 28407 4847 28463
rect 4903 28407 4989 28463
rect 5045 28407 5131 28463
rect 5187 28407 5273 28463
rect 5329 28407 5415 28463
rect 5471 28407 5557 28463
rect 5613 28407 5699 28463
rect 5755 28407 5841 28463
rect 5897 28407 5983 28463
rect 6039 28407 6125 28463
rect 6181 28407 6267 28463
rect 6323 28407 6409 28463
rect 6465 28407 6551 28463
rect 6607 28407 6693 28463
rect 6749 28407 6835 28463
rect 6891 28407 6977 28463
rect 7033 28407 7119 28463
rect 7175 28407 7261 28463
rect 7317 28407 7403 28463
rect 7459 28407 7545 28463
rect 7601 28407 7687 28463
rect 7743 28407 7829 28463
rect 7885 28407 7971 28463
rect 8027 28407 8113 28463
rect 8169 28407 8255 28463
rect 8311 28407 8397 28463
rect 8453 28407 8539 28463
rect 8595 28407 8681 28463
rect 8737 28407 8823 28463
rect 8879 28407 8965 28463
rect 9021 28407 9107 28463
rect 9163 28407 9249 28463
rect 9305 28407 9391 28463
rect 9447 28407 9533 28463
rect 9589 28407 9675 28463
rect 9731 28407 9817 28463
rect 9873 28407 9959 28463
rect 10015 28407 10101 28463
rect 10157 28407 10243 28463
rect 10299 28407 10385 28463
rect 10441 28407 10527 28463
rect 10583 28407 10669 28463
rect 10725 28407 10811 28463
rect 10867 28407 10953 28463
rect 11009 28407 11095 28463
rect 11151 28407 11237 28463
rect 11293 28407 11379 28463
rect 11435 28407 11521 28463
rect 11577 28407 11663 28463
rect 11719 28407 11805 28463
rect 11861 28407 11947 28463
rect 12003 28407 12089 28463
rect 12145 28407 12231 28463
rect 12287 28407 12373 28463
rect 12429 28407 12515 28463
rect 12571 28407 12657 28463
rect 12713 28407 12799 28463
rect 12855 28407 12941 28463
rect 12997 28407 13083 28463
rect 13139 28407 13225 28463
rect 13281 28407 13367 28463
rect 13423 28407 13509 28463
rect 13565 28407 13651 28463
rect 13707 28407 13793 28463
rect 13849 28407 13935 28463
rect 13991 28407 14077 28463
rect 14133 28407 14219 28463
rect 14275 28407 14361 28463
rect 14417 28407 14503 28463
rect 14559 28407 14645 28463
rect 14701 28407 14787 28463
rect 14843 28407 15000 28463
rect 0 28321 15000 28407
rect 0 28265 161 28321
rect 217 28265 303 28321
rect 359 28265 445 28321
rect 501 28265 587 28321
rect 643 28265 729 28321
rect 785 28265 871 28321
rect 927 28265 1013 28321
rect 1069 28265 1155 28321
rect 1211 28265 1297 28321
rect 1353 28265 1439 28321
rect 1495 28265 1581 28321
rect 1637 28265 1723 28321
rect 1779 28265 1865 28321
rect 1921 28265 2007 28321
rect 2063 28265 2149 28321
rect 2205 28265 2291 28321
rect 2347 28265 2433 28321
rect 2489 28265 2575 28321
rect 2631 28265 2717 28321
rect 2773 28265 2859 28321
rect 2915 28265 3001 28321
rect 3057 28265 3143 28321
rect 3199 28265 3285 28321
rect 3341 28265 3427 28321
rect 3483 28265 3569 28321
rect 3625 28265 3711 28321
rect 3767 28265 3853 28321
rect 3909 28265 3995 28321
rect 4051 28265 4137 28321
rect 4193 28265 4279 28321
rect 4335 28265 4421 28321
rect 4477 28265 4563 28321
rect 4619 28265 4705 28321
rect 4761 28265 4847 28321
rect 4903 28265 4989 28321
rect 5045 28265 5131 28321
rect 5187 28265 5273 28321
rect 5329 28265 5415 28321
rect 5471 28265 5557 28321
rect 5613 28265 5699 28321
rect 5755 28265 5841 28321
rect 5897 28265 5983 28321
rect 6039 28265 6125 28321
rect 6181 28265 6267 28321
rect 6323 28265 6409 28321
rect 6465 28265 6551 28321
rect 6607 28265 6693 28321
rect 6749 28265 6835 28321
rect 6891 28265 6977 28321
rect 7033 28265 7119 28321
rect 7175 28265 7261 28321
rect 7317 28265 7403 28321
rect 7459 28265 7545 28321
rect 7601 28265 7687 28321
rect 7743 28265 7829 28321
rect 7885 28265 7971 28321
rect 8027 28265 8113 28321
rect 8169 28265 8255 28321
rect 8311 28265 8397 28321
rect 8453 28265 8539 28321
rect 8595 28265 8681 28321
rect 8737 28265 8823 28321
rect 8879 28265 8965 28321
rect 9021 28265 9107 28321
rect 9163 28265 9249 28321
rect 9305 28265 9391 28321
rect 9447 28265 9533 28321
rect 9589 28265 9675 28321
rect 9731 28265 9817 28321
rect 9873 28265 9959 28321
rect 10015 28265 10101 28321
rect 10157 28265 10243 28321
rect 10299 28265 10385 28321
rect 10441 28265 10527 28321
rect 10583 28265 10669 28321
rect 10725 28265 10811 28321
rect 10867 28265 10953 28321
rect 11009 28265 11095 28321
rect 11151 28265 11237 28321
rect 11293 28265 11379 28321
rect 11435 28265 11521 28321
rect 11577 28265 11663 28321
rect 11719 28265 11805 28321
rect 11861 28265 11947 28321
rect 12003 28265 12089 28321
rect 12145 28265 12231 28321
rect 12287 28265 12373 28321
rect 12429 28265 12515 28321
rect 12571 28265 12657 28321
rect 12713 28265 12799 28321
rect 12855 28265 12941 28321
rect 12997 28265 13083 28321
rect 13139 28265 13225 28321
rect 13281 28265 13367 28321
rect 13423 28265 13509 28321
rect 13565 28265 13651 28321
rect 13707 28265 13793 28321
rect 13849 28265 13935 28321
rect 13991 28265 14077 28321
rect 14133 28265 14219 28321
rect 14275 28265 14361 28321
rect 14417 28265 14503 28321
rect 14559 28265 14645 28321
rect 14701 28265 14787 28321
rect 14843 28265 15000 28321
rect 0 28179 15000 28265
rect 0 28123 161 28179
rect 217 28123 303 28179
rect 359 28123 445 28179
rect 501 28123 587 28179
rect 643 28123 729 28179
rect 785 28123 871 28179
rect 927 28123 1013 28179
rect 1069 28123 1155 28179
rect 1211 28123 1297 28179
rect 1353 28123 1439 28179
rect 1495 28123 1581 28179
rect 1637 28123 1723 28179
rect 1779 28123 1865 28179
rect 1921 28123 2007 28179
rect 2063 28123 2149 28179
rect 2205 28123 2291 28179
rect 2347 28123 2433 28179
rect 2489 28123 2575 28179
rect 2631 28123 2717 28179
rect 2773 28123 2859 28179
rect 2915 28123 3001 28179
rect 3057 28123 3143 28179
rect 3199 28123 3285 28179
rect 3341 28123 3427 28179
rect 3483 28123 3569 28179
rect 3625 28123 3711 28179
rect 3767 28123 3853 28179
rect 3909 28123 3995 28179
rect 4051 28123 4137 28179
rect 4193 28123 4279 28179
rect 4335 28123 4421 28179
rect 4477 28123 4563 28179
rect 4619 28123 4705 28179
rect 4761 28123 4847 28179
rect 4903 28123 4989 28179
rect 5045 28123 5131 28179
rect 5187 28123 5273 28179
rect 5329 28123 5415 28179
rect 5471 28123 5557 28179
rect 5613 28123 5699 28179
rect 5755 28123 5841 28179
rect 5897 28123 5983 28179
rect 6039 28123 6125 28179
rect 6181 28123 6267 28179
rect 6323 28123 6409 28179
rect 6465 28123 6551 28179
rect 6607 28123 6693 28179
rect 6749 28123 6835 28179
rect 6891 28123 6977 28179
rect 7033 28123 7119 28179
rect 7175 28123 7261 28179
rect 7317 28123 7403 28179
rect 7459 28123 7545 28179
rect 7601 28123 7687 28179
rect 7743 28123 7829 28179
rect 7885 28123 7971 28179
rect 8027 28123 8113 28179
rect 8169 28123 8255 28179
rect 8311 28123 8397 28179
rect 8453 28123 8539 28179
rect 8595 28123 8681 28179
rect 8737 28123 8823 28179
rect 8879 28123 8965 28179
rect 9021 28123 9107 28179
rect 9163 28123 9249 28179
rect 9305 28123 9391 28179
rect 9447 28123 9533 28179
rect 9589 28123 9675 28179
rect 9731 28123 9817 28179
rect 9873 28123 9959 28179
rect 10015 28123 10101 28179
rect 10157 28123 10243 28179
rect 10299 28123 10385 28179
rect 10441 28123 10527 28179
rect 10583 28123 10669 28179
rect 10725 28123 10811 28179
rect 10867 28123 10953 28179
rect 11009 28123 11095 28179
rect 11151 28123 11237 28179
rect 11293 28123 11379 28179
rect 11435 28123 11521 28179
rect 11577 28123 11663 28179
rect 11719 28123 11805 28179
rect 11861 28123 11947 28179
rect 12003 28123 12089 28179
rect 12145 28123 12231 28179
rect 12287 28123 12373 28179
rect 12429 28123 12515 28179
rect 12571 28123 12657 28179
rect 12713 28123 12799 28179
rect 12855 28123 12941 28179
rect 12997 28123 13083 28179
rect 13139 28123 13225 28179
rect 13281 28123 13367 28179
rect 13423 28123 13509 28179
rect 13565 28123 13651 28179
rect 13707 28123 13793 28179
rect 13849 28123 13935 28179
rect 13991 28123 14077 28179
rect 14133 28123 14219 28179
rect 14275 28123 14361 28179
rect 14417 28123 14503 28179
rect 14559 28123 14645 28179
rect 14701 28123 14787 28179
rect 14843 28123 15000 28179
rect 0 28037 15000 28123
rect 0 27981 161 28037
rect 217 27981 303 28037
rect 359 27981 445 28037
rect 501 27981 587 28037
rect 643 27981 729 28037
rect 785 27981 871 28037
rect 927 27981 1013 28037
rect 1069 27981 1155 28037
rect 1211 27981 1297 28037
rect 1353 27981 1439 28037
rect 1495 27981 1581 28037
rect 1637 27981 1723 28037
rect 1779 27981 1865 28037
rect 1921 27981 2007 28037
rect 2063 27981 2149 28037
rect 2205 27981 2291 28037
rect 2347 27981 2433 28037
rect 2489 27981 2575 28037
rect 2631 27981 2717 28037
rect 2773 27981 2859 28037
rect 2915 27981 3001 28037
rect 3057 27981 3143 28037
rect 3199 27981 3285 28037
rect 3341 27981 3427 28037
rect 3483 27981 3569 28037
rect 3625 27981 3711 28037
rect 3767 27981 3853 28037
rect 3909 27981 3995 28037
rect 4051 27981 4137 28037
rect 4193 27981 4279 28037
rect 4335 27981 4421 28037
rect 4477 27981 4563 28037
rect 4619 27981 4705 28037
rect 4761 27981 4847 28037
rect 4903 27981 4989 28037
rect 5045 27981 5131 28037
rect 5187 27981 5273 28037
rect 5329 27981 5415 28037
rect 5471 27981 5557 28037
rect 5613 27981 5699 28037
rect 5755 27981 5841 28037
rect 5897 27981 5983 28037
rect 6039 27981 6125 28037
rect 6181 27981 6267 28037
rect 6323 27981 6409 28037
rect 6465 27981 6551 28037
rect 6607 27981 6693 28037
rect 6749 27981 6835 28037
rect 6891 27981 6977 28037
rect 7033 27981 7119 28037
rect 7175 27981 7261 28037
rect 7317 27981 7403 28037
rect 7459 27981 7545 28037
rect 7601 27981 7687 28037
rect 7743 27981 7829 28037
rect 7885 27981 7971 28037
rect 8027 27981 8113 28037
rect 8169 27981 8255 28037
rect 8311 27981 8397 28037
rect 8453 27981 8539 28037
rect 8595 27981 8681 28037
rect 8737 27981 8823 28037
rect 8879 27981 8965 28037
rect 9021 27981 9107 28037
rect 9163 27981 9249 28037
rect 9305 27981 9391 28037
rect 9447 27981 9533 28037
rect 9589 27981 9675 28037
rect 9731 27981 9817 28037
rect 9873 27981 9959 28037
rect 10015 27981 10101 28037
rect 10157 27981 10243 28037
rect 10299 27981 10385 28037
rect 10441 27981 10527 28037
rect 10583 27981 10669 28037
rect 10725 27981 10811 28037
rect 10867 27981 10953 28037
rect 11009 27981 11095 28037
rect 11151 27981 11237 28037
rect 11293 27981 11379 28037
rect 11435 27981 11521 28037
rect 11577 27981 11663 28037
rect 11719 27981 11805 28037
rect 11861 27981 11947 28037
rect 12003 27981 12089 28037
rect 12145 27981 12231 28037
rect 12287 27981 12373 28037
rect 12429 27981 12515 28037
rect 12571 27981 12657 28037
rect 12713 27981 12799 28037
rect 12855 27981 12941 28037
rect 12997 27981 13083 28037
rect 13139 27981 13225 28037
rect 13281 27981 13367 28037
rect 13423 27981 13509 28037
rect 13565 27981 13651 28037
rect 13707 27981 13793 28037
rect 13849 27981 13935 28037
rect 13991 27981 14077 28037
rect 14133 27981 14219 28037
rect 14275 27981 14361 28037
rect 14417 27981 14503 28037
rect 14559 27981 14645 28037
rect 14701 27981 14787 28037
rect 14843 27981 15000 28037
rect 0 27895 15000 27981
rect 0 27839 161 27895
rect 217 27839 303 27895
rect 359 27839 445 27895
rect 501 27839 587 27895
rect 643 27839 729 27895
rect 785 27839 871 27895
rect 927 27839 1013 27895
rect 1069 27839 1155 27895
rect 1211 27839 1297 27895
rect 1353 27839 1439 27895
rect 1495 27839 1581 27895
rect 1637 27839 1723 27895
rect 1779 27839 1865 27895
rect 1921 27839 2007 27895
rect 2063 27839 2149 27895
rect 2205 27839 2291 27895
rect 2347 27839 2433 27895
rect 2489 27839 2575 27895
rect 2631 27839 2717 27895
rect 2773 27839 2859 27895
rect 2915 27839 3001 27895
rect 3057 27839 3143 27895
rect 3199 27839 3285 27895
rect 3341 27839 3427 27895
rect 3483 27839 3569 27895
rect 3625 27839 3711 27895
rect 3767 27839 3853 27895
rect 3909 27839 3995 27895
rect 4051 27839 4137 27895
rect 4193 27839 4279 27895
rect 4335 27839 4421 27895
rect 4477 27839 4563 27895
rect 4619 27839 4705 27895
rect 4761 27839 4847 27895
rect 4903 27839 4989 27895
rect 5045 27839 5131 27895
rect 5187 27839 5273 27895
rect 5329 27839 5415 27895
rect 5471 27839 5557 27895
rect 5613 27839 5699 27895
rect 5755 27839 5841 27895
rect 5897 27839 5983 27895
rect 6039 27839 6125 27895
rect 6181 27839 6267 27895
rect 6323 27839 6409 27895
rect 6465 27839 6551 27895
rect 6607 27839 6693 27895
rect 6749 27839 6835 27895
rect 6891 27839 6977 27895
rect 7033 27839 7119 27895
rect 7175 27839 7261 27895
rect 7317 27839 7403 27895
rect 7459 27839 7545 27895
rect 7601 27839 7687 27895
rect 7743 27839 7829 27895
rect 7885 27839 7971 27895
rect 8027 27839 8113 27895
rect 8169 27839 8255 27895
rect 8311 27839 8397 27895
rect 8453 27839 8539 27895
rect 8595 27839 8681 27895
rect 8737 27839 8823 27895
rect 8879 27839 8965 27895
rect 9021 27839 9107 27895
rect 9163 27839 9249 27895
rect 9305 27839 9391 27895
rect 9447 27839 9533 27895
rect 9589 27839 9675 27895
rect 9731 27839 9817 27895
rect 9873 27839 9959 27895
rect 10015 27839 10101 27895
rect 10157 27839 10243 27895
rect 10299 27839 10385 27895
rect 10441 27839 10527 27895
rect 10583 27839 10669 27895
rect 10725 27839 10811 27895
rect 10867 27839 10953 27895
rect 11009 27839 11095 27895
rect 11151 27839 11237 27895
rect 11293 27839 11379 27895
rect 11435 27839 11521 27895
rect 11577 27839 11663 27895
rect 11719 27839 11805 27895
rect 11861 27839 11947 27895
rect 12003 27839 12089 27895
rect 12145 27839 12231 27895
rect 12287 27839 12373 27895
rect 12429 27839 12515 27895
rect 12571 27839 12657 27895
rect 12713 27839 12799 27895
rect 12855 27839 12941 27895
rect 12997 27839 13083 27895
rect 13139 27839 13225 27895
rect 13281 27839 13367 27895
rect 13423 27839 13509 27895
rect 13565 27839 13651 27895
rect 13707 27839 13793 27895
rect 13849 27839 13935 27895
rect 13991 27839 14077 27895
rect 14133 27839 14219 27895
rect 14275 27839 14361 27895
rect 14417 27839 14503 27895
rect 14559 27839 14645 27895
rect 14701 27839 14787 27895
rect 14843 27839 15000 27895
rect 0 27753 15000 27839
rect 0 27697 161 27753
rect 217 27697 303 27753
rect 359 27697 445 27753
rect 501 27697 587 27753
rect 643 27697 729 27753
rect 785 27697 871 27753
rect 927 27697 1013 27753
rect 1069 27697 1155 27753
rect 1211 27697 1297 27753
rect 1353 27697 1439 27753
rect 1495 27697 1581 27753
rect 1637 27697 1723 27753
rect 1779 27697 1865 27753
rect 1921 27697 2007 27753
rect 2063 27697 2149 27753
rect 2205 27697 2291 27753
rect 2347 27697 2433 27753
rect 2489 27697 2575 27753
rect 2631 27697 2717 27753
rect 2773 27697 2859 27753
rect 2915 27697 3001 27753
rect 3057 27697 3143 27753
rect 3199 27697 3285 27753
rect 3341 27697 3427 27753
rect 3483 27697 3569 27753
rect 3625 27697 3711 27753
rect 3767 27697 3853 27753
rect 3909 27697 3995 27753
rect 4051 27697 4137 27753
rect 4193 27697 4279 27753
rect 4335 27697 4421 27753
rect 4477 27697 4563 27753
rect 4619 27697 4705 27753
rect 4761 27697 4847 27753
rect 4903 27697 4989 27753
rect 5045 27697 5131 27753
rect 5187 27697 5273 27753
rect 5329 27697 5415 27753
rect 5471 27697 5557 27753
rect 5613 27697 5699 27753
rect 5755 27697 5841 27753
rect 5897 27697 5983 27753
rect 6039 27697 6125 27753
rect 6181 27697 6267 27753
rect 6323 27697 6409 27753
rect 6465 27697 6551 27753
rect 6607 27697 6693 27753
rect 6749 27697 6835 27753
rect 6891 27697 6977 27753
rect 7033 27697 7119 27753
rect 7175 27697 7261 27753
rect 7317 27697 7403 27753
rect 7459 27697 7545 27753
rect 7601 27697 7687 27753
rect 7743 27697 7829 27753
rect 7885 27697 7971 27753
rect 8027 27697 8113 27753
rect 8169 27697 8255 27753
rect 8311 27697 8397 27753
rect 8453 27697 8539 27753
rect 8595 27697 8681 27753
rect 8737 27697 8823 27753
rect 8879 27697 8965 27753
rect 9021 27697 9107 27753
rect 9163 27697 9249 27753
rect 9305 27697 9391 27753
rect 9447 27697 9533 27753
rect 9589 27697 9675 27753
rect 9731 27697 9817 27753
rect 9873 27697 9959 27753
rect 10015 27697 10101 27753
rect 10157 27697 10243 27753
rect 10299 27697 10385 27753
rect 10441 27697 10527 27753
rect 10583 27697 10669 27753
rect 10725 27697 10811 27753
rect 10867 27697 10953 27753
rect 11009 27697 11095 27753
rect 11151 27697 11237 27753
rect 11293 27697 11379 27753
rect 11435 27697 11521 27753
rect 11577 27697 11663 27753
rect 11719 27697 11805 27753
rect 11861 27697 11947 27753
rect 12003 27697 12089 27753
rect 12145 27697 12231 27753
rect 12287 27697 12373 27753
rect 12429 27697 12515 27753
rect 12571 27697 12657 27753
rect 12713 27697 12799 27753
rect 12855 27697 12941 27753
rect 12997 27697 13083 27753
rect 13139 27697 13225 27753
rect 13281 27697 13367 27753
rect 13423 27697 13509 27753
rect 13565 27697 13651 27753
rect 13707 27697 13793 27753
rect 13849 27697 13935 27753
rect 13991 27697 14077 27753
rect 14133 27697 14219 27753
rect 14275 27697 14361 27753
rect 14417 27697 14503 27753
rect 14559 27697 14645 27753
rect 14701 27697 14787 27753
rect 14843 27697 15000 27753
rect 0 27611 15000 27697
rect 0 27555 161 27611
rect 217 27555 303 27611
rect 359 27555 445 27611
rect 501 27555 587 27611
rect 643 27555 729 27611
rect 785 27555 871 27611
rect 927 27555 1013 27611
rect 1069 27555 1155 27611
rect 1211 27555 1297 27611
rect 1353 27555 1439 27611
rect 1495 27555 1581 27611
rect 1637 27555 1723 27611
rect 1779 27555 1865 27611
rect 1921 27555 2007 27611
rect 2063 27555 2149 27611
rect 2205 27555 2291 27611
rect 2347 27555 2433 27611
rect 2489 27555 2575 27611
rect 2631 27555 2717 27611
rect 2773 27555 2859 27611
rect 2915 27555 3001 27611
rect 3057 27555 3143 27611
rect 3199 27555 3285 27611
rect 3341 27555 3427 27611
rect 3483 27555 3569 27611
rect 3625 27555 3711 27611
rect 3767 27555 3853 27611
rect 3909 27555 3995 27611
rect 4051 27555 4137 27611
rect 4193 27555 4279 27611
rect 4335 27555 4421 27611
rect 4477 27555 4563 27611
rect 4619 27555 4705 27611
rect 4761 27555 4847 27611
rect 4903 27555 4989 27611
rect 5045 27555 5131 27611
rect 5187 27555 5273 27611
rect 5329 27555 5415 27611
rect 5471 27555 5557 27611
rect 5613 27555 5699 27611
rect 5755 27555 5841 27611
rect 5897 27555 5983 27611
rect 6039 27555 6125 27611
rect 6181 27555 6267 27611
rect 6323 27555 6409 27611
rect 6465 27555 6551 27611
rect 6607 27555 6693 27611
rect 6749 27555 6835 27611
rect 6891 27555 6977 27611
rect 7033 27555 7119 27611
rect 7175 27555 7261 27611
rect 7317 27555 7403 27611
rect 7459 27555 7545 27611
rect 7601 27555 7687 27611
rect 7743 27555 7829 27611
rect 7885 27555 7971 27611
rect 8027 27555 8113 27611
rect 8169 27555 8255 27611
rect 8311 27555 8397 27611
rect 8453 27555 8539 27611
rect 8595 27555 8681 27611
rect 8737 27555 8823 27611
rect 8879 27555 8965 27611
rect 9021 27555 9107 27611
rect 9163 27555 9249 27611
rect 9305 27555 9391 27611
rect 9447 27555 9533 27611
rect 9589 27555 9675 27611
rect 9731 27555 9817 27611
rect 9873 27555 9959 27611
rect 10015 27555 10101 27611
rect 10157 27555 10243 27611
rect 10299 27555 10385 27611
rect 10441 27555 10527 27611
rect 10583 27555 10669 27611
rect 10725 27555 10811 27611
rect 10867 27555 10953 27611
rect 11009 27555 11095 27611
rect 11151 27555 11237 27611
rect 11293 27555 11379 27611
rect 11435 27555 11521 27611
rect 11577 27555 11663 27611
rect 11719 27555 11805 27611
rect 11861 27555 11947 27611
rect 12003 27555 12089 27611
rect 12145 27555 12231 27611
rect 12287 27555 12373 27611
rect 12429 27555 12515 27611
rect 12571 27555 12657 27611
rect 12713 27555 12799 27611
rect 12855 27555 12941 27611
rect 12997 27555 13083 27611
rect 13139 27555 13225 27611
rect 13281 27555 13367 27611
rect 13423 27555 13509 27611
rect 13565 27555 13651 27611
rect 13707 27555 13793 27611
rect 13849 27555 13935 27611
rect 13991 27555 14077 27611
rect 14133 27555 14219 27611
rect 14275 27555 14361 27611
rect 14417 27555 14503 27611
rect 14559 27555 14645 27611
rect 14701 27555 14787 27611
rect 14843 27555 15000 27611
rect 0 27469 15000 27555
rect 0 27413 161 27469
rect 217 27413 303 27469
rect 359 27413 445 27469
rect 501 27413 587 27469
rect 643 27413 729 27469
rect 785 27413 871 27469
rect 927 27413 1013 27469
rect 1069 27413 1155 27469
rect 1211 27413 1297 27469
rect 1353 27413 1439 27469
rect 1495 27413 1581 27469
rect 1637 27413 1723 27469
rect 1779 27413 1865 27469
rect 1921 27413 2007 27469
rect 2063 27413 2149 27469
rect 2205 27413 2291 27469
rect 2347 27413 2433 27469
rect 2489 27413 2575 27469
rect 2631 27413 2717 27469
rect 2773 27413 2859 27469
rect 2915 27413 3001 27469
rect 3057 27413 3143 27469
rect 3199 27413 3285 27469
rect 3341 27413 3427 27469
rect 3483 27413 3569 27469
rect 3625 27413 3711 27469
rect 3767 27413 3853 27469
rect 3909 27413 3995 27469
rect 4051 27413 4137 27469
rect 4193 27413 4279 27469
rect 4335 27413 4421 27469
rect 4477 27413 4563 27469
rect 4619 27413 4705 27469
rect 4761 27413 4847 27469
rect 4903 27413 4989 27469
rect 5045 27413 5131 27469
rect 5187 27413 5273 27469
rect 5329 27413 5415 27469
rect 5471 27413 5557 27469
rect 5613 27413 5699 27469
rect 5755 27413 5841 27469
rect 5897 27413 5983 27469
rect 6039 27413 6125 27469
rect 6181 27413 6267 27469
rect 6323 27413 6409 27469
rect 6465 27413 6551 27469
rect 6607 27413 6693 27469
rect 6749 27413 6835 27469
rect 6891 27413 6977 27469
rect 7033 27413 7119 27469
rect 7175 27413 7261 27469
rect 7317 27413 7403 27469
rect 7459 27413 7545 27469
rect 7601 27413 7687 27469
rect 7743 27413 7829 27469
rect 7885 27413 7971 27469
rect 8027 27413 8113 27469
rect 8169 27413 8255 27469
rect 8311 27413 8397 27469
rect 8453 27413 8539 27469
rect 8595 27413 8681 27469
rect 8737 27413 8823 27469
rect 8879 27413 8965 27469
rect 9021 27413 9107 27469
rect 9163 27413 9249 27469
rect 9305 27413 9391 27469
rect 9447 27413 9533 27469
rect 9589 27413 9675 27469
rect 9731 27413 9817 27469
rect 9873 27413 9959 27469
rect 10015 27413 10101 27469
rect 10157 27413 10243 27469
rect 10299 27413 10385 27469
rect 10441 27413 10527 27469
rect 10583 27413 10669 27469
rect 10725 27413 10811 27469
rect 10867 27413 10953 27469
rect 11009 27413 11095 27469
rect 11151 27413 11237 27469
rect 11293 27413 11379 27469
rect 11435 27413 11521 27469
rect 11577 27413 11663 27469
rect 11719 27413 11805 27469
rect 11861 27413 11947 27469
rect 12003 27413 12089 27469
rect 12145 27413 12231 27469
rect 12287 27413 12373 27469
rect 12429 27413 12515 27469
rect 12571 27413 12657 27469
rect 12713 27413 12799 27469
rect 12855 27413 12941 27469
rect 12997 27413 13083 27469
rect 13139 27413 13225 27469
rect 13281 27413 13367 27469
rect 13423 27413 13509 27469
rect 13565 27413 13651 27469
rect 13707 27413 13793 27469
rect 13849 27413 13935 27469
rect 13991 27413 14077 27469
rect 14133 27413 14219 27469
rect 14275 27413 14361 27469
rect 14417 27413 14503 27469
rect 14559 27413 14645 27469
rect 14701 27413 14787 27469
rect 14843 27413 15000 27469
rect 0 27327 15000 27413
rect 0 27271 161 27327
rect 217 27271 303 27327
rect 359 27271 445 27327
rect 501 27271 587 27327
rect 643 27271 729 27327
rect 785 27271 871 27327
rect 927 27271 1013 27327
rect 1069 27271 1155 27327
rect 1211 27271 1297 27327
rect 1353 27271 1439 27327
rect 1495 27271 1581 27327
rect 1637 27271 1723 27327
rect 1779 27271 1865 27327
rect 1921 27271 2007 27327
rect 2063 27271 2149 27327
rect 2205 27271 2291 27327
rect 2347 27271 2433 27327
rect 2489 27271 2575 27327
rect 2631 27271 2717 27327
rect 2773 27271 2859 27327
rect 2915 27271 3001 27327
rect 3057 27271 3143 27327
rect 3199 27271 3285 27327
rect 3341 27271 3427 27327
rect 3483 27271 3569 27327
rect 3625 27271 3711 27327
rect 3767 27271 3853 27327
rect 3909 27271 3995 27327
rect 4051 27271 4137 27327
rect 4193 27271 4279 27327
rect 4335 27271 4421 27327
rect 4477 27271 4563 27327
rect 4619 27271 4705 27327
rect 4761 27271 4847 27327
rect 4903 27271 4989 27327
rect 5045 27271 5131 27327
rect 5187 27271 5273 27327
rect 5329 27271 5415 27327
rect 5471 27271 5557 27327
rect 5613 27271 5699 27327
rect 5755 27271 5841 27327
rect 5897 27271 5983 27327
rect 6039 27271 6125 27327
rect 6181 27271 6267 27327
rect 6323 27271 6409 27327
rect 6465 27271 6551 27327
rect 6607 27271 6693 27327
rect 6749 27271 6835 27327
rect 6891 27271 6977 27327
rect 7033 27271 7119 27327
rect 7175 27271 7261 27327
rect 7317 27271 7403 27327
rect 7459 27271 7545 27327
rect 7601 27271 7687 27327
rect 7743 27271 7829 27327
rect 7885 27271 7971 27327
rect 8027 27271 8113 27327
rect 8169 27271 8255 27327
rect 8311 27271 8397 27327
rect 8453 27271 8539 27327
rect 8595 27271 8681 27327
rect 8737 27271 8823 27327
rect 8879 27271 8965 27327
rect 9021 27271 9107 27327
rect 9163 27271 9249 27327
rect 9305 27271 9391 27327
rect 9447 27271 9533 27327
rect 9589 27271 9675 27327
rect 9731 27271 9817 27327
rect 9873 27271 9959 27327
rect 10015 27271 10101 27327
rect 10157 27271 10243 27327
rect 10299 27271 10385 27327
rect 10441 27271 10527 27327
rect 10583 27271 10669 27327
rect 10725 27271 10811 27327
rect 10867 27271 10953 27327
rect 11009 27271 11095 27327
rect 11151 27271 11237 27327
rect 11293 27271 11379 27327
rect 11435 27271 11521 27327
rect 11577 27271 11663 27327
rect 11719 27271 11805 27327
rect 11861 27271 11947 27327
rect 12003 27271 12089 27327
rect 12145 27271 12231 27327
rect 12287 27271 12373 27327
rect 12429 27271 12515 27327
rect 12571 27271 12657 27327
rect 12713 27271 12799 27327
rect 12855 27271 12941 27327
rect 12997 27271 13083 27327
rect 13139 27271 13225 27327
rect 13281 27271 13367 27327
rect 13423 27271 13509 27327
rect 13565 27271 13651 27327
rect 13707 27271 13793 27327
rect 13849 27271 13935 27327
rect 13991 27271 14077 27327
rect 14133 27271 14219 27327
rect 14275 27271 14361 27327
rect 14417 27271 14503 27327
rect 14559 27271 14645 27327
rect 14701 27271 14787 27327
rect 14843 27271 15000 27327
rect 0 27185 15000 27271
rect 0 27129 161 27185
rect 217 27129 303 27185
rect 359 27129 445 27185
rect 501 27129 587 27185
rect 643 27129 729 27185
rect 785 27129 871 27185
rect 927 27129 1013 27185
rect 1069 27129 1155 27185
rect 1211 27129 1297 27185
rect 1353 27129 1439 27185
rect 1495 27129 1581 27185
rect 1637 27129 1723 27185
rect 1779 27129 1865 27185
rect 1921 27129 2007 27185
rect 2063 27129 2149 27185
rect 2205 27129 2291 27185
rect 2347 27129 2433 27185
rect 2489 27129 2575 27185
rect 2631 27129 2717 27185
rect 2773 27129 2859 27185
rect 2915 27129 3001 27185
rect 3057 27129 3143 27185
rect 3199 27129 3285 27185
rect 3341 27129 3427 27185
rect 3483 27129 3569 27185
rect 3625 27129 3711 27185
rect 3767 27129 3853 27185
rect 3909 27129 3995 27185
rect 4051 27129 4137 27185
rect 4193 27129 4279 27185
rect 4335 27129 4421 27185
rect 4477 27129 4563 27185
rect 4619 27129 4705 27185
rect 4761 27129 4847 27185
rect 4903 27129 4989 27185
rect 5045 27129 5131 27185
rect 5187 27129 5273 27185
rect 5329 27129 5415 27185
rect 5471 27129 5557 27185
rect 5613 27129 5699 27185
rect 5755 27129 5841 27185
rect 5897 27129 5983 27185
rect 6039 27129 6125 27185
rect 6181 27129 6267 27185
rect 6323 27129 6409 27185
rect 6465 27129 6551 27185
rect 6607 27129 6693 27185
rect 6749 27129 6835 27185
rect 6891 27129 6977 27185
rect 7033 27129 7119 27185
rect 7175 27129 7261 27185
rect 7317 27129 7403 27185
rect 7459 27129 7545 27185
rect 7601 27129 7687 27185
rect 7743 27129 7829 27185
rect 7885 27129 7971 27185
rect 8027 27129 8113 27185
rect 8169 27129 8255 27185
rect 8311 27129 8397 27185
rect 8453 27129 8539 27185
rect 8595 27129 8681 27185
rect 8737 27129 8823 27185
rect 8879 27129 8965 27185
rect 9021 27129 9107 27185
rect 9163 27129 9249 27185
rect 9305 27129 9391 27185
rect 9447 27129 9533 27185
rect 9589 27129 9675 27185
rect 9731 27129 9817 27185
rect 9873 27129 9959 27185
rect 10015 27129 10101 27185
rect 10157 27129 10243 27185
rect 10299 27129 10385 27185
rect 10441 27129 10527 27185
rect 10583 27129 10669 27185
rect 10725 27129 10811 27185
rect 10867 27129 10953 27185
rect 11009 27129 11095 27185
rect 11151 27129 11237 27185
rect 11293 27129 11379 27185
rect 11435 27129 11521 27185
rect 11577 27129 11663 27185
rect 11719 27129 11805 27185
rect 11861 27129 11947 27185
rect 12003 27129 12089 27185
rect 12145 27129 12231 27185
rect 12287 27129 12373 27185
rect 12429 27129 12515 27185
rect 12571 27129 12657 27185
rect 12713 27129 12799 27185
rect 12855 27129 12941 27185
rect 12997 27129 13083 27185
rect 13139 27129 13225 27185
rect 13281 27129 13367 27185
rect 13423 27129 13509 27185
rect 13565 27129 13651 27185
rect 13707 27129 13793 27185
rect 13849 27129 13935 27185
rect 13991 27129 14077 27185
rect 14133 27129 14219 27185
rect 14275 27129 14361 27185
rect 14417 27129 14503 27185
rect 14559 27129 14645 27185
rect 14701 27129 14787 27185
rect 14843 27129 15000 27185
rect 0 27043 15000 27129
rect 0 26987 161 27043
rect 217 26987 303 27043
rect 359 26987 445 27043
rect 501 26987 587 27043
rect 643 26987 729 27043
rect 785 26987 871 27043
rect 927 26987 1013 27043
rect 1069 26987 1155 27043
rect 1211 26987 1297 27043
rect 1353 26987 1439 27043
rect 1495 26987 1581 27043
rect 1637 26987 1723 27043
rect 1779 26987 1865 27043
rect 1921 26987 2007 27043
rect 2063 26987 2149 27043
rect 2205 26987 2291 27043
rect 2347 26987 2433 27043
rect 2489 26987 2575 27043
rect 2631 26987 2717 27043
rect 2773 26987 2859 27043
rect 2915 26987 3001 27043
rect 3057 26987 3143 27043
rect 3199 26987 3285 27043
rect 3341 26987 3427 27043
rect 3483 26987 3569 27043
rect 3625 26987 3711 27043
rect 3767 26987 3853 27043
rect 3909 26987 3995 27043
rect 4051 26987 4137 27043
rect 4193 26987 4279 27043
rect 4335 26987 4421 27043
rect 4477 26987 4563 27043
rect 4619 26987 4705 27043
rect 4761 26987 4847 27043
rect 4903 26987 4989 27043
rect 5045 26987 5131 27043
rect 5187 26987 5273 27043
rect 5329 26987 5415 27043
rect 5471 26987 5557 27043
rect 5613 26987 5699 27043
rect 5755 26987 5841 27043
rect 5897 26987 5983 27043
rect 6039 26987 6125 27043
rect 6181 26987 6267 27043
rect 6323 26987 6409 27043
rect 6465 26987 6551 27043
rect 6607 26987 6693 27043
rect 6749 26987 6835 27043
rect 6891 26987 6977 27043
rect 7033 26987 7119 27043
rect 7175 26987 7261 27043
rect 7317 26987 7403 27043
rect 7459 26987 7545 27043
rect 7601 26987 7687 27043
rect 7743 26987 7829 27043
rect 7885 26987 7971 27043
rect 8027 26987 8113 27043
rect 8169 26987 8255 27043
rect 8311 26987 8397 27043
rect 8453 26987 8539 27043
rect 8595 26987 8681 27043
rect 8737 26987 8823 27043
rect 8879 26987 8965 27043
rect 9021 26987 9107 27043
rect 9163 26987 9249 27043
rect 9305 26987 9391 27043
rect 9447 26987 9533 27043
rect 9589 26987 9675 27043
rect 9731 26987 9817 27043
rect 9873 26987 9959 27043
rect 10015 26987 10101 27043
rect 10157 26987 10243 27043
rect 10299 26987 10385 27043
rect 10441 26987 10527 27043
rect 10583 26987 10669 27043
rect 10725 26987 10811 27043
rect 10867 26987 10953 27043
rect 11009 26987 11095 27043
rect 11151 26987 11237 27043
rect 11293 26987 11379 27043
rect 11435 26987 11521 27043
rect 11577 26987 11663 27043
rect 11719 26987 11805 27043
rect 11861 26987 11947 27043
rect 12003 26987 12089 27043
rect 12145 26987 12231 27043
rect 12287 26987 12373 27043
rect 12429 26987 12515 27043
rect 12571 26987 12657 27043
rect 12713 26987 12799 27043
rect 12855 26987 12941 27043
rect 12997 26987 13083 27043
rect 13139 26987 13225 27043
rect 13281 26987 13367 27043
rect 13423 26987 13509 27043
rect 13565 26987 13651 27043
rect 13707 26987 13793 27043
rect 13849 26987 13935 27043
rect 13991 26987 14077 27043
rect 14133 26987 14219 27043
rect 14275 26987 14361 27043
rect 14417 26987 14503 27043
rect 14559 26987 14645 27043
rect 14701 26987 14787 27043
rect 14843 26987 15000 27043
rect 0 26901 15000 26987
rect 0 26845 161 26901
rect 217 26845 303 26901
rect 359 26845 445 26901
rect 501 26845 587 26901
rect 643 26845 729 26901
rect 785 26845 871 26901
rect 927 26845 1013 26901
rect 1069 26845 1155 26901
rect 1211 26845 1297 26901
rect 1353 26845 1439 26901
rect 1495 26845 1581 26901
rect 1637 26845 1723 26901
rect 1779 26845 1865 26901
rect 1921 26845 2007 26901
rect 2063 26845 2149 26901
rect 2205 26845 2291 26901
rect 2347 26845 2433 26901
rect 2489 26845 2575 26901
rect 2631 26845 2717 26901
rect 2773 26845 2859 26901
rect 2915 26845 3001 26901
rect 3057 26845 3143 26901
rect 3199 26845 3285 26901
rect 3341 26845 3427 26901
rect 3483 26845 3569 26901
rect 3625 26845 3711 26901
rect 3767 26845 3853 26901
rect 3909 26845 3995 26901
rect 4051 26845 4137 26901
rect 4193 26845 4279 26901
rect 4335 26845 4421 26901
rect 4477 26845 4563 26901
rect 4619 26845 4705 26901
rect 4761 26845 4847 26901
rect 4903 26845 4989 26901
rect 5045 26845 5131 26901
rect 5187 26845 5273 26901
rect 5329 26845 5415 26901
rect 5471 26845 5557 26901
rect 5613 26845 5699 26901
rect 5755 26845 5841 26901
rect 5897 26845 5983 26901
rect 6039 26845 6125 26901
rect 6181 26845 6267 26901
rect 6323 26845 6409 26901
rect 6465 26845 6551 26901
rect 6607 26845 6693 26901
rect 6749 26845 6835 26901
rect 6891 26845 6977 26901
rect 7033 26845 7119 26901
rect 7175 26845 7261 26901
rect 7317 26845 7403 26901
rect 7459 26845 7545 26901
rect 7601 26845 7687 26901
rect 7743 26845 7829 26901
rect 7885 26845 7971 26901
rect 8027 26845 8113 26901
rect 8169 26845 8255 26901
rect 8311 26845 8397 26901
rect 8453 26845 8539 26901
rect 8595 26845 8681 26901
rect 8737 26845 8823 26901
rect 8879 26845 8965 26901
rect 9021 26845 9107 26901
rect 9163 26845 9249 26901
rect 9305 26845 9391 26901
rect 9447 26845 9533 26901
rect 9589 26845 9675 26901
rect 9731 26845 9817 26901
rect 9873 26845 9959 26901
rect 10015 26845 10101 26901
rect 10157 26845 10243 26901
rect 10299 26845 10385 26901
rect 10441 26845 10527 26901
rect 10583 26845 10669 26901
rect 10725 26845 10811 26901
rect 10867 26845 10953 26901
rect 11009 26845 11095 26901
rect 11151 26845 11237 26901
rect 11293 26845 11379 26901
rect 11435 26845 11521 26901
rect 11577 26845 11663 26901
rect 11719 26845 11805 26901
rect 11861 26845 11947 26901
rect 12003 26845 12089 26901
rect 12145 26845 12231 26901
rect 12287 26845 12373 26901
rect 12429 26845 12515 26901
rect 12571 26845 12657 26901
rect 12713 26845 12799 26901
rect 12855 26845 12941 26901
rect 12997 26845 13083 26901
rect 13139 26845 13225 26901
rect 13281 26845 13367 26901
rect 13423 26845 13509 26901
rect 13565 26845 13651 26901
rect 13707 26845 13793 26901
rect 13849 26845 13935 26901
rect 13991 26845 14077 26901
rect 14133 26845 14219 26901
rect 14275 26845 14361 26901
rect 14417 26845 14503 26901
rect 14559 26845 14645 26901
rect 14701 26845 14787 26901
rect 14843 26845 15000 26901
rect 0 26800 15000 26845
rect 0 26563 15000 26600
rect 0 26507 161 26563
rect 217 26507 303 26563
rect 359 26507 445 26563
rect 501 26507 587 26563
rect 643 26507 729 26563
rect 785 26507 871 26563
rect 927 26507 1013 26563
rect 1069 26507 1155 26563
rect 1211 26507 1297 26563
rect 1353 26507 1439 26563
rect 1495 26507 1581 26563
rect 1637 26507 1723 26563
rect 1779 26507 1865 26563
rect 1921 26507 2007 26563
rect 2063 26507 2149 26563
rect 2205 26507 2291 26563
rect 2347 26507 2433 26563
rect 2489 26507 2575 26563
rect 2631 26507 2717 26563
rect 2773 26507 2859 26563
rect 2915 26507 3001 26563
rect 3057 26507 3143 26563
rect 3199 26507 3285 26563
rect 3341 26507 3427 26563
rect 3483 26507 3569 26563
rect 3625 26507 3711 26563
rect 3767 26507 3853 26563
rect 3909 26507 3995 26563
rect 4051 26507 4137 26563
rect 4193 26507 4279 26563
rect 4335 26507 4421 26563
rect 4477 26507 4563 26563
rect 4619 26507 4705 26563
rect 4761 26507 4847 26563
rect 4903 26507 4989 26563
rect 5045 26507 5131 26563
rect 5187 26507 5273 26563
rect 5329 26507 5415 26563
rect 5471 26507 5557 26563
rect 5613 26507 5699 26563
rect 5755 26507 5841 26563
rect 5897 26507 5983 26563
rect 6039 26507 6125 26563
rect 6181 26507 6267 26563
rect 6323 26507 6409 26563
rect 6465 26507 6551 26563
rect 6607 26507 6693 26563
rect 6749 26507 6835 26563
rect 6891 26507 6977 26563
rect 7033 26507 7119 26563
rect 7175 26507 7261 26563
rect 7317 26507 7403 26563
rect 7459 26507 7545 26563
rect 7601 26507 7687 26563
rect 7743 26507 7829 26563
rect 7885 26507 7971 26563
rect 8027 26507 8113 26563
rect 8169 26507 8255 26563
rect 8311 26507 8397 26563
rect 8453 26507 8539 26563
rect 8595 26507 8681 26563
rect 8737 26507 8823 26563
rect 8879 26507 8965 26563
rect 9021 26507 9107 26563
rect 9163 26507 9249 26563
rect 9305 26507 9391 26563
rect 9447 26507 9533 26563
rect 9589 26507 9675 26563
rect 9731 26507 9817 26563
rect 9873 26507 9959 26563
rect 10015 26507 10101 26563
rect 10157 26507 10243 26563
rect 10299 26507 10385 26563
rect 10441 26507 10527 26563
rect 10583 26507 10669 26563
rect 10725 26507 10811 26563
rect 10867 26507 10953 26563
rect 11009 26507 11095 26563
rect 11151 26507 11237 26563
rect 11293 26507 11379 26563
rect 11435 26507 11521 26563
rect 11577 26507 11663 26563
rect 11719 26507 11805 26563
rect 11861 26507 11947 26563
rect 12003 26507 12089 26563
rect 12145 26507 12231 26563
rect 12287 26507 12373 26563
rect 12429 26507 12515 26563
rect 12571 26507 12657 26563
rect 12713 26507 12799 26563
rect 12855 26507 12941 26563
rect 12997 26507 13083 26563
rect 13139 26507 13225 26563
rect 13281 26507 13367 26563
rect 13423 26507 13509 26563
rect 13565 26507 13651 26563
rect 13707 26507 13793 26563
rect 13849 26507 13935 26563
rect 13991 26507 14077 26563
rect 14133 26507 14219 26563
rect 14275 26507 14361 26563
rect 14417 26507 14503 26563
rect 14559 26507 14645 26563
rect 14701 26507 14787 26563
rect 14843 26507 15000 26563
rect 0 26421 15000 26507
rect 0 26365 161 26421
rect 217 26365 303 26421
rect 359 26365 445 26421
rect 501 26365 587 26421
rect 643 26365 729 26421
rect 785 26365 871 26421
rect 927 26365 1013 26421
rect 1069 26365 1155 26421
rect 1211 26365 1297 26421
rect 1353 26365 1439 26421
rect 1495 26365 1581 26421
rect 1637 26365 1723 26421
rect 1779 26365 1865 26421
rect 1921 26365 2007 26421
rect 2063 26365 2149 26421
rect 2205 26365 2291 26421
rect 2347 26365 2433 26421
rect 2489 26365 2575 26421
rect 2631 26365 2717 26421
rect 2773 26365 2859 26421
rect 2915 26365 3001 26421
rect 3057 26365 3143 26421
rect 3199 26365 3285 26421
rect 3341 26365 3427 26421
rect 3483 26365 3569 26421
rect 3625 26365 3711 26421
rect 3767 26365 3853 26421
rect 3909 26365 3995 26421
rect 4051 26365 4137 26421
rect 4193 26365 4279 26421
rect 4335 26365 4421 26421
rect 4477 26365 4563 26421
rect 4619 26365 4705 26421
rect 4761 26365 4847 26421
rect 4903 26365 4989 26421
rect 5045 26365 5131 26421
rect 5187 26365 5273 26421
rect 5329 26365 5415 26421
rect 5471 26365 5557 26421
rect 5613 26365 5699 26421
rect 5755 26365 5841 26421
rect 5897 26365 5983 26421
rect 6039 26365 6125 26421
rect 6181 26365 6267 26421
rect 6323 26365 6409 26421
rect 6465 26365 6551 26421
rect 6607 26365 6693 26421
rect 6749 26365 6835 26421
rect 6891 26365 6977 26421
rect 7033 26365 7119 26421
rect 7175 26365 7261 26421
rect 7317 26365 7403 26421
rect 7459 26365 7545 26421
rect 7601 26365 7687 26421
rect 7743 26365 7829 26421
rect 7885 26365 7971 26421
rect 8027 26365 8113 26421
rect 8169 26365 8255 26421
rect 8311 26365 8397 26421
rect 8453 26365 8539 26421
rect 8595 26365 8681 26421
rect 8737 26365 8823 26421
rect 8879 26365 8965 26421
rect 9021 26365 9107 26421
rect 9163 26365 9249 26421
rect 9305 26365 9391 26421
rect 9447 26365 9533 26421
rect 9589 26365 9675 26421
rect 9731 26365 9817 26421
rect 9873 26365 9959 26421
rect 10015 26365 10101 26421
rect 10157 26365 10243 26421
rect 10299 26365 10385 26421
rect 10441 26365 10527 26421
rect 10583 26365 10669 26421
rect 10725 26365 10811 26421
rect 10867 26365 10953 26421
rect 11009 26365 11095 26421
rect 11151 26365 11237 26421
rect 11293 26365 11379 26421
rect 11435 26365 11521 26421
rect 11577 26365 11663 26421
rect 11719 26365 11805 26421
rect 11861 26365 11947 26421
rect 12003 26365 12089 26421
rect 12145 26365 12231 26421
rect 12287 26365 12373 26421
rect 12429 26365 12515 26421
rect 12571 26365 12657 26421
rect 12713 26365 12799 26421
rect 12855 26365 12941 26421
rect 12997 26365 13083 26421
rect 13139 26365 13225 26421
rect 13281 26365 13367 26421
rect 13423 26365 13509 26421
rect 13565 26365 13651 26421
rect 13707 26365 13793 26421
rect 13849 26365 13935 26421
rect 13991 26365 14077 26421
rect 14133 26365 14219 26421
rect 14275 26365 14361 26421
rect 14417 26365 14503 26421
rect 14559 26365 14645 26421
rect 14701 26365 14787 26421
rect 14843 26365 15000 26421
rect 0 26279 15000 26365
rect 0 26223 161 26279
rect 217 26223 303 26279
rect 359 26223 445 26279
rect 501 26223 587 26279
rect 643 26223 729 26279
rect 785 26223 871 26279
rect 927 26223 1013 26279
rect 1069 26223 1155 26279
rect 1211 26223 1297 26279
rect 1353 26223 1439 26279
rect 1495 26223 1581 26279
rect 1637 26223 1723 26279
rect 1779 26223 1865 26279
rect 1921 26223 2007 26279
rect 2063 26223 2149 26279
rect 2205 26223 2291 26279
rect 2347 26223 2433 26279
rect 2489 26223 2575 26279
rect 2631 26223 2717 26279
rect 2773 26223 2859 26279
rect 2915 26223 3001 26279
rect 3057 26223 3143 26279
rect 3199 26223 3285 26279
rect 3341 26223 3427 26279
rect 3483 26223 3569 26279
rect 3625 26223 3711 26279
rect 3767 26223 3853 26279
rect 3909 26223 3995 26279
rect 4051 26223 4137 26279
rect 4193 26223 4279 26279
rect 4335 26223 4421 26279
rect 4477 26223 4563 26279
rect 4619 26223 4705 26279
rect 4761 26223 4847 26279
rect 4903 26223 4989 26279
rect 5045 26223 5131 26279
rect 5187 26223 5273 26279
rect 5329 26223 5415 26279
rect 5471 26223 5557 26279
rect 5613 26223 5699 26279
rect 5755 26223 5841 26279
rect 5897 26223 5983 26279
rect 6039 26223 6125 26279
rect 6181 26223 6267 26279
rect 6323 26223 6409 26279
rect 6465 26223 6551 26279
rect 6607 26223 6693 26279
rect 6749 26223 6835 26279
rect 6891 26223 6977 26279
rect 7033 26223 7119 26279
rect 7175 26223 7261 26279
rect 7317 26223 7403 26279
rect 7459 26223 7545 26279
rect 7601 26223 7687 26279
rect 7743 26223 7829 26279
rect 7885 26223 7971 26279
rect 8027 26223 8113 26279
rect 8169 26223 8255 26279
rect 8311 26223 8397 26279
rect 8453 26223 8539 26279
rect 8595 26223 8681 26279
rect 8737 26223 8823 26279
rect 8879 26223 8965 26279
rect 9021 26223 9107 26279
rect 9163 26223 9249 26279
rect 9305 26223 9391 26279
rect 9447 26223 9533 26279
rect 9589 26223 9675 26279
rect 9731 26223 9817 26279
rect 9873 26223 9959 26279
rect 10015 26223 10101 26279
rect 10157 26223 10243 26279
rect 10299 26223 10385 26279
rect 10441 26223 10527 26279
rect 10583 26223 10669 26279
rect 10725 26223 10811 26279
rect 10867 26223 10953 26279
rect 11009 26223 11095 26279
rect 11151 26223 11237 26279
rect 11293 26223 11379 26279
rect 11435 26223 11521 26279
rect 11577 26223 11663 26279
rect 11719 26223 11805 26279
rect 11861 26223 11947 26279
rect 12003 26223 12089 26279
rect 12145 26223 12231 26279
rect 12287 26223 12373 26279
rect 12429 26223 12515 26279
rect 12571 26223 12657 26279
rect 12713 26223 12799 26279
rect 12855 26223 12941 26279
rect 12997 26223 13083 26279
rect 13139 26223 13225 26279
rect 13281 26223 13367 26279
rect 13423 26223 13509 26279
rect 13565 26223 13651 26279
rect 13707 26223 13793 26279
rect 13849 26223 13935 26279
rect 13991 26223 14077 26279
rect 14133 26223 14219 26279
rect 14275 26223 14361 26279
rect 14417 26223 14503 26279
rect 14559 26223 14645 26279
rect 14701 26223 14787 26279
rect 14843 26223 15000 26279
rect 0 26137 15000 26223
rect 0 26081 161 26137
rect 217 26081 303 26137
rect 359 26081 445 26137
rect 501 26081 587 26137
rect 643 26081 729 26137
rect 785 26081 871 26137
rect 927 26081 1013 26137
rect 1069 26081 1155 26137
rect 1211 26081 1297 26137
rect 1353 26081 1439 26137
rect 1495 26081 1581 26137
rect 1637 26081 1723 26137
rect 1779 26081 1865 26137
rect 1921 26081 2007 26137
rect 2063 26081 2149 26137
rect 2205 26081 2291 26137
rect 2347 26081 2433 26137
rect 2489 26081 2575 26137
rect 2631 26081 2717 26137
rect 2773 26081 2859 26137
rect 2915 26081 3001 26137
rect 3057 26081 3143 26137
rect 3199 26081 3285 26137
rect 3341 26081 3427 26137
rect 3483 26081 3569 26137
rect 3625 26081 3711 26137
rect 3767 26081 3853 26137
rect 3909 26081 3995 26137
rect 4051 26081 4137 26137
rect 4193 26081 4279 26137
rect 4335 26081 4421 26137
rect 4477 26081 4563 26137
rect 4619 26081 4705 26137
rect 4761 26081 4847 26137
rect 4903 26081 4989 26137
rect 5045 26081 5131 26137
rect 5187 26081 5273 26137
rect 5329 26081 5415 26137
rect 5471 26081 5557 26137
rect 5613 26081 5699 26137
rect 5755 26081 5841 26137
rect 5897 26081 5983 26137
rect 6039 26081 6125 26137
rect 6181 26081 6267 26137
rect 6323 26081 6409 26137
rect 6465 26081 6551 26137
rect 6607 26081 6693 26137
rect 6749 26081 6835 26137
rect 6891 26081 6977 26137
rect 7033 26081 7119 26137
rect 7175 26081 7261 26137
rect 7317 26081 7403 26137
rect 7459 26081 7545 26137
rect 7601 26081 7687 26137
rect 7743 26081 7829 26137
rect 7885 26081 7971 26137
rect 8027 26081 8113 26137
rect 8169 26081 8255 26137
rect 8311 26081 8397 26137
rect 8453 26081 8539 26137
rect 8595 26081 8681 26137
rect 8737 26081 8823 26137
rect 8879 26081 8965 26137
rect 9021 26081 9107 26137
rect 9163 26081 9249 26137
rect 9305 26081 9391 26137
rect 9447 26081 9533 26137
rect 9589 26081 9675 26137
rect 9731 26081 9817 26137
rect 9873 26081 9959 26137
rect 10015 26081 10101 26137
rect 10157 26081 10243 26137
rect 10299 26081 10385 26137
rect 10441 26081 10527 26137
rect 10583 26081 10669 26137
rect 10725 26081 10811 26137
rect 10867 26081 10953 26137
rect 11009 26081 11095 26137
rect 11151 26081 11237 26137
rect 11293 26081 11379 26137
rect 11435 26081 11521 26137
rect 11577 26081 11663 26137
rect 11719 26081 11805 26137
rect 11861 26081 11947 26137
rect 12003 26081 12089 26137
rect 12145 26081 12231 26137
rect 12287 26081 12373 26137
rect 12429 26081 12515 26137
rect 12571 26081 12657 26137
rect 12713 26081 12799 26137
rect 12855 26081 12941 26137
rect 12997 26081 13083 26137
rect 13139 26081 13225 26137
rect 13281 26081 13367 26137
rect 13423 26081 13509 26137
rect 13565 26081 13651 26137
rect 13707 26081 13793 26137
rect 13849 26081 13935 26137
rect 13991 26081 14077 26137
rect 14133 26081 14219 26137
rect 14275 26081 14361 26137
rect 14417 26081 14503 26137
rect 14559 26081 14645 26137
rect 14701 26081 14787 26137
rect 14843 26081 15000 26137
rect 0 25995 15000 26081
rect 0 25939 161 25995
rect 217 25939 303 25995
rect 359 25939 445 25995
rect 501 25939 587 25995
rect 643 25939 729 25995
rect 785 25939 871 25995
rect 927 25939 1013 25995
rect 1069 25939 1155 25995
rect 1211 25939 1297 25995
rect 1353 25939 1439 25995
rect 1495 25939 1581 25995
rect 1637 25939 1723 25995
rect 1779 25939 1865 25995
rect 1921 25939 2007 25995
rect 2063 25939 2149 25995
rect 2205 25939 2291 25995
rect 2347 25939 2433 25995
rect 2489 25939 2575 25995
rect 2631 25939 2717 25995
rect 2773 25939 2859 25995
rect 2915 25939 3001 25995
rect 3057 25939 3143 25995
rect 3199 25939 3285 25995
rect 3341 25939 3427 25995
rect 3483 25939 3569 25995
rect 3625 25939 3711 25995
rect 3767 25939 3853 25995
rect 3909 25939 3995 25995
rect 4051 25939 4137 25995
rect 4193 25939 4279 25995
rect 4335 25939 4421 25995
rect 4477 25939 4563 25995
rect 4619 25939 4705 25995
rect 4761 25939 4847 25995
rect 4903 25939 4989 25995
rect 5045 25939 5131 25995
rect 5187 25939 5273 25995
rect 5329 25939 5415 25995
rect 5471 25939 5557 25995
rect 5613 25939 5699 25995
rect 5755 25939 5841 25995
rect 5897 25939 5983 25995
rect 6039 25939 6125 25995
rect 6181 25939 6267 25995
rect 6323 25939 6409 25995
rect 6465 25939 6551 25995
rect 6607 25939 6693 25995
rect 6749 25939 6835 25995
rect 6891 25939 6977 25995
rect 7033 25939 7119 25995
rect 7175 25939 7261 25995
rect 7317 25939 7403 25995
rect 7459 25939 7545 25995
rect 7601 25939 7687 25995
rect 7743 25939 7829 25995
rect 7885 25939 7971 25995
rect 8027 25939 8113 25995
rect 8169 25939 8255 25995
rect 8311 25939 8397 25995
rect 8453 25939 8539 25995
rect 8595 25939 8681 25995
rect 8737 25939 8823 25995
rect 8879 25939 8965 25995
rect 9021 25939 9107 25995
rect 9163 25939 9249 25995
rect 9305 25939 9391 25995
rect 9447 25939 9533 25995
rect 9589 25939 9675 25995
rect 9731 25939 9817 25995
rect 9873 25939 9959 25995
rect 10015 25939 10101 25995
rect 10157 25939 10243 25995
rect 10299 25939 10385 25995
rect 10441 25939 10527 25995
rect 10583 25939 10669 25995
rect 10725 25939 10811 25995
rect 10867 25939 10953 25995
rect 11009 25939 11095 25995
rect 11151 25939 11237 25995
rect 11293 25939 11379 25995
rect 11435 25939 11521 25995
rect 11577 25939 11663 25995
rect 11719 25939 11805 25995
rect 11861 25939 11947 25995
rect 12003 25939 12089 25995
rect 12145 25939 12231 25995
rect 12287 25939 12373 25995
rect 12429 25939 12515 25995
rect 12571 25939 12657 25995
rect 12713 25939 12799 25995
rect 12855 25939 12941 25995
rect 12997 25939 13083 25995
rect 13139 25939 13225 25995
rect 13281 25939 13367 25995
rect 13423 25939 13509 25995
rect 13565 25939 13651 25995
rect 13707 25939 13793 25995
rect 13849 25939 13935 25995
rect 13991 25939 14077 25995
rect 14133 25939 14219 25995
rect 14275 25939 14361 25995
rect 14417 25939 14503 25995
rect 14559 25939 14645 25995
rect 14701 25939 14787 25995
rect 14843 25939 15000 25995
rect 0 25853 15000 25939
rect 0 25797 161 25853
rect 217 25797 303 25853
rect 359 25797 445 25853
rect 501 25797 587 25853
rect 643 25797 729 25853
rect 785 25797 871 25853
rect 927 25797 1013 25853
rect 1069 25797 1155 25853
rect 1211 25797 1297 25853
rect 1353 25797 1439 25853
rect 1495 25797 1581 25853
rect 1637 25797 1723 25853
rect 1779 25797 1865 25853
rect 1921 25797 2007 25853
rect 2063 25797 2149 25853
rect 2205 25797 2291 25853
rect 2347 25797 2433 25853
rect 2489 25797 2575 25853
rect 2631 25797 2717 25853
rect 2773 25797 2859 25853
rect 2915 25797 3001 25853
rect 3057 25797 3143 25853
rect 3199 25797 3285 25853
rect 3341 25797 3427 25853
rect 3483 25797 3569 25853
rect 3625 25797 3711 25853
rect 3767 25797 3853 25853
rect 3909 25797 3995 25853
rect 4051 25797 4137 25853
rect 4193 25797 4279 25853
rect 4335 25797 4421 25853
rect 4477 25797 4563 25853
rect 4619 25797 4705 25853
rect 4761 25797 4847 25853
rect 4903 25797 4989 25853
rect 5045 25797 5131 25853
rect 5187 25797 5273 25853
rect 5329 25797 5415 25853
rect 5471 25797 5557 25853
rect 5613 25797 5699 25853
rect 5755 25797 5841 25853
rect 5897 25797 5983 25853
rect 6039 25797 6125 25853
rect 6181 25797 6267 25853
rect 6323 25797 6409 25853
rect 6465 25797 6551 25853
rect 6607 25797 6693 25853
rect 6749 25797 6835 25853
rect 6891 25797 6977 25853
rect 7033 25797 7119 25853
rect 7175 25797 7261 25853
rect 7317 25797 7403 25853
rect 7459 25797 7545 25853
rect 7601 25797 7687 25853
rect 7743 25797 7829 25853
rect 7885 25797 7971 25853
rect 8027 25797 8113 25853
rect 8169 25797 8255 25853
rect 8311 25797 8397 25853
rect 8453 25797 8539 25853
rect 8595 25797 8681 25853
rect 8737 25797 8823 25853
rect 8879 25797 8965 25853
rect 9021 25797 9107 25853
rect 9163 25797 9249 25853
rect 9305 25797 9391 25853
rect 9447 25797 9533 25853
rect 9589 25797 9675 25853
rect 9731 25797 9817 25853
rect 9873 25797 9959 25853
rect 10015 25797 10101 25853
rect 10157 25797 10243 25853
rect 10299 25797 10385 25853
rect 10441 25797 10527 25853
rect 10583 25797 10669 25853
rect 10725 25797 10811 25853
rect 10867 25797 10953 25853
rect 11009 25797 11095 25853
rect 11151 25797 11237 25853
rect 11293 25797 11379 25853
rect 11435 25797 11521 25853
rect 11577 25797 11663 25853
rect 11719 25797 11805 25853
rect 11861 25797 11947 25853
rect 12003 25797 12089 25853
rect 12145 25797 12231 25853
rect 12287 25797 12373 25853
rect 12429 25797 12515 25853
rect 12571 25797 12657 25853
rect 12713 25797 12799 25853
rect 12855 25797 12941 25853
rect 12997 25797 13083 25853
rect 13139 25797 13225 25853
rect 13281 25797 13367 25853
rect 13423 25797 13509 25853
rect 13565 25797 13651 25853
rect 13707 25797 13793 25853
rect 13849 25797 13935 25853
rect 13991 25797 14077 25853
rect 14133 25797 14219 25853
rect 14275 25797 14361 25853
rect 14417 25797 14503 25853
rect 14559 25797 14645 25853
rect 14701 25797 14787 25853
rect 14843 25797 15000 25853
rect 0 25711 15000 25797
rect 0 25655 161 25711
rect 217 25655 303 25711
rect 359 25655 445 25711
rect 501 25655 587 25711
rect 643 25655 729 25711
rect 785 25655 871 25711
rect 927 25655 1013 25711
rect 1069 25655 1155 25711
rect 1211 25655 1297 25711
rect 1353 25655 1439 25711
rect 1495 25655 1581 25711
rect 1637 25655 1723 25711
rect 1779 25655 1865 25711
rect 1921 25655 2007 25711
rect 2063 25655 2149 25711
rect 2205 25655 2291 25711
rect 2347 25655 2433 25711
rect 2489 25655 2575 25711
rect 2631 25655 2717 25711
rect 2773 25655 2859 25711
rect 2915 25655 3001 25711
rect 3057 25655 3143 25711
rect 3199 25655 3285 25711
rect 3341 25655 3427 25711
rect 3483 25655 3569 25711
rect 3625 25655 3711 25711
rect 3767 25655 3853 25711
rect 3909 25655 3995 25711
rect 4051 25655 4137 25711
rect 4193 25655 4279 25711
rect 4335 25655 4421 25711
rect 4477 25655 4563 25711
rect 4619 25655 4705 25711
rect 4761 25655 4847 25711
rect 4903 25655 4989 25711
rect 5045 25655 5131 25711
rect 5187 25655 5273 25711
rect 5329 25655 5415 25711
rect 5471 25655 5557 25711
rect 5613 25655 5699 25711
rect 5755 25655 5841 25711
rect 5897 25655 5983 25711
rect 6039 25655 6125 25711
rect 6181 25655 6267 25711
rect 6323 25655 6409 25711
rect 6465 25655 6551 25711
rect 6607 25655 6693 25711
rect 6749 25655 6835 25711
rect 6891 25655 6977 25711
rect 7033 25655 7119 25711
rect 7175 25655 7261 25711
rect 7317 25655 7403 25711
rect 7459 25655 7545 25711
rect 7601 25655 7687 25711
rect 7743 25655 7829 25711
rect 7885 25655 7971 25711
rect 8027 25655 8113 25711
rect 8169 25655 8255 25711
rect 8311 25655 8397 25711
rect 8453 25655 8539 25711
rect 8595 25655 8681 25711
rect 8737 25655 8823 25711
rect 8879 25655 8965 25711
rect 9021 25655 9107 25711
rect 9163 25655 9249 25711
rect 9305 25655 9391 25711
rect 9447 25655 9533 25711
rect 9589 25655 9675 25711
rect 9731 25655 9817 25711
rect 9873 25655 9959 25711
rect 10015 25655 10101 25711
rect 10157 25655 10243 25711
rect 10299 25655 10385 25711
rect 10441 25655 10527 25711
rect 10583 25655 10669 25711
rect 10725 25655 10811 25711
rect 10867 25655 10953 25711
rect 11009 25655 11095 25711
rect 11151 25655 11237 25711
rect 11293 25655 11379 25711
rect 11435 25655 11521 25711
rect 11577 25655 11663 25711
rect 11719 25655 11805 25711
rect 11861 25655 11947 25711
rect 12003 25655 12089 25711
rect 12145 25655 12231 25711
rect 12287 25655 12373 25711
rect 12429 25655 12515 25711
rect 12571 25655 12657 25711
rect 12713 25655 12799 25711
rect 12855 25655 12941 25711
rect 12997 25655 13083 25711
rect 13139 25655 13225 25711
rect 13281 25655 13367 25711
rect 13423 25655 13509 25711
rect 13565 25655 13651 25711
rect 13707 25655 13793 25711
rect 13849 25655 13935 25711
rect 13991 25655 14077 25711
rect 14133 25655 14219 25711
rect 14275 25655 14361 25711
rect 14417 25655 14503 25711
rect 14559 25655 14645 25711
rect 14701 25655 14787 25711
rect 14843 25655 15000 25711
rect 0 25569 15000 25655
rect 0 25513 161 25569
rect 217 25513 303 25569
rect 359 25513 445 25569
rect 501 25513 587 25569
rect 643 25513 729 25569
rect 785 25513 871 25569
rect 927 25513 1013 25569
rect 1069 25513 1155 25569
rect 1211 25513 1297 25569
rect 1353 25513 1439 25569
rect 1495 25513 1581 25569
rect 1637 25513 1723 25569
rect 1779 25513 1865 25569
rect 1921 25513 2007 25569
rect 2063 25513 2149 25569
rect 2205 25513 2291 25569
rect 2347 25513 2433 25569
rect 2489 25513 2575 25569
rect 2631 25513 2717 25569
rect 2773 25513 2859 25569
rect 2915 25513 3001 25569
rect 3057 25513 3143 25569
rect 3199 25513 3285 25569
rect 3341 25513 3427 25569
rect 3483 25513 3569 25569
rect 3625 25513 3711 25569
rect 3767 25513 3853 25569
rect 3909 25513 3995 25569
rect 4051 25513 4137 25569
rect 4193 25513 4279 25569
rect 4335 25513 4421 25569
rect 4477 25513 4563 25569
rect 4619 25513 4705 25569
rect 4761 25513 4847 25569
rect 4903 25513 4989 25569
rect 5045 25513 5131 25569
rect 5187 25513 5273 25569
rect 5329 25513 5415 25569
rect 5471 25513 5557 25569
rect 5613 25513 5699 25569
rect 5755 25513 5841 25569
rect 5897 25513 5983 25569
rect 6039 25513 6125 25569
rect 6181 25513 6267 25569
rect 6323 25513 6409 25569
rect 6465 25513 6551 25569
rect 6607 25513 6693 25569
rect 6749 25513 6835 25569
rect 6891 25513 6977 25569
rect 7033 25513 7119 25569
rect 7175 25513 7261 25569
rect 7317 25513 7403 25569
rect 7459 25513 7545 25569
rect 7601 25513 7687 25569
rect 7743 25513 7829 25569
rect 7885 25513 7971 25569
rect 8027 25513 8113 25569
rect 8169 25513 8255 25569
rect 8311 25513 8397 25569
rect 8453 25513 8539 25569
rect 8595 25513 8681 25569
rect 8737 25513 8823 25569
rect 8879 25513 8965 25569
rect 9021 25513 9107 25569
rect 9163 25513 9249 25569
rect 9305 25513 9391 25569
rect 9447 25513 9533 25569
rect 9589 25513 9675 25569
rect 9731 25513 9817 25569
rect 9873 25513 9959 25569
rect 10015 25513 10101 25569
rect 10157 25513 10243 25569
rect 10299 25513 10385 25569
rect 10441 25513 10527 25569
rect 10583 25513 10669 25569
rect 10725 25513 10811 25569
rect 10867 25513 10953 25569
rect 11009 25513 11095 25569
rect 11151 25513 11237 25569
rect 11293 25513 11379 25569
rect 11435 25513 11521 25569
rect 11577 25513 11663 25569
rect 11719 25513 11805 25569
rect 11861 25513 11947 25569
rect 12003 25513 12089 25569
rect 12145 25513 12231 25569
rect 12287 25513 12373 25569
rect 12429 25513 12515 25569
rect 12571 25513 12657 25569
rect 12713 25513 12799 25569
rect 12855 25513 12941 25569
rect 12997 25513 13083 25569
rect 13139 25513 13225 25569
rect 13281 25513 13367 25569
rect 13423 25513 13509 25569
rect 13565 25513 13651 25569
rect 13707 25513 13793 25569
rect 13849 25513 13935 25569
rect 13991 25513 14077 25569
rect 14133 25513 14219 25569
rect 14275 25513 14361 25569
rect 14417 25513 14503 25569
rect 14559 25513 14645 25569
rect 14701 25513 14787 25569
rect 14843 25513 15000 25569
rect 0 25427 15000 25513
rect 0 25371 161 25427
rect 217 25371 303 25427
rect 359 25371 445 25427
rect 501 25371 587 25427
rect 643 25371 729 25427
rect 785 25371 871 25427
rect 927 25371 1013 25427
rect 1069 25371 1155 25427
rect 1211 25371 1297 25427
rect 1353 25371 1439 25427
rect 1495 25371 1581 25427
rect 1637 25371 1723 25427
rect 1779 25371 1865 25427
rect 1921 25371 2007 25427
rect 2063 25371 2149 25427
rect 2205 25371 2291 25427
rect 2347 25371 2433 25427
rect 2489 25371 2575 25427
rect 2631 25371 2717 25427
rect 2773 25371 2859 25427
rect 2915 25371 3001 25427
rect 3057 25371 3143 25427
rect 3199 25371 3285 25427
rect 3341 25371 3427 25427
rect 3483 25371 3569 25427
rect 3625 25371 3711 25427
rect 3767 25371 3853 25427
rect 3909 25371 3995 25427
rect 4051 25371 4137 25427
rect 4193 25371 4279 25427
rect 4335 25371 4421 25427
rect 4477 25371 4563 25427
rect 4619 25371 4705 25427
rect 4761 25371 4847 25427
rect 4903 25371 4989 25427
rect 5045 25371 5131 25427
rect 5187 25371 5273 25427
rect 5329 25371 5415 25427
rect 5471 25371 5557 25427
rect 5613 25371 5699 25427
rect 5755 25371 5841 25427
rect 5897 25371 5983 25427
rect 6039 25371 6125 25427
rect 6181 25371 6267 25427
rect 6323 25371 6409 25427
rect 6465 25371 6551 25427
rect 6607 25371 6693 25427
rect 6749 25371 6835 25427
rect 6891 25371 6977 25427
rect 7033 25371 7119 25427
rect 7175 25371 7261 25427
rect 7317 25371 7403 25427
rect 7459 25371 7545 25427
rect 7601 25371 7687 25427
rect 7743 25371 7829 25427
rect 7885 25371 7971 25427
rect 8027 25371 8113 25427
rect 8169 25371 8255 25427
rect 8311 25371 8397 25427
rect 8453 25371 8539 25427
rect 8595 25371 8681 25427
rect 8737 25371 8823 25427
rect 8879 25371 8965 25427
rect 9021 25371 9107 25427
rect 9163 25371 9249 25427
rect 9305 25371 9391 25427
rect 9447 25371 9533 25427
rect 9589 25371 9675 25427
rect 9731 25371 9817 25427
rect 9873 25371 9959 25427
rect 10015 25371 10101 25427
rect 10157 25371 10243 25427
rect 10299 25371 10385 25427
rect 10441 25371 10527 25427
rect 10583 25371 10669 25427
rect 10725 25371 10811 25427
rect 10867 25371 10953 25427
rect 11009 25371 11095 25427
rect 11151 25371 11237 25427
rect 11293 25371 11379 25427
rect 11435 25371 11521 25427
rect 11577 25371 11663 25427
rect 11719 25371 11805 25427
rect 11861 25371 11947 25427
rect 12003 25371 12089 25427
rect 12145 25371 12231 25427
rect 12287 25371 12373 25427
rect 12429 25371 12515 25427
rect 12571 25371 12657 25427
rect 12713 25371 12799 25427
rect 12855 25371 12941 25427
rect 12997 25371 13083 25427
rect 13139 25371 13225 25427
rect 13281 25371 13367 25427
rect 13423 25371 13509 25427
rect 13565 25371 13651 25427
rect 13707 25371 13793 25427
rect 13849 25371 13935 25427
rect 13991 25371 14077 25427
rect 14133 25371 14219 25427
rect 14275 25371 14361 25427
rect 14417 25371 14503 25427
rect 14559 25371 14645 25427
rect 14701 25371 14787 25427
rect 14843 25371 15000 25427
rect 0 25285 15000 25371
rect 0 25229 161 25285
rect 217 25229 303 25285
rect 359 25229 445 25285
rect 501 25229 587 25285
rect 643 25229 729 25285
rect 785 25229 871 25285
rect 927 25229 1013 25285
rect 1069 25229 1155 25285
rect 1211 25229 1297 25285
rect 1353 25229 1439 25285
rect 1495 25229 1581 25285
rect 1637 25229 1723 25285
rect 1779 25229 1865 25285
rect 1921 25229 2007 25285
rect 2063 25229 2149 25285
rect 2205 25229 2291 25285
rect 2347 25229 2433 25285
rect 2489 25229 2575 25285
rect 2631 25229 2717 25285
rect 2773 25229 2859 25285
rect 2915 25229 3001 25285
rect 3057 25229 3143 25285
rect 3199 25229 3285 25285
rect 3341 25229 3427 25285
rect 3483 25229 3569 25285
rect 3625 25229 3711 25285
rect 3767 25229 3853 25285
rect 3909 25229 3995 25285
rect 4051 25229 4137 25285
rect 4193 25229 4279 25285
rect 4335 25229 4421 25285
rect 4477 25229 4563 25285
rect 4619 25229 4705 25285
rect 4761 25229 4847 25285
rect 4903 25229 4989 25285
rect 5045 25229 5131 25285
rect 5187 25229 5273 25285
rect 5329 25229 5415 25285
rect 5471 25229 5557 25285
rect 5613 25229 5699 25285
rect 5755 25229 5841 25285
rect 5897 25229 5983 25285
rect 6039 25229 6125 25285
rect 6181 25229 6267 25285
rect 6323 25229 6409 25285
rect 6465 25229 6551 25285
rect 6607 25229 6693 25285
rect 6749 25229 6835 25285
rect 6891 25229 6977 25285
rect 7033 25229 7119 25285
rect 7175 25229 7261 25285
rect 7317 25229 7403 25285
rect 7459 25229 7545 25285
rect 7601 25229 7687 25285
rect 7743 25229 7829 25285
rect 7885 25229 7971 25285
rect 8027 25229 8113 25285
rect 8169 25229 8255 25285
rect 8311 25229 8397 25285
rect 8453 25229 8539 25285
rect 8595 25229 8681 25285
rect 8737 25229 8823 25285
rect 8879 25229 8965 25285
rect 9021 25229 9107 25285
rect 9163 25229 9249 25285
rect 9305 25229 9391 25285
rect 9447 25229 9533 25285
rect 9589 25229 9675 25285
rect 9731 25229 9817 25285
rect 9873 25229 9959 25285
rect 10015 25229 10101 25285
rect 10157 25229 10243 25285
rect 10299 25229 10385 25285
rect 10441 25229 10527 25285
rect 10583 25229 10669 25285
rect 10725 25229 10811 25285
rect 10867 25229 10953 25285
rect 11009 25229 11095 25285
rect 11151 25229 11237 25285
rect 11293 25229 11379 25285
rect 11435 25229 11521 25285
rect 11577 25229 11663 25285
rect 11719 25229 11805 25285
rect 11861 25229 11947 25285
rect 12003 25229 12089 25285
rect 12145 25229 12231 25285
rect 12287 25229 12373 25285
rect 12429 25229 12515 25285
rect 12571 25229 12657 25285
rect 12713 25229 12799 25285
rect 12855 25229 12941 25285
rect 12997 25229 13083 25285
rect 13139 25229 13225 25285
rect 13281 25229 13367 25285
rect 13423 25229 13509 25285
rect 13565 25229 13651 25285
rect 13707 25229 13793 25285
rect 13849 25229 13935 25285
rect 13991 25229 14077 25285
rect 14133 25229 14219 25285
rect 14275 25229 14361 25285
rect 14417 25229 14503 25285
rect 14559 25229 14645 25285
rect 14701 25229 14787 25285
rect 14843 25229 15000 25285
rect 0 25200 15000 25229
rect 0 24963 15000 25000
rect 0 24907 161 24963
rect 217 24907 303 24963
rect 359 24907 445 24963
rect 501 24907 587 24963
rect 643 24907 729 24963
rect 785 24907 871 24963
rect 927 24907 1013 24963
rect 1069 24907 1155 24963
rect 1211 24907 1297 24963
rect 1353 24907 1439 24963
rect 1495 24907 1581 24963
rect 1637 24907 1723 24963
rect 1779 24907 1865 24963
rect 1921 24907 2007 24963
rect 2063 24907 2149 24963
rect 2205 24907 2291 24963
rect 2347 24907 2433 24963
rect 2489 24907 2575 24963
rect 2631 24907 2717 24963
rect 2773 24907 2859 24963
rect 2915 24907 3001 24963
rect 3057 24907 3143 24963
rect 3199 24907 3285 24963
rect 3341 24907 3427 24963
rect 3483 24907 3569 24963
rect 3625 24907 3711 24963
rect 3767 24907 3853 24963
rect 3909 24907 3995 24963
rect 4051 24907 4137 24963
rect 4193 24907 4279 24963
rect 4335 24907 4421 24963
rect 4477 24907 4563 24963
rect 4619 24907 4705 24963
rect 4761 24907 4847 24963
rect 4903 24907 4989 24963
rect 5045 24907 5131 24963
rect 5187 24907 5273 24963
rect 5329 24907 5415 24963
rect 5471 24907 5557 24963
rect 5613 24907 5699 24963
rect 5755 24907 5841 24963
rect 5897 24907 5983 24963
rect 6039 24907 6125 24963
rect 6181 24907 6267 24963
rect 6323 24907 6409 24963
rect 6465 24907 6551 24963
rect 6607 24907 6693 24963
rect 6749 24907 6835 24963
rect 6891 24907 6977 24963
rect 7033 24907 7119 24963
rect 7175 24907 7261 24963
rect 7317 24907 7403 24963
rect 7459 24907 7545 24963
rect 7601 24907 7687 24963
rect 7743 24907 7829 24963
rect 7885 24907 7971 24963
rect 8027 24907 8113 24963
rect 8169 24907 8255 24963
rect 8311 24907 8397 24963
rect 8453 24907 8539 24963
rect 8595 24907 8681 24963
rect 8737 24907 8823 24963
rect 8879 24907 8965 24963
rect 9021 24907 9107 24963
rect 9163 24907 9249 24963
rect 9305 24907 9391 24963
rect 9447 24907 9533 24963
rect 9589 24907 9675 24963
rect 9731 24907 9817 24963
rect 9873 24907 9959 24963
rect 10015 24907 10101 24963
rect 10157 24907 10243 24963
rect 10299 24907 10385 24963
rect 10441 24907 10527 24963
rect 10583 24907 10669 24963
rect 10725 24907 10811 24963
rect 10867 24907 10953 24963
rect 11009 24907 11095 24963
rect 11151 24907 11237 24963
rect 11293 24907 11379 24963
rect 11435 24907 11521 24963
rect 11577 24907 11663 24963
rect 11719 24907 11805 24963
rect 11861 24907 11947 24963
rect 12003 24907 12089 24963
rect 12145 24907 12231 24963
rect 12287 24907 12373 24963
rect 12429 24907 12515 24963
rect 12571 24907 12657 24963
rect 12713 24907 12799 24963
rect 12855 24907 12941 24963
rect 12997 24907 13083 24963
rect 13139 24907 13225 24963
rect 13281 24907 13367 24963
rect 13423 24907 13509 24963
rect 13565 24907 13651 24963
rect 13707 24907 13793 24963
rect 13849 24907 13935 24963
rect 13991 24907 14077 24963
rect 14133 24907 14219 24963
rect 14275 24907 14361 24963
rect 14417 24907 14503 24963
rect 14559 24907 14645 24963
rect 14701 24907 14787 24963
rect 14843 24907 15000 24963
rect 0 24821 15000 24907
rect 0 24765 161 24821
rect 217 24765 303 24821
rect 359 24765 445 24821
rect 501 24765 587 24821
rect 643 24765 729 24821
rect 785 24765 871 24821
rect 927 24765 1013 24821
rect 1069 24765 1155 24821
rect 1211 24765 1297 24821
rect 1353 24765 1439 24821
rect 1495 24765 1581 24821
rect 1637 24765 1723 24821
rect 1779 24765 1865 24821
rect 1921 24765 2007 24821
rect 2063 24765 2149 24821
rect 2205 24765 2291 24821
rect 2347 24765 2433 24821
rect 2489 24765 2575 24821
rect 2631 24765 2717 24821
rect 2773 24765 2859 24821
rect 2915 24765 3001 24821
rect 3057 24765 3143 24821
rect 3199 24765 3285 24821
rect 3341 24765 3427 24821
rect 3483 24765 3569 24821
rect 3625 24765 3711 24821
rect 3767 24765 3853 24821
rect 3909 24765 3995 24821
rect 4051 24765 4137 24821
rect 4193 24765 4279 24821
rect 4335 24765 4421 24821
rect 4477 24765 4563 24821
rect 4619 24765 4705 24821
rect 4761 24765 4847 24821
rect 4903 24765 4989 24821
rect 5045 24765 5131 24821
rect 5187 24765 5273 24821
rect 5329 24765 5415 24821
rect 5471 24765 5557 24821
rect 5613 24765 5699 24821
rect 5755 24765 5841 24821
rect 5897 24765 5983 24821
rect 6039 24765 6125 24821
rect 6181 24765 6267 24821
rect 6323 24765 6409 24821
rect 6465 24765 6551 24821
rect 6607 24765 6693 24821
rect 6749 24765 6835 24821
rect 6891 24765 6977 24821
rect 7033 24765 7119 24821
rect 7175 24765 7261 24821
rect 7317 24765 7403 24821
rect 7459 24765 7545 24821
rect 7601 24765 7687 24821
rect 7743 24765 7829 24821
rect 7885 24765 7971 24821
rect 8027 24765 8113 24821
rect 8169 24765 8255 24821
rect 8311 24765 8397 24821
rect 8453 24765 8539 24821
rect 8595 24765 8681 24821
rect 8737 24765 8823 24821
rect 8879 24765 8965 24821
rect 9021 24765 9107 24821
rect 9163 24765 9249 24821
rect 9305 24765 9391 24821
rect 9447 24765 9533 24821
rect 9589 24765 9675 24821
rect 9731 24765 9817 24821
rect 9873 24765 9959 24821
rect 10015 24765 10101 24821
rect 10157 24765 10243 24821
rect 10299 24765 10385 24821
rect 10441 24765 10527 24821
rect 10583 24765 10669 24821
rect 10725 24765 10811 24821
rect 10867 24765 10953 24821
rect 11009 24765 11095 24821
rect 11151 24765 11237 24821
rect 11293 24765 11379 24821
rect 11435 24765 11521 24821
rect 11577 24765 11663 24821
rect 11719 24765 11805 24821
rect 11861 24765 11947 24821
rect 12003 24765 12089 24821
rect 12145 24765 12231 24821
rect 12287 24765 12373 24821
rect 12429 24765 12515 24821
rect 12571 24765 12657 24821
rect 12713 24765 12799 24821
rect 12855 24765 12941 24821
rect 12997 24765 13083 24821
rect 13139 24765 13225 24821
rect 13281 24765 13367 24821
rect 13423 24765 13509 24821
rect 13565 24765 13651 24821
rect 13707 24765 13793 24821
rect 13849 24765 13935 24821
rect 13991 24765 14077 24821
rect 14133 24765 14219 24821
rect 14275 24765 14361 24821
rect 14417 24765 14503 24821
rect 14559 24765 14645 24821
rect 14701 24765 14787 24821
rect 14843 24765 15000 24821
rect 0 24679 15000 24765
rect 0 24623 161 24679
rect 217 24623 303 24679
rect 359 24623 445 24679
rect 501 24623 587 24679
rect 643 24623 729 24679
rect 785 24623 871 24679
rect 927 24623 1013 24679
rect 1069 24623 1155 24679
rect 1211 24623 1297 24679
rect 1353 24623 1439 24679
rect 1495 24623 1581 24679
rect 1637 24623 1723 24679
rect 1779 24623 1865 24679
rect 1921 24623 2007 24679
rect 2063 24623 2149 24679
rect 2205 24623 2291 24679
rect 2347 24623 2433 24679
rect 2489 24623 2575 24679
rect 2631 24623 2717 24679
rect 2773 24623 2859 24679
rect 2915 24623 3001 24679
rect 3057 24623 3143 24679
rect 3199 24623 3285 24679
rect 3341 24623 3427 24679
rect 3483 24623 3569 24679
rect 3625 24623 3711 24679
rect 3767 24623 3853 24679
rect 3909 24623 3995 24679
rect 4051 24623 4137 24679
rect 4193 24623 4279 24679
rect 4335 24623 4421 24679
rect 4477 24623 4563 24679
rect 4619 24623 4705 24679
rect 4761 24623 4847 24679
rect 4903 24623 4989 24679
rect 5045 24623 5131 24679
rect 5187 24623 5273 24679
rect 5329 24623 5415 24679
rect 5471 24623 5557 24679
rect 5613 24623 5699 24679
rect 5755 24623 5841 24679
rect 5897 24623 5983 24679
rect 6039 24623 6125 24679
rect 6181 24623 6267 24679
rect 6323 24623 6409 24679
rect 6465 24623 6551 24679
rect 6607 24623 6693 24679
rect 6749 24623 6835 24679
rect 6891 24623 6977 24679
rect 7033 24623 7119 24679
rect 7175 24623 7261 24679
rect 7317 24623 7403 24679
rect 7459 24623 7545 24679
rect 7601 24623 7687 24679
rect 7743 24623 7829 24679
rect 7885 24623 7971 24679
rect 8027 24623 8113 24679
rect 8169 24623 8255 24679
rect 8311 24623 8397 24679
rect 8453 24623 8539 24679
rect 8595 24623 8681 24679
rect 8737 24623 8823 24679
rect 8879 24623 8965 24679
rect 9021 24623 9107 24679
rect 9163 24623 9249 24679
rect 9305 24623 9391 24679
rect 9447 24623 9533 24679
rect 9589 24623 9675 24679
rect 9731 24623 9817 24679
rect 9873 24623 9959 24679
rect 10015 24623 10101 24679
rect 10157 24623 10243 24679
rect 10299 24623 10385 24679
rect 10441 24623 10527 24679
rect 10583 24623 10669 24679
rect 10725 24623 10811 24679
rect 10867 24623 10953 24679
rect 11009 24623 11095 24679
rect 11151 24623 11237 24679
rect 11293 24623 11379 24679
rect 11435 24623 11521 24679
rect 11577 24623 11663 24679
rect 11719 24623 11805 24679
rect 11861 24623 11947 24679
rect 12003 24623 12089 24679
rect 12145 24623 12231 24679
rect 12287 24623 12373 24679
rect 12429 24623 12515 24679
rect 12571 24623 12657 24679
rect 12713 24623 12799 24679
rect 12855 24623 12941 24679
rect 12997 24623 13083 24679
rect 13139 24623 13225 24679
rect 13281 24623 13367 24679
rect 13423 24623 13509 24679
rect 13565 24623 13651 24679
rect 13707 24623 13793 24679
rect 13849 24623 13935 24679
rect 13991 24623 14077 24679
rect 14133 24623 14219 24679
rect 14275 24623 14361 24679
rect 14417 24623 14503 24679
rect 14559 24623 14645 24679
rect 14701 24623 14787 24679
rect 14843 24623 15000 24679
rect 0 24537 15000 24623
rect 0 24481 161 24537
rect 217 24481 303 24537
rect 359 24481 445 24537
rect 501 24481 587 24537
rect 643 24481 729 24537
rect 785 24481 871 24537
rect 927 24481 1013 24537
rect 1069 24481 1155 24537
rect 1211 24481 1297 24537
rect 1353 24481 1439 24537
rect 1495 24481 1581 24537
rect 1637 24481 1723 24537
rect 1779 24481 1865 24537
rect 1921 24481 2007 24537
rect 2063 24481 2149 24537
rect 2205 24481 2291 24537
rect 2347 24481 2433 24537
rect 2489 24481 2575 24537
rect 2631 24481 2717 24537
rect 2773 24481 2859 24537
rect 2915 24481 3001 24537
rect 3057 24481 3143 24537
rect 3199 24481 3285 24537
rect 3341 24481 3427 24537
rect 3483 24481 3569 24537
rect 3625 24481 3711 24537
rect 3767 24481 3853 24537
rect 3909 24481 3995 24537
rect 4051 24481 4137 24537
rect 4193 24481 4279 24537
rect 4335 24481 4421 24537
rect 4477 24481 4563 24537
rect 4619 24481 4705 24537
rect 4761 24481 4847 24537
rect 4903 24481 4989 24537
rect 5045 24481 5131 24537
rect 5187 24481 5273 24537
rect 5329 24481 5415 24537
rect 5471 24481 5557 24537
rect 5613 24481 5699 24537
rect 5755 24481 5841 24537
rect 5897 24481 5983 24537
rect 6039 24481 6125 24537
rect 6181 24481 6267 24537
rect 6323 24481 6409 24537
rect 6465 24481 6551 24537
rect 6607 24481 6693 24537
rect 6749 24481 6835 24537
rect 6891 24481 6977 24537
rect 7033 24481 7119 24537
rect 7175 24481 7261 24537
rect 7317 24481 7403 24537
rect 7459 24481 7545 24537
rect 7601 24481 7687 24537
rect 7743 24481 7829 24537
rect 7885 24481 7971 24537
rect 8027 24481 8113 24537
rect 8169 24481 8255 24537
rect 8311 24481 8397 24537
rect 8453 24481 8539 24537
rect 8595 24481 8681 24537
rect 8737 24481 8823 24537
rect 8879 24481 8965 24537
rect 9021 24481 9107 24537
rect 9163 24481 9249 24537
rect 9305 24481 9391 24537
rect 9447 24481 9533 24537
rect 9589 24481 9675 24537
rect 9731 24481 9817 24537
rect 9873 24481 9959 24537
rect 10015 24481 10101 24537
rect 10157 24481 10243 24537
rect 10299 24481 10385 24537
rect 10441 24481 10527 24537
rect 10583 24481 10669 24537
rect 10725 24481 10811 24537
rect 10867 24481 10953 24537
rect 11009 24481 11095 24537
rect 11151 24481 11237 24537
rect 11293 24481 11379 24537
rect 11435 24481 11521 24537
rect 11577 24481 11663 24537
rect 11719 24481 11805 24537
rect 11861 24481 11947 24537
rect 12003 24481 12089 24537
rect 12145 24481 12231 24537
rect 12287 24481 12373 24537
rect 12429 24481 12515 24537
rect 12571 24481 12657 24537
rect 12713 24481 12799 24537
rect 12855 24481 12941 24537
rect 12997 24481 13083 24537
rect 13139 24481 13225 24537
rect 13281 24481 13367 24537
rect 13423 24481 13509 24537
rect 13565 24481 13651 24537
rect 13707 24481 13793 24537
rect 13849 24481 13935 24537
rect 13991 24481 14077 24537
rect 14133 24481 14219 24537
rect 14275 24481 14361 24537
rect 14417 24481 14503 24537
rect 14559 24481 14645 24537
rect 14701 24481 14787 24537
rect 14843 24481 15000 24537
rect 0 24395 15000 24481
rect 0 24339 161 24395
rect 217 24339 303 24395
rect 359 24339 445 24395
rect 501 24339 587 24395
rect 643 24339 729 24395
rect 785 24339 871 24395
rect 927 24339 1013 24395
rect 1069 24339 1155 24395
rect 1211 24339 1297 24395
rect 1353 24339 1439 24395
rect 1495 24339 1581 24395
rect 1637 24339 1723 24395
rect 1779 24339 1865 24395
rect 1921 24339 2007 24395
rect 2063 24339 2149 24395
rect 2205 24339 2291 24395
rect 2347 24339 2433 24395
rect 2489 24339 2575 24395
rect 2631 24339 2717 24395
rect 2773 24339 2859 24395
rect 2915 24339 3001 24395
rect 3057 24339 3143 24395
rect 3199 24339 3285 24395
rect 3341 24339 3427 24395
rect 3483 24339 3569 24395
rect 3625 24339 3711 24395
rect 3767 24339 3853 24395
rect 3909 24339 3995 24395
rect 4051 24339 4137 24395
rect 4193 24339 4279 24395
rect 4335 24339 4421 24395
rect 4477 24339 4563 24395
rect 4619 24339 4705 24395
rect 4761 24339 4847 24395
rect 4903 24339 4989 24395
rect 5045 24339 5131 24395
rect 5187 24339 5273 24395
rect 5329 24339 5415 24395
rect 5471 24339 5557 24395
rect 5613 24339 5699 24395
rect 5755 24339 5841 24395
rect 5897 24339 5983 24395
rect 6039 24339 6125 24395
rect 6181 24339 6267 24395
rect 6323 24339 6409 24395
rect 6465 24339 6551 24395
rect 6607 24339 6693 24395
rect 6749 24339 6835 24395
rect 6891 24339 6977 24395
rect 7033 24339 7119 24395
rect 7175 24339 7261 24395
rect 7317 24339 7403 24395
rect 7459 24339 7545 24395
rect 7601 24339 7687 24395
rect 7743 24339 7829 24395
rect 7885 24339 7971 24395
rect 8027 24339 8113 24395
rect 8169 24339 8255 24395
rect 8311 24339 8397 24395
rect 8453 24339 8539 24395
rect 8595 24339 8681 24395
rect 8737 24339 8823 24395
rect 8879 24339 8965 24395
rect 9021 24339 9107 24395
rect 9163 24339 9249 24395
rect 9305 24339 9391 24395
rect 9447 24339 9533 24395
rect 9589 24339 9675 24395
rect 9731 24339 9817 24395
rect 9873 24339 9959 24395
rect 10015 24339 10101 24395
rect 10157 24339 10243 24395
rect 10299 24339 10385 24395
rect 10441 24339 10527 24395
rect 10583 24339 10669 24395
rect 10725 24339 10811 24395
rect 10867 24339 10953 24395
rect 11009 24339 11095 24395
rect 11151 24339 11237 24395
rect 11293 24339 11379 24395
rect 11435 24339 11521 24395
rect 11577 24339 11663 24395
rect 11719 24339 11805 24395
rect 11861 24339 11947 24395
rect 12003 24339 12089 24395
rect 12145 24339 12231 24395
rect 12287 24339 12373 24395
rect 12429 24339 12515 24395
rect 12571 24339 12657 24395
rect 12713 24339 12799 24395
rect 12855 24339 12941 24395
rect 12997 24339 13083 24395
rect 13139 24339 13225 24395
rect 13281 24339 13367 24395
rect 13423 24339 13509 24395
rect 13565 24339 13651 24395
rect 13707 24339 13793 24395
rect 13849 24339 13935 24395
rect 13991 24339 14077 24395
rect 14133 24339 14219 24395
rect 14275 24339 14361 24395
rect 14417 24339 14503 24395
rect 14559 24339 14645 24395
rect 14701 24339 14787 24395
rect 14843 24339 15000 24395
rect 0 24253 15000 24339
rect 0 24197 161 24253
rect 217 24197 303 24253
rect 359 24197 445 24253
rect 501 24197 587 24253
rect 643 24197 729 24253
rect 785 24197 871 24253
rect 927 24197 1013 24253
rect 1069 24197 1155 24253
rect 1211 24197 1297 24253
rect 1353 24197 1439 24253
rect 1495 24197 1581 24253
rect 1637 24197 1723 24253
rect 1779 24197 1865 24253
rect 1921 24197 2007 24253
rect 2063 24197 2149 24253
rect 2205 24197 2291 24253
rect 2347 24197 2433 24253
rect 2489 24197 2575 24253
rect 2631 24197 2717 24253
rect 2773 24197 2859 24253
rect 2915 24197 3001 24253
rect 3057 24197 3143 24253
rect 3199 24197 3285 24253
rect 3341 24197 3427 24253
rect 3483 24197 3569 24253
rect 3625 24197 3711 24253
rect 3767 24197 3853 24253
rect 3909 24197 3995 24253
rect 4051 24197 4137 24253
rect 4193 24197 4279 24253
rect 4335 24197 4421 24253
rect 4477 24197 4563 24253
rect 4619 24197 4705 24253
rect 4761 24197 4847 24253
rect 4903 24197 4989 24253
rect 5045 24197 5131 24253
rect 5187 24197 5273 24253
rect 5329 24197 5415 24253
rect 5471 24197 5557 24253
rect 5613 24197 5699 24253
rect 5755 24197 5841 24253
rect 5897 24197 5983 24253
rect 6039 24197 6125 24253
rect 6181 24197 6267 24253
rect 6323 24197 6409 24253
rect 6465 24197 6551 24253
rect 6607 24197 6693 24253
rect 6749 24197 6835 24253
rect 6891 24197 6977 24253
rect 7033 24197 7119 24253
rect 7175 24197 7261 24253
rect 7317 24197 7403 24253
rect 7459 24197 7545 24253
rect 7601 24197 7687 24253
rect 7743 24197 7829 24253
rect 7885 24197 7971 24253
rect 8027 24197 8113 24253
rect 8169 24197 8255 24253
rect 8311 24197 8397 24253
rect 8453 24197 8539 24253
rect 8595 24197 8681 24253
rect 8737 24197 8823 24253
rect 8879 24197 8965 24253
rect 9021 24197 9107 24253
rect 9163 24197 9249 24253
rect 9305 24197 9391 24253
rect 9447 24197 9533 24253
rect 9589 24197 9675 24253
rect 9731 24197 9817 24253
rect 9873 24197 9959 24253
rect 10015 24197 10101 24253
rect 10157 24197 10243 24253
rect 10299 24197 10385 24253
rect 10441 24197 10527 24253
rect 10583 24197 10669 24253
rect 10725 24197 10811 24253
rect 10867 24197 10953 24253
rect 11009 24197 11095 24253
rect 11151 24197 11237 24253
rect 11293 24197 11379 24253
rect 11435 24197 11521 24253
rect 11577 24197 11663 24253
rect 11719 24197 11805 24253
rect 11861 24197 11947 24253
rect 12003 24197 12089 24253
rect 12145 24197 12231 24253
rect 12287 24197 12373 24253
rect 12429 24197 12515 24253
rect 12571 24197 12657 24253
rect 12713 24197 12799 24253
rect 12855 24197 12941 24253
rect 12997 24197 13083 24253
rect 13139 24197 13225 24253
rect 13281 24197 13367 24253
rect 13423 24197 13509 24253
rect 13565 24197 13651 24253
rect 13707 24197 13793 24253
rect 13849 24197 13935 24253
rect 13991 24197 14077 24253
rect 14133 24197 14219 24253
rect 14275 24197 14361 24253
rect 14417 24197 14503 24253
rect 14559 24197 14645 24253
rect 14701 24197 14787 24253
rect 14843 24197 15000 24253
rect 0 24111 15000 24197
rect 0 24055 161 24111
rect 217 24055 303 24111
rect 359 24055 445 24111
rect 501 24055 587 24111
rect 643 24055 729 24111
rect 785 24055 871 24111
rect 927 24055 1013 24111
rect 1069 24055 1155 24111
rect 1211 24055 1297 24111
rect 1353 24055 1439 24111
rect 1495 24055 1581 24111
rect 1637 24055 1723 24111
rect 1779 24055 1865 24111
rect 1921 24055 2007 24111
rect 2063 24055 2149 24111
rect 2205 24055 2291 24111
rect 2347 24055 2433 24111
rect 2489 24055 2575 24111
rect 2631 24055 2717 24111
rect 2773 24055 2859 24111
rect 2915 24055 3001 24111
rect 3057 24055 3143 24111
rect 3199 24055 3285 24111
rect 3341 24055 3427 24111
rect 3483 24055 3569 24111
rect 3625 24055 3711 24111
rect 3767 24055 3853 24111
rect 3909 24055 3995 24111
rect 4051 24055 4137 24111
rect 4193 24055 4279 24111
rect 4335 24055 4421 24111
rect 4477 24055 4563 24111
rect 4619 24055 4705 24111
rect 4761 24055 4847 24111
rect 4903 24055 4989 24111
rect 5045 24055 5131 24111
rect 5187 24055 5273 24111
rect 5329 24055 5415 24111
rect 5471 24055 5557 24111
rect 5613 24055 5699 24111
rect 5755 24055 5841 24111
rect 5897 24055 5983 24111
rect 6039 24055 6125 24111
rect 6181 24055 6267 24111
rect 6323 24055 6409 24111
rect 6465 24055 6551 24111
rect 6607 24055 6693 24111
rect 6749 24055 6835 24111
rect 6891 24055 6977 24111
rect 7033 24055 7119 24111
rect 7175 24055 7261 24111
rect 7317 24055 7403 24111
rect 7459 24055 7545 24111
rect 7601 24055 7687 24111
rect 7743 24055 7829 24111
rect 7885 24055 7971 24111
rect 8027 24055 8113 24111
rect 8169 24055 8255 24111
rect 8311 24055 8397 24111
rect 8453 24055 8539 24111
rect 8595 24055 8681 24111
rect 8737 24055 8823 24111
rect 8879 24055 8965 24111
rect 9021 24055 9107 24111
rect 9163 24055 9249 24111
rect 9305 24055 9391 24111
rect 9447 24055 9533 24111
rect 9589 24055 9675 24111
rect 9731 24055 9817 24111
rect 9873 24055 9959 24111
rect 10015 24055 10101 24111
rect 10157 24055 10243 24111
rect 10299 24055 10385 24111
rect 10441 24055 10527 24111
rect 10583 24055 10669 24111
rect 10725 24055 10811 24111
rect 10867 24055 10953 24111
rect 11009 24055 11095 24111
rect 11151 24055 11237 24111
rect 11293 24055 11379 24111
rect 11435 24055 11521 24111
rect 11577 24055 11663 24111
rect 11719 24055 11805 24111
rect 11861 24055 11947 24111
rect 12003 24055 12089 24111
rect 12145 24055 12231 24111
rect 12287 24055 12373 24111
rect 12429 24055 12515 24111
rect 12571 24055 12657 24111
rect 12713 24055 12799 24111
rect 12855 24055 12941 24111
rect 12997 24055 13083 24111
rect 13139 24055 13225 24111
rect 13281 24055 13367 24111
rect 13423 24055 13509 24111
rect 13565 24055 13651 24111
rect 13707 24055 13793 24111
rect 13849 24055 13935 24111
rect 13991 24055 14077 24111
rect 14133 24055 14219 24111
rect 14275 24055 14361 24111
rect 14417 24055 14503 24111
rect 14559 24055 14645 24111
rect 14701 24055 14787 24111
rect 14843 24055 15000 24111
rect 0 23969 15000 24055
rect 0 23913 161 23969
rect 217 23913 303 23969
rect 359 23913 445 23969
rect 501 23913 587 23969
rect 643 23913 729 23969
rect 785 23913 871 23969
rect 927 23913 1013 23969
rect 1069 23913 1155 23969
rect 1211 23913 1297 23969
rect 1353 23913 1439 23969
rect 1495 23913 1581 23969
rect 1637 23913 1723 23969
rect 1779 23913 1865 23969
rect 1921 23913 2007 23969
rect 2063 23913 2149 23969
rect 2205 23913 2291 23969
rect 2347 23913 2433 23969
rect 2489 23913 2575 23969
rect 2631 23913 2717 23969
rect 2773 23913 2859 23969
rect 2915 23913 3001 23969
rect 3057 23913 3143 23969
rect 3199 23913 3285 23969
rect 3341 23913 3427 23969
rect 3483 23913 3569 23969
rect 3625 23913 3711 23969
rect 3767 23913 3853 23969
rect 3909 23913 3995 23969
rect 4051 23913 4137 23969
rect 4193 23913 4279 23969
rect 4335 23913 4421 23969
rect 4477 23913 4563 23969
rect 4619 23913 4705 23969
rect 4761 23913 4847 23969
rect 4903 23913 4989 23969
rect 5045 23913 5131 23969
rect 5187 23913 5273 23969
rect 5329 23913 5415 23969
rect 5471 23913 5557 23969
rect 5613 23913 5699 23969
rect 5755 23913 5841 23969
rect 5897 23913 5983 23969
rect 6039 23913 6125 23969
rect 6181 23913 6267 23969
rect 6323 23913 6409 23969
rect 6465 23913 6551 23969
rect 6607 23913 6693 23969
rect 6749 23913 6835 23969
rect 6891 23913 6977 23969
rect 7033 23913 7119 23969
rect 7175 23913 7261 23969
rect 7317 23913 7403 23969
rect 7459 23913 7545 23969
rect 7601 23913 7687 23969
rect 7743 23913 7829 23969
rect 7885 23913 7971 23969
rect 8027 23913 8113 23969
rect 8169 23913 8255 23969
rect 8311 23913 8397 23969
rect 8453 23913 8539 23969
rect 8595 23913 8681 23969
rect 8737 23913 8823 23969
rect 8879 23913 8965 23969
rect 9021 23913 9107 23969
rect 9163 23913 9249 23969
rect 9305 23913 9391 23969
rect 9447 23913 9533 23969
rect 9589 23913 9675 23969
rect 9731 23913 9817 23969
rect 9873 23913 9959 23969
rect 10015 23913 10101 23969
rect 10157 23913 10243 23969
rect 10299 23913 10385 23969
rect 10441 23913 10527 23969
rect 10583 23913 10669 23969
rect 10725 23913 10811 23969
rect 10867 23913 10953 23969
rect 11009 23913 11095 23969
rect 11151 23913 11237 23969
rect 11293 23913 11379 23969
rect 11435 23913 11521 23969
rect 11577 23913 11663 23969
rect 11719 23913 11805 23969
rect 11861 23913 11947 23969
rect 12003 23913 12089 23969
rect 12145 23913 12231 23969
rect 12287 23913 12373 23969
rect 12429 23913 12515 23969
rect 12571 23913 12657 23969
rect 12713 23913 12799 23969
rect 12855 23913 12941 23969
rect 12997 23913 13083 23969
rect 13139 23913 13225 23969
rect 13281 23913 13367 23969
rect 13423 23913 13509 23969
rect 13565 23913 13651 23969
rect 13707 23913 13793 23969
rect 13849 23913 13935 23969
rect 13991 23913 14077 23969
rect 14133 23913 14219 23969
rect 14275 23913 14361 23969
rect 14417 23913 14503 23969
rect 14559 23913 14645 23969
rect 14701 23913 14787 23969
rect 14843 23913 15000 23969
rect 0 23827 15000 23913
rect 0 23771 161 23827
rect 217 23771 303 23827
rect 359 23771 445 23827
rect 501 23771 587 23827
rect 643 23771 729 23827
rect 785 23771 871 23827
rect 927 23771 1013 23827
rect 1069 23771 1155 23827
rect 1211 23771 1297 23827
rect 1353 23771 1439 23827
rect 1495 23771 1581 23827
rect 1637 23771 1723 23827
rect 1779 23771 1865 23827
rect 1921 23771 2007 23827
rect 2063 23771 2149 23827
rect 2205 23771 2291 23827
rect 2347 23771 2433 23827
rect 2489 23771 2575 23827
rect 2631 23771 2717 23827
rect 2773 23771 2859 23827
rect 2915 23771 3001 23827
rect 3057 23771 3143 23827
rect 3199 23771 3285 23827
rect 3341 23771 3427 23827
rect 3483 23771 3569 23827
rect 3625 23771 3711 23827
rect 3767 23771 3853 23827
rect 3909 23771 3995 23827
rect 4051 23771 4137 23827
rect 4193 23771 4279 23827
rect 4335 23771 4421 23827
rect 4477 23771 4563 23827
rect 4619 23771 4705 23827
rect 4761 23771 4847 23827
rect 4903 23771 4989 23827
rect 5045 23771 5131 23827
rect 5187 23771 5273 23827
rect 5329 23771 5415 23827
rect 5471 23771 5557 23827
rect 5613 23771 5699 23827
rect 5755 23771 5841 23827
rect 5897 23771 5983 23827
rect 6039 23771 6125 23827
rect 6181 23771 6267 23827
rect 6323 23771 6409 23827
rect 6465 23771 6551 23827
rect 6607 23771 6693 23827
rect 6749 23771 6835 23827
rect 6891 23771 6977 23827
rect 7033 23771 7119 23827
rect 7175 23771 7261 23827
rect 7317 23771 7403 23827
rect 7459 23771 7545 23827
rect 7601 23771 7687 23827
rect 7743 23771 7829 23827
rect 7885 23771 7971 23827
rect 8027 23771 8113 23827
rect 8169 23771 8255 23827
rect 8311 23771 8397 23827
rect 8453 23771 8539 23827
rect 8595 23771 8681 23827
rect 8737 23771 8823 23827
rect 8879 23771 8965 23827
rect 9021 23771 9107 23827
rect 9163 23771 9249 23827
rect 9305 23771 9391 23827
rect 9447 23771 9533 23827
rect 9589 23771 9675 23827
rect 9731 23771 9817 23827
rect 9873 23771 9959 23827
rect 10015 23771 10101 23827
rect 10157 23771 10243 23827
rect 10299 23771 10385 23827
rect 10441 23771 10527 23827
rect 10583 23771 10669 23827
rect 10725 23771 10811 23827
rect 10867 23771 10953 23827
rect 11009 23771 11095 23827
rect 11151 23771 11237 23827
rect 11293 23771 11379 23827
rect 11435 23771 11521 23827
rect 11577 23771 11663 23827
rect 11719 23771 11805 23827
rect 11861 23771 11947 23827
rect 12003 23771 12089 23827
rect 12145 23771 12231 23827
rect 12287 23771 12373 23827
rect 12429 23771 12515 23827
rect 12571 23771 12657 23827
rect 12713 23771 12799 23827
rect 12855 23771 12941 23827
rect 12997 23771 13083 23827
rect 13139 23771 13225 23827
rect 13281 23771 13367 23827
rect 13423 23771 13509 23827
rect 13565 23771 13651 23827
rect 13707 23771 13793 23827
rect 13849 23771 13935 23827
rect 13991 23771 14077 23827
rect 14133 23771 14219 23827
rect 14275 23771 14361 23827
rect 14417 23771 14503 23827
rect 14559 23771 14645 23827
rect 14701 23771 14787 23827
rect 14843 23771 15000 23827
rect 0 23685 15000 23771
rect 0 23629 161 23685
rect 217 23629 303 23685
rect 359 23629 445 23685
rect 501 23629 587 23685
rect 643 23629 729 23685
rect 785 23629 871 23685
rect 927 23629 1013 23685
rect 1069 23629 1155 23685
rect 1211 23629 1297 23685
rect 1353 23629 1439 23685
rect 1495 23629 1581 23685
rect 1637 23629 1723 23685
rect 1779 23629 1865 23685
rect 1921 23629 2007 23685
rect 2063 23629 2149 23685
rect 2205 23629 2291 23685
rect 2347 23629 2433 23685
rect 2489 23629 2575 23685
rect 2631 23629 2717 23685
rect 2773 23629 2859 23685
rect 2915 23629 3001 23685
rect 3057 23629 3143 23685
rect 3199 23629 3285 23685
rect 3341 23629 3427 23685
rect 3483 23629 3569 23685
rect 3625 23629 3711 23685
rect 3767 23629 3853 23685
rect 3909 23629 3995 23685
rect 4051 23629 4137 23685
rect 4193 23629 4279 23685
rect 4335 23629 4421 23685
rect 4477 23629 4563 23685
rect 4619 23629 4705 23685
rect 4761 23629 4847 23685
rect 4903 23629 4989 23685
rect 5045 23629 5131 23685
rect 5187 23629 5273 23685
rect 5329 23629 5415 23685
rect 5471 23629 5557 23685
rect 5613 23629 5699 23685
rect 5755 23629 5841 23685
rect 5897 23629 5983 23685
rect 6039 23629 6125 23685
rect 6181 23629 6267 23685
rect 6323 23629 6409 23685
rect 6465 23629 6551 23685
rect 6607 23629 6693 23685
rect 6749 23629 6835 23685
rect 6891 23629 6977 23685
rect 7033 23629 7119 23685
rect 7175 23629 7261 23685
rect 7317 23629 7403 23685
rect 7459 23629 7545 23685
rect 7601 23629 7687 23685
rect 7743 23629 7829 23685
rect 7885 23629 7971 23685
rect 8027 23629 8113 23685
rect 8169 23629 8255 23685
rect 8311 23629 8397 23685
rect 8453 23629 8539 23685
rect 8595 23629 8681 23685
rect 8737 23629 8823 23685
rect 8879 23629 8965 23685
rect 9021 23629 9107 23685
rect 9163 23629 9249 23685
rect 9305 23629 9391 23685
rect 9447 23629 9533 23685
rect 9589 23629 9675 23685
rect 9731 23629 9817 23685
rect 9873 23629 9959 23685
rect 10015 23629 10101 23685
rect 10157 23629 10243 23685
rect 10299 23629 10385 23685
rect 10441 23629 10527 23685
rect 10583 23629 10669 23685
rect 10725 23629 10811 23685
rect 10867 23629 10953 23685
rect 11009 23629 11095 23685
rect 11151 23629 11237 23685
rect 11293 23629 11379 23685
rect 11435 23629 11521 23685
rect 11577 23629 11663 23685
rect 11719 23629 11805 23685
rect 11861 23629 11947 23685
rect 12003 23629 12089 23685
rect 12145 23629 12231 23685
rect 12287 23629 12373 23685
rect 12429 23629 12515 23685
rect 12571 23629 12657 23685
rect 12713 23629 12799 23685
rect 12855 23629 12941 23685
rect 12997 23629 13083 23685
rect 13139 23629 13225 23685
rect 13281 23629 13367 23685
rect 13423 23629 13509 23685
rect 13565 23629 13651 23685
rect 13707 23629 13793 23685
rect 13849 23629 13935 23685
rect 13991 23629 14077 23685
rect 14133 23629 14219 23685
rect 14275 23629 14361 23685
rect 14417 23629 14503 23685
rect 14559 23629 14645 23685
rect 14701 23629 14787 23685
rect 14843 23629 15000 23685
rect 0 23600 15000 23629
rect 0 23341 15000 23400
rect 0 23285 161 23341
rect 217 23285 303 23341
rect 359 23285 445 23341
rect 501 23285 587 23341
rect 643 23285 729 23341
rect 785 23285 871 23341
rect 927 23285 1013 23341
rect 1069 23285 1155 23341
rect 1211 23285 1297 23341
rect 1353 23285 1439 23341
rect 1495 23285 1581 23341
rect 1637 23285 1723 23341
rect 1779 23285 1865 23341
rect 1921 23285 2007 23341
rect 2063 23285 2149 23341
rect 2205 23285 2291 23341
rect 2347 23285 2433 23341
rect 2489 23285 2575 23341
rect 2631 23285 2717 23341
rect 2773 23285 2859 23341
rect 2915 23285 3001 23341
rect 3057 23285 3143 23341
rect 3199 23285 3285 23341
rect 3341 23285 3427 23341
rect 3483 23285 3569 23341
rect 3625 23285 3711 23341
rect 3767 23285 3853 23341
rect 3909 23285 3995 23341
rect 4051 23285 4137 23341
rect 4193 23285 4279 23341
rect 4335 23285 4421 23341
rect 4477 23285 4563 23341
rect 4619 23285 4705 23341
rect 4761 23285 4847 23341
rect 4903 23285 4989 23341
rect 5045 23285 5131 23341
rect 5187 23285 5273 23341
rect 5329 23285 5415 23341
rect 5471 23285 5557 23341
rect 5613 23285 5699 23341
rect 5755 23285 5841 23341
rect 5897 23285 5983 23341
rect 6039 23285 6125 23341
rect 6181 23285 6267 23341
rect 6323 23285 6409 23341
rect 6465 23285 6551 23341
rect 6607 23285 6693 23341
rect 6749 23285 6835 23341
rect 6891 23285 6977 23341
rect 7033 23285 7119 23341
rect 7175 23285 7261 23341
rect 7317 23285 7403 23341
rect 7459 23285 7545 23341
rect 7601 23285 7687 23341
rect 7743 23285 7829 23341
rect 7885 23285 7971 23341
rect 8027 23285 8113 23341
rect 8169 23285 8255 23341
rect 8311 23285 8397 23341
rect 8453 23285 8539 23341
rect 8595 23285 8681 23341
rect 8737 23285 8823 23341
rect 8879 23285 8965 23341
rect 9021 23285 9107 23341
rect 9163 23285 9249 23341
rect 9305 23285 9391 23341
rect 9447 23285 9533 23341
rect 9589 23285 9675 23341
rect 9731 23285 9817 23341
rect 9873 23285 9959 23341
rect 10015 23285 10101 23341
rect 10157 23285 10243 23341
rect 10299 23285 10385 23341
rect 10441 23285 10527 23341
rect 10583 23285 10669 23341
rect 10725 23285 10811 23341
rect 10867 23285 10953 23341
rect 11009 23285 11095 23341
rect 11151 23285 11237 23341
rect 11293 23285 11379 23341
rect 11435 23285 11521 23341
rect 11577 23285 11663 23341
rect 11719 23285 11805 23341
rect 11861 23285 11947 23341
rect 12003 23285 12089 23341
rect 12145 23285 12231 23341
rect 12287 23285 12373 23341
rect 12429 23285 12515 23341
rect 12571 23285 12657 23341
rect 12713 23285 12799 23341
rect 12855 23285 12941 23341
rect 12997 23285 13083 23341
rect 13139 23285 13225 23341
rect 13281 23285 13367 23341
rect 13423 23285 13509 23341
rect 13565 23285 13651 23341
rect 13707 23285 13793 23341
rect 13849 23285 13935 23341
rect 13991 23285 14077 23341
rect 14133 23285 14219 23341
rect 14275 23285 14361 23341
rect 14417 23285 14503 23341
rect 14559 23285 14645 23341
rect 14701 23285 14787 23341
rect 14843 23285 15000 23341
rect 0 23199 15000 23285
rect 0 23143 161 23199
rect 217 23143 303 23199
rect 359 23143 445 23199
rect 501 23143 587 23199
rect 643 23143 729 23199
rect 785 23143 871 23199
rect 927 23143 1013 23199
rect 1069 23143 1155 23199
rect 1211 23143 1297 23199
rect 1353 23143 1439 23199
rect 1495 23143 1581 23199
rect 1637 23143 1723 23199
rect 1779 23143 1865 23199
rect 1921 23143 2007 23199
rect 2063 23143 2149 23199
rect 2205 23143 2291 23199
rect 2347 23143 2433 23199
rect 2489 23143 2575 23199
rect 2631 23143 2717 23199
rect 2773 23143 2859 23199
rect 2915 23143 3001 23199
rect 3057 23143 3143 23199
rect 3199 23143 3285 23199
rect 3341 23143 3427 23199
rect 3483 23143 3569 23199
rect 3625 23143 3711 23199
rect 3767 23143 3853 23199
rect 3909 23143 3995 23199
rect 4051 23143 4137 23199
rect 4193 23143 4279 23199
rect 4335 23143 4421 23199
rect 4477 23143 4563 23199
rect 4619 23143 4705 23199
rect 4761 23143 4847 23199
rect 4903 23143 4989 23199
rect 5045 23143 5131 23199
rect 5187 23143 5273 23199
rect 5329 23143 5415 23199
rect 5471 23143 5557 23199
rect 5613 23143 5699 23199
rect 5755 23143 5841 23199
rect 5897 23143 5983 23199
rect 6039 23143 6125 23199
rect 6181 23143 6267 23199
rect 6323 23143 6409 23199
rect 6465 23143 6551 23199
rect 6607 23143 6693 23199
rect 6749 23143 6835 23199
rect 6891 23143 6977 23199
rect 7033 23143 7119 23199
rect 7175 23143 7261 23199
rect 7317 23143 7403 23199
rect 7459 23143 7545 23199
rect 7601 23143 7687 23199
rect 7743 23143 7829 23199
rect 7885 23143 7971 23199
rect 8027 23143 8113 23199
rect 8169 23143 8255 23199
rect 8311 23143 8397 23199
rect 8453 23143 8539 23199
rect 8595 23143 8681 23199
rect 8737 23143 8823 23199
rect 8879 23143 8965 23199
rect 9021 23143 9107 23199
rect 9163 23143 9249 23199
rect 9305 23143 9391 23199
rect 9447 23143 9533 23199
rect 9589 23143 9675 23199
rect 9731 23143 9817 23199
rect 9873 23143 9959 23199
rect 10015 23143 10101 23199
rect 10157 23143 10243 23199
rect 10299 23143 10385 23199
rect 10441 23143 10527 23199
rect 10583 23143 10669 23199
rect 10725 23143 10811 23199
rect 10867 23143 10953 23199
rect 11009 23143 11095 23199
rect 11151 23143 11237 23199
rect 11293 23143 11379 23199
rect 11435 23143 11521 23199
rect 11577 23143 11663 23199
rect 11719 23143 11805 23199
rect 11861 23143 11947 23199
rect 12003 23143 12089 23199
rect 12145 23143 12231 23199
rect 12287 23143 12373 23199
rect 12429 23143 12515 23199
rect 12571 23143 12657 23199
rect 12713 23143 12799 23199
rect 12855 23143 12941 23199
rect 12997 23143 13083 23199
rect 13139 23143 13225 23199
rect 13281 23143 13367 23199
rect 13423 23143 13509 23199
rect 13565 23143 13651 23199
rect 13707 23143 13793 23199
rect 13849 23143 13935 23199
rect 13991 23143 14077 23199
rect 14133 23143 14219 23199
rect 14275 23143 14361 23199
rect 14417 23143 14503 23199
rect 14559 23143 14645 23199
rect 14701 23143 14787 23199
rect 14843 23143 15000 23199
rect 0 23057 15000 23143
rect 0 23001 161 23057
rect 217 23001 303 23057
rect 359 23001 445 23057
rect 501 23001 587 23057
rect 643 23001 729 23057
rect 785 23001 871 23057
rect 927 23001 1013 23057
rect 1069 23001 1155 23057
rect 1211 23001 1297 23057
rect 1353 23001 1439 23057
rect 1495 23001 1581 23057
rect 1637 23001 1723 23057
rect 1779 23001 1865 23057
rect 1921 23001 2007 23057
rect 2063 23001 2149 23057
rect 2205 23001 2291 23057
rect 2347 23001 2433 23057
rect 2489 23001 2575 23057
rect 2631 23001 2717 23057
rect 2773 23001 2859 23057
rect 2915 23001 3001 23057
rect 3057 23001 3143 23057
rect 3199 23001 3285 23057
rect 3341 23001 3427 23057
rect 3483 23001 3569 23057
rect 3625 23001 3711 23057
rect 3767 23001 3853 23057
rect 3909 23001 3995 23057
rect 4051 23001 4137 23057
rect 4193 23001 4279 23057
rect 4335 23001 4421 23057
rect 4477 23001 4563 23057
rect 4619 23001 4705 23057
rect 4761 23001 4847 23057
rect 4903 23001 4989 23057
rect 5045 23001 5131 23057
rect 5187 23001 5273 23057
rect 5329 23001 5415 23057
rect 5471 23001 5557 23057
rect 5613 23001 5699 23057
rect 5755 23001 5841 23057
rect 5897 23001 5983 23057
rect 6039 23001 6125 23057
rect 6181 23001 6267 23057
rect 6323 23001 6409 23057
rect 6465 23001 6551 23057
rect 6607 23001 6693 23057
rect 6749 23001 6835 23057
rect 6891 23001 6977 23057
rect 7033 23001 7119 23057
rect 7175 23001 7261 23057
rect 7317 23001 7403 23057
rect 7459 23001 7545 23057
rect 7601 23001 7687 23057
rect 7743 23001 7829 23057
rect 7885 23001 7971 23057
rect 8027 23001 8113 23057
rect 8169 23001 8255 23057
rect 8311 23001 8397 23057
rect 8453 23001 8539 23057
rect 8595 23001 8681 23057
rect 8737 23001 8823 23057
rect 8879 23001 8965 23057
rect 9021 23001 9107 23057
rect 9163 23001 9249 23057
rect 9305 23001 9391 23057
rect 9447 23001 9533 23057
rect 9589 23001 9675 23057
rect 9731 23001 9817 23057
rect 9873 23001 9959 23057
rect 10015 23001 10101 23057
rect 10157 23001 10243 23057
rect 10299 23001 10385 23057
rect 10441 23001 10527 23057
rect 10583 23001 10669 23057
rect 10725 23001 10811 23057
rect 10867 23001 10953 23057
rect 11009 23001 11095 23057
rect 11151 23001 11237 23057
rect 11293 23001 11379 23057
rect 11435 23001 11521 23057
rect 11577 23001 11663 23057
rect 11719 23001 11805 23057
rect 11861 23001 11947 23057
rect 12003 23001 12089 23057
rect 12145 23001 12231 23057
rect 12287 23001 12373 23057
rect 12429 23001 12515 23057
rect 12571 23001 12657 23057
rect 12713 23001 12799 23057
rect 12855 23001 12941 23057
rect 12997 23001 13083 23057
rect 13139 23001 13225 23057
rect 13281 23001 13367 23057
rect 13423 23001 13509 23057
rect 13565 23001 13651 23057
rect 13707 23001 13793 23057
rect 13849 23001 13935 23057
rect 13991 23001 14077 23057
rect 14133 23001 14219 23057
rect 14275 23001 14361 23057
rect 14417 23001 14503 23057
rect 14559 23001 14645 23057
rect 14701 23001 14787 23057
rect 14843 23001 15000 23057
rect 0 22915 15000 23001
rect 0 22859 161 22915
rect 217 22859 303 22915
rect 359 22859 445 22915
rect 501 22859 587 22915
rect 643 22859 729 22915
rect 785 22859 871 22915
rect 927 22859 1013 22915
rect 1069 22859 1155 22915
rect 1211 22859 1297 22915
rect 1353 22859 1439 22915
rect 1495 22859 1581 22915
rect 1637 22859 1723 22915
rect 1779 22859 1865 22915
rect 1921 22859 2007 22915
rect 2063 22859 2149 22915
rect 2205 22859 2291 22915
rect 2347 22859 2433 22915
rect 2489 22859 2575 22915
rect 2631 22859 2717 22915
rect 2773 22859 2859 22915
rect 2915 22859 3001 22915
rect 3057 22859 3143 22915
rect 3199 22859 3285 22915
rect 3341 22859 3427 22915
rect 3483 22859 3569 22915
rect 3625 22859 3711 22915
rect 3767 22859 3853 22915
rect 3909 22859 3995 22915
rect 4051 22859 4137 22915
rect 4193 22859 4279 22915
rect 4335 22859 4421 22915
rect 4477 22859 4563 22915
rect 4619 22859 4705 22915
rect 4761 22859 4847 22915
rect 4903 22859 4989 22915
rect 5045 22859 5131 22915
rect 5187 22859 5273 22915
rect 5329 22859 5415 22915
rect 5471 22859 5557 22915
rect 5613 22859 5699 22915
rect 5755 22859 5841 22915
rect 5897 22859 5983 22915
rect 6039 22859 6125 22915
rect 6181 22859 6267 22915
rect 6323 22859 6409 22915
rect 6465 22859 6551 22915
rect 6607 22859 6693 22915
rect 6749 22859 6835 22915
rect 6891 22859 6977 22915
rect 7033 22859 7119 22915
rect 7175 22859 7261 22915
rect 7317 22859 7403 22915
rect 7459 22859 7545 22915
rect 7601 22859 7687 22915
rect 7743 22859 7829 22915
rect 7885 22859 7971 22915
rect 8027 22859 8113 22915
rect 8169 22859 8255 22915
rect 8311 22859 8397 22915
rect 8453 22859 8539 22915
rect 8595 22859 8681 22915
rect 8737 22859 8823 22915
rect 8879 22859 8965 22915
rect 9021 22859 9107 22915
rect 9163 22859 9249 22915
rect 9305 22859 9391 22915
rect 9447 22859 9533 22915
rect 9589 22859 9675 22915
rect 9731 22859 9817 22915
rect 9873 22859 9959 22915
rect 10015 22859 10101 22915
rect 10157 22859 10243 22915
rect 10299 22859 10385 22915
rect 10441 22859 10527 22915
rect 10583 22859 10669 22915
rect 10725 22859 10811 22915
rect 10867 22859 10953 22915
rect 11009 22859 11095 22915
rect 11151 22859 11237 22915
rect 11293 22859 11379 22915
rect 11435 22859 11521 22915
rect 11577 22859 11663 22915
rect 11719 22859 11805 22915
rect 11861 22859 11947 22915
rect 12003 22859 12089 22915
rect 12145 22859 12231 22915
rect 12287 22859 12373 22915
rect 12429 22859 12515 22915
rect 12571 22859 12657 22915
rect 12713 22859 12799 22915
rect 12855 22859 12941 22915
rect 12997 22859 13083 22915
rect 13139 22859 13225 22915
rect 13281 22859 13367 22915
rect 13423 22859 13509 22915
rect 13565 22859 13651 22915
rect 13707 22859 13793 22915
rect 13849 22859 13935 22915
rect 13991 22859 14077 22915
rect 14133 22859 14219 22915
rect 14275 22859 14361 22915
rect 14417 22859 14503 22915
rect 14559 22859 14645 22915
rect 14701 22859 14787 22915
rect 14843 22859 15000 22915
rect 0 22773 15000 22859
rect 0 22717 161 22773
rect 217 22717 303 22773
rect 359 22717 445 22773
rect 501 22717 587 22773
rect 643 22717 729 22773
rect 785 22717 871 22773
rect 927 22717 1013 22773
rect 1069 22717 1155 22773
rect 1211 22717 1297 22773
rect 1353 22717 1439 22773
rect 1495 22717 1581 22773
rect 1637 22717 1723 22773
rect 1779 22717 1865 22773
rect 1921 22717 2007 22773
rect 2063 22717 2149 22773
rect 2205 22717 2291 22773
rect 2347 22717 2433 22773
rect 2489 22717 2575 22773
rect 2631 22717 2717 22773
rect 2773 22717 2859 22773
rect 2915 22717 3001 22773
rect 3057 22717 3143 22773
rect 3199 22717 3285 22773
rect 3341 22717 3427 22773
rect 3483 22717 3569 22773
rect 3625 22717 3711 22773
rect 3767 22717 3853 22773
rect 3909 22717 3995 22773
rect 4051 22717 4137 22773
rect 4193 22717 4279 22773
rect 4335 22717 4421 22773
rect 4477 22717 4563 22773
rect 4619 22717 4705 22773
rect 4761 22717 4847 22773
rect 4903 22717 4989 22773
rect 5045 22717 5131 22773
rect 5187 22717 5273 22773
rect 5329 22717 5415 22773
rect 5471 22717 5557 22773
rect 5613 22717 5699 22773
rect 5755 22717 5841 22773
rect 5897 22717 5983 22773
rect 6039 22717 6125 22773
rect 6181 22717 6267 22773
rect 6323 22717 6409 22773
rect 6465 22717 6551 22773
rect 6607 22717 6693 22773
rect 6749 22717 6835 22773
rect 6891 22717 6977 22773
rect 7033 22717 7119 22773
rect 7175 22717 7261 22773
rect 7317 22717 7403 22773
rect 7459 22717 7545 22773
rect 7601 22717 7687 22773
rect 7743 22717 7829 22773
rect 7885 22717 7971 22773
rect 8027 22717 8113 22773
rect 8169 22717 8255 22773
rect 8311 22717 8397 22773
rect 8453 22717 8539 22773
rect 8595 22717 8681 22773
rect 8737 22717 8823 22773
rect 8879 22717 8965 22773
rect 9021 22717 9107 22773
rect 9163 22717 9249 22773
rect 9305 22717 9391 22773
rect 9447 22717 9533 22773
rect 9589 22717 9675 22773
rect 9731 22717 9817 22773
rect 9873 22717 9959 22773
rect 10015 22717 10101 22773
rect 10157 22717 10243 22773
rect 10299 22717 10385 22773
rect 10441 22717 10527 22773
rect 10583 22717 10669 22773
rect 10725 22717 10811 22773
rect 10867 22717 10953 22773
rect 11009 22717 11095 22773
rect 11151 22717 11237 22773
rect 11293 22717 11379 22773
rect 11435 22717 11521 22773
rect 11577 22717 11663 22773
rect 11719 22717 11805 22773
rect 11861 22717 11947 22773
rect 12003 22717 12089 22773
rect 12145 22717 12231 22773
rect 12287 22717 12373 22773
rect 12429 22717 12515 22773
rect 12571 22717 12657 22773
rect 12713 22717 12799 22773
rect 12855 22717 12941 22773
rect 12997 22717 13083 22773
rect 13139 22717 13225 22773
rect 13281 22717 13367 22773
rect 13423 22717 13509 22773
rect 13565 22717 13651 22773
rect 13707 22717 13793 22773
rect 13849 22717 13935 22773
rect 13991 22717 14077 22773
rect 14133 22717 14219 22773
rect 14275 22717 14361 22773
rect 14417 22717 14503 22773
rect 14559 22717 14645 22773
rect 14701 22717 14787 22773
rect 14843 22717 15000 22773
rect 0 22631 15000 22717
rect 0 22575 161 22631
rect 217 22575 303 22631
rect 359 22575 445 22631
rect 501 22575 587 22631
rect 643 22575 729 22631
rect 785 22575 871 22631
rect 927 22575 1013 22631
rect 1069 22575 1155 22631
rect 1211 22575 1297 22631
rect 1353 22575 1439 22631
rect 1495 22575 1581 22631
rect 1637 22575 1723 22631
rect 1779 22575 1865 22631
rect 1921 22575 2007 22631
rect 2063 22575 2149 22631
rect 2205 22575 2291 22631
rect 2347 22575 2433 22631
rect 2489 22575 2575 22631
rect 2631 22575 2717 22631
rect 2773 22575 2859 22631
rect 2915 22575 3001 22631
rect 3057 22575 3143 22631
rect 3199 22575 3285 22631
rect 3341 22575 3427 22631
rect 3483 22575 3569 22631
rect 3625 22575 3711 22631
rect 3767 22575 3853 22631
rect 3909 22575 3995 22631
rect 4051 22575 4137 22631
rect 4193 22575 4279 22631
rect 4335 22575 4421 22631
rect 4477 22575 4563 22631
rect 4619 22575 4705 22631
rect 4761 22575 4847 22631
rect 4903 22575 4989 22631
rect 5045 22575 5131 22631
rect 5187 22575 5273 22631
rect 5329 22575 5415 22631
rect 5471 22575 5557 22631
rect 5613 22575 5699 22631
rect 5755 22575 5841 22631
rect 5897 22575 5983 22631
rect 6039 22575 6125 22631
rect 6181 22575 6267 22631
rect 6323 22575 6409 22631
rect 6465 22575 6551 22631
rect 6607 22575 6693 22631
rect 6749 22575 6835 22631
rect 6891 22575 6977 22631
rect 7033 22575 7119 22631
rect 7175 22575 7261 22631
rect 7317 22575 7403 22631
rect 7459 22575 7545 22631
rect 7601 22575 7687 22631
rect 7743 22575 7829 22631
rect 7885 22575 7971 22631
rect 8027 22575 8113 22631
rect 8169 22575 8255 22631
rect 8311 22575 8397 22631
rect 8453 22575 8539 22631
rect 8595 22575 8681 22631
rect 8737 22575 8823 22631
rect 8879 22575 8965 22631
rect 9021 22575 9107 22631
rect 9163 22575 9249 22631
rect 9305 22575 9391 22631
rect 9447 22575 9533 22631
rect 9589 22575 9675 22631
rect 9731 22575 9817 22631
rect 9873 22575 9959 22631
rect 10015 22575 10101 22631
rect 10157 22575 10243 22631
rect 10299 22575 10385 22631
rect 10441 22575 10527 22631
rect 10583 22575 10669 22631
rect 10725 22575 10811 22631
rect 10867 22575 10953 22631
rect 11009 22575 11095 22631
rect 11151 22575 11237 22631
rect 11293 22575 11379 22631
rect 11435 22575 11521 22631
rect 11577 22575 11663 22631
rect 11719 22575 11805 22631
rect 11861 22575 11947 22631
rect 12003 22575 12089 22631
rect 12145 22575 12231 22631
rect 12287 22575 12373 22631
rect 12429 22575 12515 22631
rect 12571 22575 12657 22631
rect 12713 22575 12799 22631
rect 12855 22575 12941 22631
rect 12997 22575 13083 22631
rect 13139 22575 13225 22631
rect 13281 22575 13367 22631
rect 13423 22575 13509 22631
rect 13565 22575 13651 22631
rect 13707 22575 13793 22631
rect 13849 22575 13935 22631
rect 13991 22575 14077 22631
rect 14133 22575 14219 22631
rect 14275 22575 14361 22631
rect 14417 22575 14503 22631
rect 14559 22575 14645 22631
rect 14701 22575 14787 22631
rect 14843 22575 15000 22631
rect 0 22489 15000 22575
rect 0 22433 161 22489
rect 217 22433 303 22489
rect 359 22433 445 22489
rect 501 22433 587 22489
rect 643 22433 729 22489
rect 785 22433 871 22489
rect 927 22433 1013 22489
rect 1069 22433 1155 22489
rect 1211 22433 1297 22489
rect 1353 22433 1439 22489
rect 1495 22433 1581 22489
rect 1637 22433 1723 22489
rect 1779 22433 1865 22489
rect 1921 22433 2007 22489
rect 2063 22433 2149 22489
rect 2205 22433 2291 22489
rect 2347 22433 2433 22489
rect 2489 22433 2575 22489
rect 2631 22433 2717 22489
rect 2773 22433 2859 22489
rect 2915 22433 3001 22489
rect 3057 22433 3143 22489
rect 3199 22433 3285 22489
rect 3341 22433 3427 22489
rect 3483 22433 3569 22489
rect 3625 22433 3711 22489
rect 3767 22433 3853 22489
rect 3909 22433 3995 22489
rect 4051 22433 4137 22489
rect 4193 22433 4279 22489
rect 4335 22433 4421 22489
rect 4477 22433 4563 22489
rect 4619 22433 4705 22489
rect 4761 22433 4847 22489
rect 4903 22433 4989 22489
rect 5045 22433 5131 22489
rect 5187 22433 5273 22489
rect 5329 22433 5415 22489
rect 5471 22433 5557 22489
rect 5613 22433 5699 22489
rect 5755 22433 5841 22489
rect 5897 22433 5983 22489
rect 6039 22433 6125 22489
rect 6181 22433 6267 22489
rect 6323 22433 6409 22489
rect 6465 22433 6551 22489
rect 6607 22433 6693 22489
rect 6749 22433 6835 22489
rect 6891 22433 6977 22489
rect 7033 22433 7119 22489
rect 7175 22433 7261 22489
rect 7317 22433 7403 22489
rect 7459 22433 7545 22489
rect 7601 22433 7687 22489
rect 7743 22433 7829 22489
rect 7885 22433 7971 22489
rect 8027 22433 8113 22489
rect 8169 22433 8255 22489
rect 8311 22433 8397 22489
rect 8453 22433 8539 22489
rect 8595 22433 8681 22489
rect 8737 22433 8823 22489
rect 8879 22433 8965 22489
rect 9021 22433 9107 22489
rect 9163 22433 9249 22489
rect 9305 22433 9391 22489
rect 9447 22433 9533 22489
rect 9589 22433 9675 22489
rect 9731 22433 9817 22489
rect 9873 22433 9959 22489
rect 10015 22433 10101 22489
rect 10157 22433 10243 22489
rect 10299 22433 10385 22489
rect 10441 22433 10527 22489
rect 10583 22433 10669 22489
rect 10725 22433 10811 22489
rect 10867 22433 10953 22489
rect 11009 22433 11095 22489
rect 11151 22433 11237 22489
rect 11293 22433 11379 22489
rect 11435 22433 11521 22489
rect 11577 22433 11663 22489
rect 11719 22433 11805 22489
rect 11861 22433 11947 22489
rect 12003 22433 12089 22489
rect 12145 22433 12231 22489
rect 12287 22433 12373 22489
rect 12429 22433 12515 22489
rect 12571 22433 12657 22489
rect 12713 22433 12799 22489
rect 12855 22433 12941 22489
rect 12997 22433 13083 22489
rect 13139 22433 13225 22489
rect 13281 22433 13367 22489
rect 13423 22433 13509 22489
rect 13565 22433 13651 22489
rect 13707 22433 13793 22489
rect 13849 22433 13935 22489
rect 13991 22433 14077 22489
rect 14133 22433 14219 22489
rect 14275 22433 14361 22489
rect 14417 22433 14503 22489
rect 14559 22433 14645 22489
rect 14701 22433 14787 22489
rect 14843 22433 15000 22489
rect 0 22347 15000 22433
rect 0 22291 161 22347
rect 217 22291 303 22347
rect 359 22291 445 22347
rect 501 22291 587 22347
rect 643 22291 729 22347
rect 785 22291 871 22347
rect 927 22291 1013 22347
rect 1069 22291 1155 22347
rect 1211 22291 1297 22347
rect 1353 22291 1439 22347
rect 1495 22291 1581 22347
rect 1637 22291 1723 22347
rect 1779 22291 1865 22347
rect 1921 22291 2007 22347
rect 2063 22291 2149 22347
rect 2205 22291 2291 22347
rect 2347 22291 2433 22347
rect 2489 22291 2575 22347
rect 2631 22291 2717 22347
rect 2773 22291 2859 22347
rect 2915 22291 3001 22347
rect 3057 22291 3143 22347
rect 3199 22291 3285 22347
rect 3341 22291 3427 22347
rect 3483 22291 3569 22347
rect 3625 22291 3711 22347
rect 3767 22291 3853 22347
rect 3909 22291 3995 22347
rect 4051 22291 4137 22347
rect 4193 22291 4279 22347
rect 4335 22291 4421 22347
rect 4477 22291 4563 22347
rect 4619 22291 4705 22347
rect 4761 22291 4847 22347
rect 4903 22291 4989 22347
rect 5045 22291 5131 22347
rect 5187 22291 5273 22347
rect 5329 22291 5415 22347
rect 5471 22291 5557 22347
rect 5613 22291 5699 22347
rect 5755 22291 5841 22347
rect 5897 22291 5983 22347
rect 6039 22291 6125 22347
rect 6181 22291 6267 22347
rect 6323 22291 6409 22347
rect 6465 22291 6551 22347
rect 6607 22291 6693 22347
rect 6749 22291 6835 22347
rect 6891 22291 6977 22347
rect 7033 22291 7119 22347
rect 7175 22291 7261 22347
rect 7317 22291 7403 22347
rect 7459 22291 7545 22347
rect 7601 22291 7687 22347
rect 7743 22291 7829 22347
rect 7885 22291 7971 22347
rect 8027 22291 8113 22347
rect 8169 22291 8255 22347
rect 8311 22291 8397 22347
rect 8453 22291 8539 22347
rect 8595 22291 8681 22347
rect 8737 22291 8823 22347
rect 8879 22291 8965 22347
rect 9021 22291 9107 22347
rect 9163 22291 9249 22347
rect 9305 22291 9391 22347
rect 9447 22291 9533 22347
rect 9589 22291 9675 22347
rect 9731 22291 9817 22347
rect 9873 22291 9959 22347
rect 10015 22291 10101 22347
rect 10157 22291 10243 22347
rect 10299 22291 10385 22347
rect 10441 22291 10527 22347
rect 10583 22291 10669 22347
rect 10725 22291 10811 22347
rect 10867 22291 10953 22347
rect 11009 22291 11095 22347
rect 11151 22291 11237 22347
rect 11293 22291 11379 22347
rect 11435 22291 11521 22347
rect 11577 22291 11663 22347
rect 11719 22291 11805 22347
rect 11861 22291 11947 22347
rect 12003 22291 12089 22347
rect 12145 22291 12231 22347
rect 12287 22291 12373 22347
rect 12429 22291 12515 22347
rect 12571 22291 12657 22347
rect 12713 22291 12799 22347
rect 12855 22291 12941 22347
rect 12997 22291 13083 22347
rect 13139 22291 13225 22347
rect 13281 22291 13367 22347
rect 13423 22291 13509 22347
rect 13565 22291 13651 22347
rect 13707 22291 13793 22347
rect 13849 22291 13935 22347
rect 13991 22291 14077 22347
rect 14133 22291 14219 22347
rect 14275 22291 14361 22347
rect 14417 22291 14503 22347
rect 14559 22291 14645 22347
rect 14701 22291 14787 22347
rect 14843 22291 15000 22347
rect 0 22205 15000 22291
rect 0 22149 161 22205
rect 217 22149 303 22205
rect 359 22149 445 22205
rect 501 22149 587 22205
rect 643 22149 729 22205
rect 785 22149 871 22205
rect 927 22149 1013 22205
rect 1069 22149 1155 22205
rect 1211 22149 1297 22205
rect 1353 22149 1439 22205
rect 1495 22149 1581 22205
rect 1637 22149 1723 22205
rect 1779 22149 1865 22205
rect 1921 22149 2007 22205
rect 2063 22149 2149 22205
rect 2205 22149 2291 22205
rect 2347 22149 2433 22205
rect 2489 22149 2575 22205
rect 2631 22149 2717 22205
rect 2773 22149 2859 22205
rect 2915 22149 3001 22205
rect 3057 22149 3143 22205
rect 3199 22149 3285 22205
rect 3341 22149 3427 22205
rect 3483 22149 3569 22205
rect 3625 22149 3711 22205
rect 3767 22149 3853 22205
rect 3909 22149 3995 22205
rect 4051 22149 4137 22205
rect 4193 22149 4279 22205
rect 4335 22149 4421 22205
rect 4477 22149 4563 22205
rect 4619 22149 4705 22205
rect 4761 22149 4847 22205
rect 4903 22149 4989 22205
rect 5045 22149 5131 22205
rect 5187 22149 5273 22205
rect 5329 22149 5415 22205
rect 5471 22149 5557 22205
rect 5613 22149 5699 22205
rect 5755 22149 5841 22205
rect 5897 22149 5983 22205
rect 6039 22149 6125 22205
rect 6181 22149 6267 22205
rect 6323 22149 6409 22205
rect 6465 22149 6551 22205
rect 6607 22149 6693 22205
rect 6749 22149 6835 22205
rect 6891 22149 6977 22205
rect 7033 22149 7119 22205
rect 7175 22149 7261 22205
rect 7317 22149 7403 22205
rect 7459 22149 7545 22205
rect 7601 22149 7687 22205
rect 7743 22149 7829 22205
rect 7885 22149 7971 22205
rect 8027 22149 8113 22205
rect 8169 22149 8255 22205
rect 8311 22149 8397 22205
rect 8453 22149 8539 22205
rect 8595 22149 8681 22205
rect 8737 22149 8823 22205
rect 8879 22149 8965 22205
rect 9021 22149 9107 22205
rect 9163 22149 9249 22205
rect 9305 22149 9391 22205
rect 9447 22149 9533 22205
rect 9589 22149 9675 22205
rect 9731 22149 9817 22205
rect 9873 22149 9959 22205
rect 10015 22149 10101 22205
rect 10157 22149 10243 22205
rect 10299 22149 10385 22205
rect 10441 22149 10527 22205
rect 10583 22149 10669 22205
rect 10725 22149 10811 22205
rect 10867 22149 10953 22205
rect 11009 22149 11095 22205
rect 11151 22149 11237 22205
rect 11293 22149 11379 22205
rect 11435 22149 11521 22205
rect 11577 22149 11663 22205
rect 11719 22149 11805 22205
rect 11861 22149 11947 22205
rect 12003 22149 12089 22205
rect 12145 22149 12231 22205
rect 12287 22149 12373 22205
rect 12429 22149 12515 22205
rect 12571 22149 12657 22205
rect 12713 22149 12799 22205
rect 12855 22149 12941 22205
rect 12997 22149 13083 22205
rect 13139 22149 13225 22205
rect 13281 22149 13367 22205
rect 13423 22149 13509 22205
rect 13565 22149 13651 22205
rect 13707 22149 13793 22205
rect 13849 22149 13935 22205
rect 13991 22149 14077 22205
rect 14133 22149 14219 22205
rect 14275 22149 14361 22205
rect 14417 22149 14503 22205
rect 14559 22149 14645 22205
rect 14701 22149 14787 22205
rect 14843 22149 15000 22205
rect 0 22063 15000 22149
rect 0 22007 161 22063
rect 217 22007 303 22063
rect 359 22007 445 22063
rect 501 22007 587 22063
rect 643 22007 729 22063
rect 785 22007 871 22063
rect 927 22007 1013 22063
rect 1069 22007 1155 22063
rect 1211 22007 1297 22063
rect 1353 22007 1439 22063
rect 1495 22007 1581 22063
rect 1637 22007 1723 22063
rect 1779 22007 1865 22063
rect 1921 22007 2007 22063
rect 2063 22007 2149 22063
rect 2205 22007 2291 22063
rect 2347 22007 2433 22063
rect 2489 22007 2575 22063
rect 2631 22007 2717 22063
rect 2773 22007 2859 22063
rect 2915 22007 3001 22063
rect 3057 22007 3143 22063
rect 3199 22007 3285 22063
rect 3341 22007 3427 22063
rect 3483 22007 3569 22063
rect 3625 22007 3711 22063
rect 3767 22007 3853 22063
rect 3909 22007 3995 22063
rect 4051 22007 4137 22063
rect 4193 22007 4279 22063
rect 4335 22007 4421 22063
rect 4477 22007 4563 22063
rect 4619 22007 4705 22063
rect 4761 22007 4847 22063
rect 4903 22007 4989 22063
rect 5045 22007 5131 22063
rect 5187 22007 5273 22063
rect 5329 22007 5415 22063
rect 5471 22007 5557 22063
rect 5613 22007 5699 22063
rect 5755 22007 5841 22063
rect 5897 22007 5983 22063
rect 6039 22007 6125 22063
rect 6181 22007 6267 22063
rect 6323 22007 6409 22063
rect 6465 22007 6551 22063
rect 6607 22007 6693 22063
rect 6749 22007 6835 22063
rect 6891 22007 6977 22063
rect 7033 22007 7119 22063
rect 7175 22007 7261 22063
rect 7317 22007 7403 22063
rect 7459 22007 7545 22063
rect 7601 22007 7687 22063
rect 7743 22007 7829 22063
rect 7885 22007 7971 22063
rect 8027 22007 8113 22063
rect 8169 22007 8255 22063
rect 8311 22007 8397 22063
rect 8453 22007 8539 22063
rect 8595 22007 8681 22063
rect 8737 22007 8823 22063
rect 8879 22007 8965 22063
rect 9021 22007 9107 22063
rect 9163 22007 9249 22063
rect 9305 22007 9391 22063
rect 9447 22007 9533 22063
rect 9589 22007 9675 22063
rect 9731 22007 9817 22063
rect 9873 22007 9959 22063
rect 10015 22007 10101 22063
rect 10157 22007 10243 22063
rect 10299 22007 10385 22063
rect 10441 22007 10527 22063
rect 10583 22007 10669 22063
rect 10725 22007 10811 22063
rect 10867 22007 10953 22063
rect 11009 22007 11095 22063
rect 11151 22007 11237 22063
rect 11293 22007 11379 22063
rect 11435 22007 11521 22063
rect 11577 22007 11663 22063
rect 11719 22007 11805 22063
rect 11861 22007 11947 22063
rect 12003 22007 12089 22063
rect 12145 22007 12231 22063
rect 12287 22007 12373 22063
rect 12429 22007 12515 22063
rect 12571 22007 12657 22063
rect 12713 22007 12799 22063
rect 12855 22007 12941 22063
rect 12997 22007 13083 22063
rect 13139 22007 13225 22063
rect 13281 22007 13367 22063
rect 13423 22007 13509 22063
rect 13565 22007 13651 22063
rect 13707 22007 13793 22063
rect 13849 22007 13935 22063
rect 13991 22007 14077 22063
rect 14133 22007 14219 22063
rect 14275 22007 14361 22063
rect 14417 22007 14503 22063
rect 14559 22007 14645 22063
rect 14701 22007 14787 22063
rect 14843 22007 15000 22063
rect 0 21921 15000 22007
rect 0 21865 161 21921
rect 217 21865 303 21921
rect 359 21865 445 21921
rect 501 21865 587 21921
rect 643 21865 729 21921
rect 785 21865 871 21921
rect 927 21865 1013 21921
rect 1069 21865 1155 21921
rect 1211 21865 1297 21921
rect 1353 21865 1439 21921
rect 1495 21865 1581 21921
rect 1637 21865 1723 21921
rect 1779 21865 1865 21921
rect 1921 21865 2007 21921
rect 2063 21865 2149 21921
rect 2205 21865 2291 21921
rect 2347 21865 2433 21921
rect 2489 21865 2575 21921
rect 2631 21865 2717 21921
rect 2773 21865 2859 21921
rect 2915 21865 3001 21921
rect 3057 21865 3143 21921
rect 3199 21865 3285 21921
rect 3341 21865 3427 21921
rect 3483 21865 3569 21921
rect 3625 21865 3711 21921
rect 3767 21865 3853 21921
rect 3909 21865 3995 21921
rect 4051 21865 4137 21921
rect 4193 21865 4279 21921
rect 4335 21865 4421 21921
rect 4477 21865 4563 21921
rect 4619 21865 4705 21921
rect 4761 21865 4847 21921
rect 4903 21865 4989 21921
rect 5045 21865 5131 21921
rect 5187 21865 5273 21921
rect 5329 21865 5415 21921
rect 5471 21865 5557 21921
rect 5613 21865 5699 21921
rect 5755 21865 5841 21921
rect 5897 21865 5983 21921
rect 6039 21865 6125 21921
rect 6181 21865 6267 21921
rect 6323 21865 6409 21921
rect 6465 21865 6551 21921
rect 6607 21865 6693 21921
rect 6749 21865 6835 21921
rect 6891 21865 6977 21921
rect 7033 21865 7119 21921
rect 7175 21865 7261 21921
rect 7317 21865 7403 21921
rect 7459 21865 7545 21921
rect 7601 21865 7687 21921
rect 7743 21865 7829 21921
rect 7885 21865 7971 21921
rect 8027 21865 8113 21921
rect 8169 21865 8255 21921
rect 8311 21865 8397 21921
rect 8453 21865 8539 21921
rect 8595 21865 8681 21921
rect 8737 21865 8823 21921
rect 8879 21865 8965 21921
rect 9021 21865 9107 21921
rect 9163 21865 9249 21921
rect 9305 21865 9391 21921
rect 9447 21865 9533 21921
rect 9589 21865 9675 21921
rect 9731 21865 9817 21921
rect 9873 21865 9959 21921
rect 10015 21865 10101 21921
rect 10157 21865 10243 21921
rect 10299 21865 10385 21921
rect 10441 21865 10527 21921
rect 10583 21865 10669 21921
rect 10725 21865 10811 21921
rect 10867 21865 10953 21921
rect 11009 21865 11095 21921
rect 11151 21865 11237 21921
rect 11293 21865 11379 21921
rect 11435 21865 11521 21921
rect 11577 21865 11663 21921
rect 11719 21865 11805 21921
rect 11861 21865 11947 21921
rect 12003 21865 12089 21921
rect 12145 21865 12231 21921
rect 12287 21865 12373 21921
rect 12429 21865 12515 21921
rect 12571 21865 12657 21921
rect 12713 21865 12799 21921
rect 12855 21865 12941 21921
rect 12997 21865 13083 21921
rect 13139 21865 13225 21921
rect 13281 21865 13367 21921
rect 13423 21865 13509 21921
rect 13565 21865 13651 21921
rect 13707 21865 13793 21921
rect 13849 21865 13935 21921
rect 13991 21865 14077 21921
rect 14133 21865 14219 21921
rect 14275 21865 14361 21921
rect 14417 21865 14503 21921
rect 14559 21865 14645 21921
rect 14701 21865 14787 21921
rect 14843 21865 15000 21921
rect 0 21779 15000 21865
rect 0 21723 161 21779
rect 217 21723 303 21779
rect 359 21723 445 21779
rect 501 21723 587 21779
rect 643 21723 729 21779
rect 785 21723 871 21779
rect 927 21723 1013 21779
rect 1069 21723 1155 21779
rect 1211 21723 1297 21779
rect 1353 21723 1439 21779
rect 1495 21723 1581 21779
rect 1637 21723 1723 21779
rect 1779 21723 1865 21779
rect 1921 21723 2007 21779
rect 2063 21723 2149 21779
rect 2205 21723 2291 21779
rect 2347 21723 2433 21779
rect 2489 21723 2575 21779
rect 2631 21723 2717 21779
rect 2773 21723 2859 21779
rect 2915 21723 3001 21779
rect 3057 21723 3143 21779
rect 3199 21723 3285 21779
rect 3341 21723 3427 21779
rect 3483 21723 3569 21779
rect 3625 21723 3711 21779
rect 3767 21723 3853 21779
rect 3909 21723 3995 21779
rect 4051 21723 4137 21779
rect 4193 21723 4279 21779
rect 4335 21723 4421 21779
rect 4477 21723 4563 21779
rect 4619 21723 4705 21779
rect 4761 21723 4847 21779
rect 4903 21723 4989 21779
rect 5045 21723 5131 21779
rect 5187 21723 5273 21779
rect 5329 21723 5415 21779
rect 5471 21723 5557 21779
rect 5613 21723 5699 21779
rect 5755 21723 5841 21779
rect 5897 21723 5983 21779
rect 6039 21723 6125 21779
rect 6181 21723 6267 21779
rect 6323 21723 6409 21779
rect 6465 21723 6551 21779
rect 6607 21723 6693 21779
rect 6749 21723 6835 21779
rect 6891 21723 6977 21779
rect 7033 21723 7119 21779
rect 7175 21723 7261 21779
rect 7317 21723 7403 21779
rect 7459 21723 7545 21779
rect 7601 21723 7687 21779
rect 7743 21723 7829 21779
rect 7885 21723 7971 21779
rect 8027 21723 8113 21779
rect 8169 21723 8255 21779
rect 8311 21723 8397 21779
rect 8453 21723 8539 21779
rect 8595 21723 8681 21779
rect 8737 21723 8823 21779
rect 8879 21723 8965 21779
rect 9021 21723 9107 21779
rect 9163 21723 9249 21779
rect 9305 21723 9391 21779
rect 9447 21723 9533 21779
rect 9589 21723 9675 21779
rect 9731 21723 9817 21779
rect 9873 21723 9959 21779
rect 10015 21723 10101 21779
rect 10157 21723 10243 21779
rect 10299 21723 10385 21779
rect 10441 21723 10527 21779
rect 10583 21723 10669 21779
rect 10725 21723 10811 21779
rect 10867 21723 10953 21779
rect 11009 21723 11095 21779
rect 11151 21723 11237 21779
rect 11293 21723 11379 21779
rect 11435 21723 11521 21779
rect 11577 21723 11663 21779
rect 11719 21723 11805 21779
rect 11861 21723 11947 21779
rect 12003 21723 12089 21779
rect 12145 21723 12231 21779
rect 12287 21723 12373 21779
rect 12429 21723 12515 21779
rect 12571 21723 12657 21779
rect 12713 21723 12799 21779
rect 12855 21723 12941 21779
rect 12997 21723 13083 21779
rect 13139 21723 13225 21779
rect 13281 21723 13367 21779
rect 13423 21723 13509 21779
rect 13565 21723 13651 21779
rect 13707 21723 13793 21779
rect 13849 21723 13935 21779
rect 13991 21723 14077 21779
rect 14133 21723 14219 21779
rect 14275 21723 14361 21779
rect 14417 21723 14503 21779
rect 14559 21723 14645 21779
rect 14701 21723 14787 21779
rect 14843 21723 15000 21779
rect 0 21637 15000 21723
rect 0 21581 161 21637
rect 217 21581 303 21637
rect 359 21581 445 21637
rect 501 21581 587 21637
rect 643 21581 729 21637
rect 785 21581 871 21637
rect 927 21581 1013 21637
rect 1069 21581 1155 21637
rect 1211 21581 1297 21637
rect 1353 21581 1439 21637
rect 1495 21581 1581 21637
rect 1637 21581 1723 21637
rect 1779 21581 1865 21637
rect 1921 21581 2007 21637
rect 2063 21581 2149 21637
rect 2205 21581 2291 21637
rect 2347 21581 2433 21637
rect 2489 21581 2575 21637
rect 2631 21581 2717 21637
rect 2773 21581 2859 21637
rect 2915 21581 3001 21637
rect 3057 21581 3143 21637
rect 3199 21581 3285 21637
rect 3341 21581 3427 21637
rect 3483 21581 3569 21637
rect 3625 21581 3711 21637
rect 3767 21581 3853 21637
rect 3909 21581 3995 21637
rect 4051 21581 4137 21637
rect 4193 21581 4279 21637
rect 4335 21581 4421 21637
rect 4477 21581 4563 21637
rect 4619 21581 4705 21637
rect 4761 21581 4847 21637
rect 4903 21581 4989 21637
rect 5045 21581 5131 21637
rect 5187 21581 5273 21637
rect 5329 21581 5415 21637
rect 5471 21581 5557 21637
rect 5613 21581 5699 21637
rect 5755 21581 5841 21637
rect 5897 21581 5983 21637
rect 6039 21581 6125 21637
rect 6181 21581 6267 21637
rect 6323 21581 6409 21637
rect 6465 21581 6551 21637
rect 6607 21581 6693 21637
rect 6749 21581 6835 21637
rect 6891 21581 6977 21637
rect 7033 21581 7119 21637
rect 7175 21581 7261 21637
rect 7317 21581 7403 21637
rect 7459 21581 7545 21637
rect 7601 21581 7687 21637
rect 7743 21581 7829 21637
rect 7885 21581 7971 21637
rect 8027 21581 8113 21637
rect 8169 21581 8255 21637
rect 8311 21581 8397 21637
rect 8453 21581 8539 21637
rect 8595 21581 8681 21637
rect 8737 21581 8823 21637
rect 8879 21581 8965 21637
rect 9021 21581 9107 21637
rect 9163 21581 9249 21637
rect 9305 21581 9391 21637
rect 9447 21581 9533 21637
rect 9589 21581 9675 21637
rect 9731 21581 9817 21637
rect 9873 21581 9959 21637
rect 10015 21581 10101 21637
rect 10157 21581 10243 21637
rect 10299 21581 10385 21637
rect 10441 21581 10527 21637
rect 10583 21581 10669 21637
rect 10725 21581 10811 21637
rect 10867 21581 10953 21637
rect 11009 21581 11095 21637
rect 11151 21581 11237 21637
rect 11293 21581 11379 21637
rect 11435 21581 11521 21637
rect 11577 21581 11663 21637
rect 11719 21581 11805 21637
rect 11861 21581 11947 21637
rect 12003 21581 12089 21637
rect 12145 21581 12231 21637
rect 12287 21581 12373 21637
rect 12429 21581 12515 21637
rect 12571 21581 12657 21637
rect 12713 21581 12799 21637
rect 12855 21581 12941 21637
rect 12997 21581 13083 21637
rect 13139 21581 13225 21637
rect 13281 21581 13367 21637
rect 13423 21581 13509 21637
rect 13565 21581 13651 21637
rect 13707 21581 13793 21637
rect 13849 21581 13935 21637
rect 13991 21581 14077 21637
rect 14133 21581 14219 21637
rect 14275 21581 14361 21637
rect 14417 21581 14503 21637
rect 14559 21581 14645 21637
rect 14701 21581 14787 21637
rect 14843 21581 15000 21637
rect 0 21495 15000 21581
rect 0 21439 161 21495
rect 217 21439 303 21495
rect 359 21439 445 21495
rect 501 21439 587 21495
rect 643 21439 729 21495
rect 785 21439 871 21495
rect 927 21439 1013 21495
rect 1069 21439 1155 21495
rect 1211 21439 1297 21495
rect 1353 21439 1439 21495
rect 1495 21439 1581 21495
rect 1637 21439 1723 21495
rect 1779 21439 1865 21495
rect 1921 21439 2007 21495
rect 2063 21439 2149 21495
rect 2205 21439 2291 21495
rect 2347 21439 2433 21495
rect 2489 21439 2575 21495
rect 2631 21439 2717 21495
rect 2773 21439 2859 21495
rect 2915 21439 3001 21495
rect 3057 21439 3143 21495
rect 3199 21439 3285 21495
rect 3341 21439 3427 21495
rect 3483 21439 3569 21495
rect 3625 21439 3711 21495
rect 3767 21439 3853 21495
rect 3909 21439 3995 21495
rect 4051 21439 4137 21495
rect 4193 21439 4279 21495
rect 4335 21439 4421 21495
rect 4477 21439 4563 21495
rect 4619 21439 4705 21495
rect 4761 21439 4847 21495
rect 4903 21439 4989 21495
rect 5045 21439 5131 21495
rect 5187 21439 5273 21495
rect 5329 21439 5415 21495
rect 5471 21439 5557 21495
rect 5613 21439 5699 21495
rect 5755 21439 5841 21495
rect 5897 21439 5983 21495
rect 6039 21439 6125 21495
rect 6181 21439 6267 21495
rect 6323 21439 6409 21495
rect 6465 21439 6551 21495
rect 6607 21439 6693 21495
rect 6749 21439 6835 21495
rect 6891 21439 6977 21495
rect 7033 21439 7119 21495
rect 7175 21439 7261 21495
rect 7317 21439 7403 21495
rect 7459 21439 7545 21495
rect 7601 21439 7687 21495
rect 7743 21439 7829 21495
rect 7885 21439 7971 21495
rect 8027 21439 8113 21495
rect 8169 21439 8255 21495
rect 8311 21439 8397 21495
rect 8453 21439 8539 21495
rect 8595 21439 8681 21495
rect 8737 21439 8823 21495
rect 8879 21439 8965 21495
rect 9021 21439 9107 21495
rect 9163 21439 9249 21495
rect 9305 21439 9391 21495
rect 9447 21439 9533 21495
rect 9589 21439 9675 21495
rect 9731 21439 9817 21495
rect 9873 21439 9959 21495
rect 10015 21439 10101 21495
rect 10157 21439 10243 21495
rect 10299 21439 10385 21495
rect 10441 21439 10527 21495
rect 10583 21439 10669 21495
rect 10725 21439 10811 21495
rect 10867 21439 10953 21495
rect 11009 21439 11095 21495
rect 11151 21439 11237 21495
rect 11293 21439 11379 21495
rect 11435 21439 11521 21495
rect 11577 21439 11663 21495
rect 11719 21439 11805 21495
rect 11861 21439 11947 21495
rect 12003 21439 12089 21495
rect 12145 21439 12231 21495
rect 12287 21439 12373 21495
rect 12429 21439 12515 21495
rect 12571 21439 12657 21495
rect 12713 21439 12799 21495
rect 12855 21439 12941 21495
rect 12997 21439 13083 21495
rect 13139 21439 13225 21495
rect 13281 21439 13367 21495
rect 13423 21439 13509 21495
rect 13565 21439 13651 21495
rect 13707 21439 13793 21495
rect 13849 21439 13935 21495
rect 13991 21439 14077 21495
rect 14133 21439 14219 21495
rect 14275 21439 14361 21495
rect 14417 21439 14503 21495
rect 14559 21439 14645 21495
rect 14701 21439 14787 21495
rect 14843 21439 15000 21495
rect 0 21353 15000 21439
rect 0 21297 161 21353
rect 217 21297 303 21353
rect 359 21297 445 21353
rect 501 21297 587 21353
rect 643 21297 729 21353
rect 785 21297 871 21353
rect 927 21297 1013 21353
rect 1069 21297 1155 21353
rect 1211 21297 1297 21353
rect 1353 21297 1439 21353
rect 1495 21297 1581 21353
rect 1637 21297 1723 21353
rect 1779 21297 1865 21353
rect 1921 21297 2007 21353
rect 2063 21297 2149 21353
rect 2205 21297 2291 21353
rect 2347 21297 2433 21353
rect 2489 21297 2575 21353
rect 2631 21297 2717 21353
rect 2773 21297 2859 21353
rect 2915 21297 3001 21353
rect 3057 21297 3143 21353
rect 3199 21297 3285 21353
rect 3341 21297 3427 21353
rect 3483 21297 3569 21353
rect 3625 21297 3711 21353
rect 3767 21297 3853 21353
rect 3909 21297 3995 21353
rect 4051 21297 4137 21353
rect 4193 21297 4279 21353
rect 4335 21297 4421 21353
rect 4477 21297 4563 21353
rect 4619 21297 4705 21353
rect 4761 21297 4847 21353
rect 4903 21297 4989 21353
rect 5045 21297 5131 21353
rect 5187 21297 5273 21353
rect 5329 21297 5415 21353
rect 5471 21297 5557 21353
rect 5613 21297 5699 21353
rect 5755 21297 5841 21353
rect 5897 21297 5983 21353
rect 6039 21297 6125 21353
rect 6181 21297 6267 21353
rect 6323 21297 6409 21353
rect 6465 21297 6551 21353
rect 6607 21297 6693 21353
rect 6749 21297 6835 21353
rect 6891 21297 6977 21353
rect 7033 21297 7119 21353
rect 7175 21297 7261 21353
rect 7317 21297 7403 21353
rect 7459 21297 7545 21353
rect 7601 21297 7687 21353
rect 7743 21297 7829 21353
rect 7885 21297 7971 21353
rect 8027 21297 8113 21353
rect 8169 21297 8255 21353
rect 8311 21297 8397 21353
rect 8453 21297 8539 21353
rect 8595 21297 8681 21353
rect 8737 21297 8823 21353
rect 8879 21297 8965 21353
rect 9021 21297 9107 21353
rect 9163 21297 9249 21353
rect 9305 21297 9391 21353
rect 9447 21297 9533 21353
rect 9589 21297 9675 21353
rect 9731 21297 9817 21353
rect 9873 21297 9959 21353
rect 10015 21297 10101 21353
rect 10157 21297 10243 21353
rect 10299 21297 10385 21353
rect 10441 21297 10527 21353
rect 10583 21297 10669 21353
rect 10725 21297 10811 21353
rect 10867 21297 10953 21353
rect 11009 21297 11095 21353
rect 11151 21297 11237 21353
rect 11293 21297 11379 21353
rect 11435 21297 11521 21353
rect 11577 21297 11663 21353
rect 11719 21297 11805 21353
rect 11861 21297 11947 21353
rect 12003 21297 12089 21353
rect 12145 21297 12231 21353
rect 12287 21297 12373 21353
rect 12429 21297 12515 21353
rect 12571 21297 12657 21353
rect 12713 21297 12799 21353
rect 12855 21297 12941 21353
rect 12997 21297 13083 21353
rect 13139 21297 13225 21353
rect 13281 21297 13367 21353
rect 13423 21297 13509 21353
rect 13565 21297 13651 21353
rect 13707 21297 13793 21353
rect 13849 21297 13935 21353
rect 13991 21297 14077 21353
rect 14133 21297 14219 21353
rect 14275 21297 14361 21353
rect 14417 21297 14503 21353
rect 14559 21297 14645 21353
rect 14701 21297 14787 21353
rect 14843 21297 15000 21353
rect 0 21211 15000 21297
rect 0 21155 161 21211
rect 217 21155 303 21211
rect 359 21155 445 21211
rect 501 21155 587 21211
rect 643 21155 729 21211
rect 785 21155 871 21211
rect 927 21155 1013 21211
rect 1069 21155 1155 21211
rect 1211 21155 1297 21211
rect 1353 21155 1439 21211
rect 1495 21155 1581 21211
rect 1637 21155 1723 21211
rect 1779 21155 1865 21211
rect 1921 21155 2007 21211
rect 2063 21155 2149 21211
rect 2205 21155 2291 21211
rect 2347 21155 2433 21211
rect 2489 21155 2575 21211
rect 2631 21155 2717 21211
rect 2773 21155 2859 21211
rect 2915 21155 3001 21211
rect 3057 21155 3143 21211
rect 3199 21155 3285 21211
rect 3341 21155 3427 21211
rect 3483 21155 3569 21211
rect 3625 21155 3711 21211
rect 3767 21155 3853 21211
rect 3909 21155 3995 21211
rect 4051 21155 4137 21211
rect 4193 21155 4279 21211
rect 4335 21155 4421 21211
rect 4477 21155 4563 21211
rect 4619 21155 4705 21211
rect 4761 21155 4847 21211
rect 4903 21155 4989 21211
rect 5045 21155 5131 21211
rect 5187 21155 5273 21211
rect 5329 21155 5415 21211
rect 5471 21155 5557 21211
rect 5613 21155 5699 21211
rect 5755 21155 5841 21211
rect 5897 21155 5983 21211
rect 6039 21155 6125 21211
rect 6181 21155 6267 21211
rect 6323 21155 6409 21211
rect 6465 21155 6551 21211
rect 6607 21155 6693 21211
rect 6749 21155 6835 21211
rect 6891 21155 6977 21211
rect 7033 21155 7119 21211
rect 7175 21155 7261 21211
rect 7317 21155 7403 21211
rect 7459 21155 7545 21211
rect 7601 21155 7687 21211
rect 7743 21155 7829 21211
rect 7885 21155 7971 21211
rect 8027 21155 8113 21211
rect 8169 21155 8255 21211
rect 8311 21155 8397 21211
rect 8453 21155 8539 21211
rect 8595 21155 8681 21211
rect 8737 21155 8823 21211
rect 8879 21155 8965 21211
rect 9021 21155 9107 21211
rect 9163 21155 9249 21211
rect 9305 21155 9391 21211
rect 9447 21155 9533 21211
rect 9589 21155 9675 21211
rect 9731 21155 9817 21211
rect 9873 21155 9959 21211
rect 10015 21155 10101 21211
rect 10157 21155 10243 21211
rect 10299 21155 10385 21211
rect 10441 21155 10527 21211
rect 10583 21155 10669 21211
rect 10725 21155 10811 21211
rect 10867 21155 10953 21211
rect 11009 21155 11095 21211
rect 11151 21155 11237 21211
rect 11293 21155 11379 21211
rect 11435 21155 11521 21211
rect 11577 21155 11663 21211
rect 11719 21155 11805 21211
rect 11861 21155 11947 21211
rect 12003 21155 12089 21211
rect 12145 21155 12231 21211
rect 12287 21155 12373 21211
rect 12429 21155 12515 21211
rect 12571 21155 12657 21211
rect 12713 21155 12799 21211
rect 12855 21155 12941 21211
rect 12997 21155 13083 21211
rect 13139 21155 13225 21211
rect 13281 21155 13367 21211
rect 13423 21155 13509 21211
rect 13565 21155 13651 21211
rect 13707 21155 13793 21211
rect 13849 21155 13935 21211
rect 13991 21155 14077 21211
rect 14133 21155 14219 21211
rect 14275 21155 14361 21211
rect 14417 21155 14503 21211
rect 14559 21155 14645 21211
rect 14701 21155 14787 21211
rect 14843 21155 15000 21211
rect 0 21069 15000 21155
rect 0 21013 161 21069
rect 217 21013 303 21069
rect 359 21013 445 21069
rect 501 21013 587 21069
rect 643 21013 729 21069
rect 785 21013 871 21069
rect 927 21013 1013 21069
rect 1069 21013 1155 21069
rect 1211 21013 1297 21069
rect 1353 21013 1439 21069
rect 1495 21013 1581 21069
rect 1637 21013 1723 21069
rect 1779 21013 1865 21069
rect 1921 21013 2007 21069
rect 2063 21013 2149 21069
rect 2205 21013 2291 21069
rect 2347 21013 2433 21069
rect 2489 21013 2575 21069
rect 2631 21013 2717 21069
rect 2773 21013 2859 21069
rect 2915 21013 3001 21069
rect 3057 21013 3143 21069
rect 3199 21013 3285 21069
rect 3341 21013 3427 21069
rect 3483 21013 3569 21069
rect 3625 21013 3711 21069
rect 3767 21013 3853 21069
rect 3909 21013 3995 21069
rect 4051 21013 4137 21069
rect 4193 21013 4279 21069
rect 4335 21013 4421 21069
rect 4477 21013 4563 21069
rect 4619 21013 4705 21069
rect 4761 21013 4847 21069
rect 4903 21013 4989 21069
rect 5045 21013 5131 21069
rect 5187 21013 5273 21069
rect 5329 21013 5415 21069
rect 5471 21013 5557 21069
rect 5613 21013 5699 21069
rect 5755 21013 5841 21069
rect 5897 21013 5983 21069
rect 6039 21013 6125 21069
rect 6181 21013 6267 21069
rect 6323 21013 6409 21069
rect 6465 21013 6551 21069
rect 6607 21013 6693 21069
rect 6749 21013 6835 21069
rect 6891 21013 6977 21069
rect 7033 21013 7119 21069
rect 7175 21013 7261 21069
rect 7317 21013 7403 21069
rect 7459 21013 7545 21069
rect 7601 21013 7687 21069
rect 7743 21013 7829 21069
rect 7885 21013 7971 21069
rect 8027 21013 8113 21069
rect 8169 21013 8255 21069
rect 8311 21013 8397 21069
rect 8453 21013 8539 21069
rect 8595 21013 8681 21069
rect 8737 21013 8823 21069
rect 8879 21013 8965 21069
rect 9021 21013 9107 21069
rect 9163 21013 9249 21069
rect 9305 21013 9391 21069
rect 9447 21013 9533 21069
rect 9589 21013 9675 21069
rect 9731 21013 9817 21069
rect 9873 21013 9959 21069
rect 10015 21013 10101 21069
rect 10157 21013 10243 21069
rect 10299 21013 10385 21069
rect 10441 21013 10527 21069
rect 10583 21013 10669 21069
rect 10725 21013 10811 21069
rect 10867 21013 10953 21069
rect 11009 21013 11095 21069
rect 11151 21013 11237 21069
rect 11293 21013 11379 21069
rect 11435 21013 11521 21069
rect 11577 21013 11663 21069
rect 11719 21013 11805 21069
rect 11861 21013 11947 21069
rect 12003 21013 12089 21069
rect 12145 21013 12231 21069
rect 12287 21013 12373 21069
rect 12429 21013 12515 21069
rect 12571 21013 12657 21069
rect 12713 21013 12799 21069
rect 12855 21013 12941 21069
rect 12997 21013 13083 21069
rect 13139 21013 13225 21069
rect 13281 21013 13367 21069
rect 13423 21013 13509 21069
rect 13565 21013 13651 21069
rect 13707 21013 13793 21069
rect 13849 21013 13935 21069
rect 13991 21013 14077 21069
rect 14133 21013 14219 21069
rect 14275 21013 14361 21069
rect 14417 21013 14503 21069
rect 14559 21013 14645 21069
rect 14701 21013 14787 21069
rect 14843 21013 15000 21069
rect 0 20927 15000 21013
rect 0 20871 161 20927
rect 217 20871 303 20927
rect 359 20871 445 20927
rect 501 20871 587 20927
rect 643 20871 729 20927
rect 785 20871 871 20927
rect 927 20871 1013 20927
rect 1069 20871 1155 20927
rect 1211 20871 1297 20927
rect 1353 20871 1439 20927
rect 1495 20871 1581 20927
rect 1637 20871 1723 20927
rect 1779 20871 1865 20927
rect 1921 20871 2007 20927
rect 2063 20871 2149 20927
rect 2205 20871 2291 20927
rect 2347 20871 2433 20927
rect 2489 20871 2575 20927
rect 2631 20871 2717 20927
rect 2773 20871 2859 20927
rect 2915 20871 3001 20927
rect 3057 20871 3143 20927
rect 3199 20871 3285 20927
rect 3341 20871 3427 20927
rect 3483 20871 3569 20927
rect 3625 20871 3711 20927
rect 3767 20871 3853 20927
rect 3909 20871 3995 20927
rect 4051 20871 4137 20927
rect 4193 20871 4279 20927
rect 4335 20871 4421 20927
rect 4477 20871 4563 20927
rect 4619 20871 4705 20927
rect 4761 20871 4847 20927
rect 4903 20871 4989 20927
rect 5045 20871 5131 20927
rect 5187 20871 5273 20927
rect 5329 20871 5415 20927
rect 5471 20871 5557 20927
rect 5613 20871 5699 20927
rect 5755 20871 5841 20927
rect 5897 20871 5983 20927
rect 6039 20871 6125 20927
rect 6181 20871 6267 20927
rect 6323 20871 6409 20927
rect 6465 20871 6551 20927
rect 6607 20871 6693 20927
rect 6749 20871 6835 20927
rect 6891 20871 6977 20927
rect 7033 20871 7119 20927
rect 7175 20871 7261 20927
rect 7317 20871 7403 20927
rect 7459 20871 7545 20927
rect 7601 20871 7687 20927
rect 7743 20871 7829 20927
rect 7885 20871 7971 20927
rect 8027 20871 8113 20927
rect 8169 20871 8255 20927
rect 8311 20871 8397 20927
rect 8453 20871 8539 20927
rect 8595 20871 8681 20927
rect 8737 20871 8823 20927
rect 8879 20871 8965 20927
rect 9021 20871 9107 20927
rect 9163 20871 9249 20927
rect 9305 20871 9391 20927
rect 9447 20871 9533 20927
rect 9589 20871 9675 20927
rect 9731 20871 9817 20927
rect 9873 20871 9959 20927
rect 10015 20871 10101 20927
rect 10157 20871 10243 20927
rect 10299 20871 10385 20927
rect 10441 20871 10527 20927
rect 10583 20871 10669 20927
rect 10725 20871 10811 20927
rect 10867 20871 10953 20927
rect 11009 20871 11095 20927
rect 11151 20871 11237 20927
rect 11293 20871 11379 20927
rect 11435 20871 11521 20927
rect 11577 20871 11663 20927
rect 11719 20871 11805 20927
rect 11861 20871 11947 20927
rect 12003 20871 12089 20927
rect 12145 20871 12231 20927
rect 12287 20871 12373 20927
rect 12429 20871 12515 20927
rect 12571 20871 12657 20927
rect 12713 20871 12799 20927
rect 12855 20871 12941 20927
rect 12997 20871 13083 20927
rect 13139 20871 13225 20927
rect 13281 20871 13367 20927
rect 13423 20871 13509 20927
rect 13565 20871 13651 20927
rect 13707 20871 13793 20927
rect 13849 20871 13935 20927
rect 13991 20871 14077 20927
rect 14133 20871 14219 20927
rect 14275 20871 14361 20927
rect 14417 20871 14503 20927
rect 14559 20871 14645 20927
rect 14701 20871 14787 20927
rect 14843 20871 15000 20927
rect 0 20785 15000 20871
rect 0 20729 161 20785
rect 217 20729 303 20785
rect 359 20729 445 20785
rect 501 20729 587 20785
rect 643 20729 729 20785
rect 785 20729 871 20785
rect 927 20729 1013 20785
rect 1069 20729 1155 20785
rect 1211 20729 1297 20785
rect 1353 20729 1439 20785
rect 1495 20729 1581 20785
rect 1637 20729 1723 20785
rect 1779 20729 1865 20785
rect 1921 20729 2007 20785
rect 2063 20729 2149 20785
rect 2205 20729 2291 20785
rect 2347 20729 2433 20785
rect 2489 20729 2575 20785
rect 2631 20729 2717 20785
rect 2773 20729 2859 20785
rect 2915 20729 3001 20785
rect 3057 20729 3143 20785
rect 3199 20729 3285 20785
rect 3341 20729 3427 20785
rect 3483 20729 3569 20785
rect 3625 20729 3711 20785
rect 3767 20729 3853 20785
rect 3909 20729 3995 20785
rect 4051 20729 4137 20785
rect 4193 20729 4279 20785
rect 4335 20729 4421 20785
rect 4477 20729 4563 20785
rect 4619 20729 4705 20785
rect 4761 20729 4847 20785
rect 4903 20729 4989 20785
rect 5045 20729 5131 20785
rect 5187 20729 5273 20785
rect 5329 20729 5415 20785
rect 5471 20729 5557 20785
rect 5613 20729 5699 20785
rect 5755 20729 5841 20785
rect 5897 20729 5983 20785
rect 6039 20729 6125 20785
rect 6181 20729 6267 20785
rect 6323 20729 6409 20785
rect 6465 20729 6551 20785
rect 6607 20729 6693 20785
rect 6749 20729 6835 20785
rect 6891 20729 6977 20785
rect 7033 20729 7119 20785
rect 7175 20729 7261 20785
rect 7317 20729 7403 20785
rect 7459 20729 7545 20785
rect 7601 20729 7687 20785
rect 7743 20729 7829 20785
rect 7885 20729 7971 20785
rect 8027 20729 8113 20785
rect 8169 20729 8255 20785
rect 8311 20729 8397 20785
rect 8453 20729 8539 20785
rect 8595 20729 8681 20785
rect 8737 20729 8823 20785
rect 8879 20729 8965 20785
rect 9021 20729 9107 20785
rect 9163 20729 9249 20785
rect 9305 20729 9391 20785
rect 9447 20729 9533 20785
rect 9589 20729 9675 20785
rect 9731 20729 9817 20785
rect 9873 20729 9959 20785
rect 10015 20729 10101 20785
rect 10157 20729 10243 20785
rect 10299 20729 10385 20785
rect 10441 20729 10527 20785
rect 10583 20729 10669 20785
rect 10725 20729 10811 20785
rect 10867 20729 10953 20785
rect 11009 20729 11095 20785
rect 11151 20729 11237 20785
rect 11293 20729 11379 20785
rect 11435 20729 11521 20785
rect 11577 20729 11663 20785
rect 11719 20729 11805 20785
rect 11861 20729 11947 20785
rect 12003 20729 12089 20785
rect 12145 20729 12231 20785
rect 12287 20729 12373 20785
rect 12429 20729 12515 20785
rect 12571 20729 12657 20785
rect 12713 20729 12799 20785
rect 12855 20729 12941 20785
rect 12997 20729 13083 20785
rect 13139 20729 13225 20785
rect 13281 20729 13367 20785
rect 13423 20729 13509 20785
rect 13565 20729 13651 20785
rect 13707 20729 13793 20785
rect 13849 20729 13935 20785
rect 13991 20729 14077 20785
rect 14133 20729 14219 20785
rect 14275 20729 14361 20785
rect 14417 20729 14503 20785
rect 14559 20729 14645 20785
rect 14701 20729 14787 20785
rect 14843 20729 15000 20785
rect 0 20643 15000 20729
rect 0 20587 161 20643
rect 217 20587 303 20643
rect 359 20587 445 20643
rect 501 20587 587 20643
rect 643 20587 729 20643
rect 785 20587 871 20643
rect 927 20587 1013 20643
rect 1069 20587 1155 20643
rect 1211 20587 1297 20643
rect 1353 20587 1439 20643
rect 1495 20587 1581 20643
rect 1637 20587 1723 20643
rect 1779 20587 1865 20643
rect 1921 20587 2007 20643
rect 2063 20587 2149 20643
rect 2205 20587 2291 20643
rect 2347 20587 2433 20643
rect 2489 20587 2575 20643
rect 2631 20587 2717 20643
rect 2773 20587 2859 20643
rect 2915 20587 3001 20643
rect 3057 20587 3143 20643
rect 3199 20587 3285 20643
rect 3341 20587 3427 20643
rect 3483 20587 3569 20643
rect 3625 20587 3711 20643
rect 3767 20587 3853 20643
rect 3909 20587 3995 20643
rect 4051 20587 4137 20643
rect 4193 20587 4279 20643
rect 4335 20587 4421 20643
rect 4477 20587 4563 20643
rect 4619 20587 4705 20643
rect 4761 20587 4847 20643
rect 4903 20587 4989 20643
rect 5045 20587 5131 20643
rect 5187 20587 5273 20643
rect 5329 20587 5415 20643
rect 5471 20587 5557 20643
rect 5613 20587 5699 20643
rect 5755 20587 5841 20643
rect 5897 20587 5983 20643
rect 6039 20587 6125 20643
rect 6181 20587 6267 20643
rect 6323 20587 6409 20643
rect 6465 20587 6551 20643
rect 6607 20587 6693 20643
rect 6749 20587 6835 20643
rect 6891 20587 6977 20643
rect 7033 20587 7119 20643
rect 7175 20587 7261 20643
rect 7317 20587 7403 20643
rect 7459 20587 7545 20643
rect 7601 20587 7687 20643
rect 7743 20587 7829 20643
rect 7885 20587 7971 20643
rect 8027 20587 8113 20643
rect 8169 20587 8255 20643
rect 8311 20587 8397 20643
rect 8453 20587 8539 20643
rect 8595 20587 8681 20643
rect 8737 20587 8823 20643
rect 8879 20587 8965 20643
rect 9021 20587 9107 20643
rect 9163 20587 9249 20643
rect 9305 20587 9391 20643
rect 9447 20587 9533 20643
rect 9589 20587 9675 20643
rect 9731 20587 9817 20643
rect 9873 20587 9959 20643
rect 10015 20587 10101 20643
rect 10157 20587 10243 20643
rect 10299 20587 10385 20643
rect 10441 20587 10527 20643
rect 10583 20587 10669 20643
rect 10725 20587 10811 20643
rect 10867 20587 10953 20643
rect 11009 20587 11095 20643
rect 11151 20587 11237 20643
rect 11293 20587 11379 20643
rect 11435 20587 11521 20643
rect 11577 20587 11663 20643
rect 11719 20587 11805 20643
rect 11861 20587 11947 20643
rect 12003 20587 12089 20643
rect 12145 20587 12231 20643
rect 12287 20587 12373 20643
rect 12429 20587 12515 20643
rect 12571 20587 12657 20643
rect 12713 20587 12799 20643
rect 12855 20587 12941 20643
rect 12997 20587 13083 20643
rect 13139 20587 13225 20643
rect 13281 20587 13367 20643
rect 13423 20587 13509 20643
rect 13565 20587 13651 20643
rect 13707 20587 13793 20643
rect 13849 20587 13935 20643
rect 13991 20587 14077 20643
rect 14133 20587 14219 20643
rect 14275 20587 14361 20643
rect 14417 20587 14503 20643
rect 14559 20587 14645 20643
rect 14701 20587 14787 20643
rect 14843 20587 15000 20643
rect 0 20501 15000 20587
rect 0 20445 161 20501
rect 217 20445 303 20501
rect 359 20445 445 20501
rect 501 20445 587 20501
rect 643 20445 729 20501
rect 785 20445 871 20501
rect 927 20445 1013 20501
rect 1069 20445 1155 20501
rect 1211 20445 1297 20501
rect 1353 20445 1439 20501
rect 1495 20445 1581 20501
rect 1637 20445 1723 20501
rect 1779 20445 1865 20501
rect 1921 20445 2007 20501
rect 2063 20445 2149 20501
rect 2205 20445 2291 20501
rect 2347 20445 2433 20501
rect 2489 20445 2575 20501
rect 2631 20445 2717 20501
rect 2773 20445 2859 20501
rect 2915 20445 3001 20501
rect 3057 20445 3143 20501
rect 3199 20445 3285 20501
rect 3341 20445 3427 20501
rect 3483 20445 3569 20501
rect 3625 20445 3711 20501
rect 3767 20445 3853 20501
rect 3909 20445 3995 20501
rect 4051 20445 4137 20501
rect 4193 20445 4279 20501
rect 4335 20445 4421 20501
rect 4477 20445 4563 20501
rect 4619 20445 4705 20501
rect 4761 20445 4847 20501
rect 4903 20445 4989 20501
rect 5045 20445 5131 20501
rect 5187 20445 5273 20501
rect 5329 20445 5415 20501
rect 5471 20445 5557 20501
rect 5613 20445 5699 20501
rect 5755 20445 5841 20501
rect 5897 20445 5983 20501
rect 6039 20445 6125 20501
rect 6181 20445 6267 20501
rect 6323 20445 6409 20501
rect 6465 20445 6551 20501
rect 6607 20445 6693 20501
rect 6749 20445 6835 20501
rect 6891 20445 6977 20501
rect 7033 20445 7119 20501
rect 7175 20445 7261 20501
rect 7317 20445 7403 20501
rect 7459 20445 7545 20501
rect 7601 20445 7687 20501
rect 7743 20445 7829 20501
rect 7885 20445 7971 20501
rect 8027 20445 8113 20501
rect 8169 20445 8255 20501
rect 8311 20445 8397 20501
rect 8453 20445 8539 20501
rect 8595 20445 8681 20501
rect 8737 20445 8823 20501
rect 8879 20445 8965 20501
rect 9021 20445 9107 20501
rect 9163 20445 9249 20501
rect 9305 20445 9391 20501
rect 9447 20445 9533 20501
rect 9589 20445 9675 20501
rect 9731 20445 9817 20501
rect 9873 20445 9959 20501
rect 10015 20445 10101 20501
rect 10157 20445 10243 20501
rect 10299 20445 10385 20501
rect 10441 20445 10527 20501
rect 10583 20445 10669 20501
rect 10725 20445 10811 20501
rect 10867 20445 10953 20501
rect 11009 20445 11095 20501
rect 11151 20445 11237 20501
rect 11293 20445 11379 20501
rect 11435 20445 11521 20501
rect 11577 20445 11663 20501
rect 11719 20445 11805 20501
rect 11861 20445 11947 20501
rect 12003 20445 12089 20501
rect 12145 20445 12231 20501
rect 12287 20445 12373 20501
rect 12429 20445 12515 20501
rect 12571 20445 12657 20501
rect 12713 20445 12799 20501
rect 12855 20445 12941 20501
rect 12997 20445 13083 20501
rect 13139 20445 13225 20501
rect 13281 20445 13367 20501
rect 13423 20445 13509 20501
rect 13565 20445 13651 20501
rect 13707 20445 13793 20501
rect 13849 20445 13935 20501
rect 13991 20445 14077 20501
rect 14133 20445 14219 20501
rect 14275 20445 14361 20501
rect 14417 20445 14503 20501
rect 14559 20445 14645 20501
rect 14701 20445 14787 20501
rect 14843 20445 15000 20501
rect 0 20400 15000 20445
rect 937 20200 3937 20400
rect 4337 20200 7337 20400
rect 7737 20200 10737 20400
rect 11137 20200 14137 20400
rect 0 20141 15000 20200
rect 0 20085 161 20141
rect 217 20085 303 20141
rect 359 20085 445 20141
rect 501 20085 587 20141
rect 643 20085 729 20141
rect 785 20085 871 20141
rect 927 20085 1013 20141
rect 1069 20085 1155 20141
rect 1211 20085 1297 20141
rect 1353 20085 1439 20141
rect 1495 20085 1581 20141
rect 1637 20085 1723 20141
rect 1779 20085 1865 20141
rect 1921 20085 2007 20141
rect 2063 20085 2149 20141
rect 2205 20085 2291 20141
rect 2347 20085 2433 20141
rect 2489 20085 2575 20141
rect 2631 20085 2717 20141
rect 2773 20085 2859 20141
rect 2915 20085 3001 20141
rect 3057 20085 3143 20141
rect 3199 20085 3285 20141
rect 3341 20085 3427 20141
rect 3483 20085 3569 20141
rect 3625 20085 3711 20141
rect 3767 20085 3853 20141
rect 3909 20085 3995 20141
rect 4051 20085 4137 20141
rect 4193 20085 4279 20141
rect 4335 20085 4421 20141
rect 4477 20085 4563 20141
rect 4619 20085 4705 20141
rect 4761 20085 4847 20141
rect 4903 20085 4989 20141
rect 5045 20085 5131 20141
rect 5187 20085 5273 20141
rect 5329 20085 5415 20141
rect 5471 20085 5557 20141
rect 5613 20085 5699 20141
rect 5755 20085 5841 20141
rect 5897 20085 5983 20141
rect 6039 20085 6125 20141
rect 6181 20085 6267 20141
rect 6323 20085 6409 20141
rect 6465 20085 6551 20141
rect 6607 20085 6693 20141
rect 6749 20085 6835 20141
rect 6891 20085 6977 20141
rect 7033 20085 7119 20141
rect 7175 20085 7261 20141
rect 7317 20085 7403 20141
rect 7459 20085 7545 20141
rect 7601 20085 7687 20141
rect 7743 20085 7829 20141
rect 7885 20085 7971 20141
rect 8027 20085 8113 20141
rect 8169 20085 8255 20141
rect 8311 20085 8397 20141
rect 8453 20085 8539 20141
rect 8595 20085 8681 20141
rect 8737 20085 8823 20141
rect 8879 20085 8965 20141
rect 9021 20085 9107 20141
rect 9163 20085 9249 20141
rect 9305 20085 9391 20141
rect 9447 20085 9533 20141
rect 9589 20085 9675 20141
rect 9731 20085 9817 20141
rect 9873 20085 9959 20141
rect 10015 20085 10101 20141
rect 10157 20085 10243 20141
rect 10299 20085 10385 20141
rect 10441 20085 10527 20141
rect 10583 20085 10669 20141
rect 10725 20085 10811 20141
rect 10867 20085 10953 20141
rect 11009 20085 11095 20141
rect 11151 20085 11237 20141
rect 11293 20085 11379 20141
rect 11435 20085 11521 20141
rect 11577 20085 11663 20141
rect 11719 20085 11805 20141
rect 11861 20085 11947 20141
rect 12003 20085 12089 20141
rect 12145 20085 12231 20141
rect 12287 20085 12373 20141
rect 12429 20085 12515 20141
rect 12571 20085 12657 20141
rect 12713 20085 12799 20141
rect 12855 20085 12941 20141
rect 12997 20085 13083 20141
rect 13139 20085 13225 20141
rect 13281 20085 13367 20141
rect 13423 20085 13509 20141
rect 13565 20085 13651 20141
rect 13707 20085 13793 20141
rect 13849 20085 13935 20141
rect 13991 20085 14077 20141
rect 14133 20085 14219 20141
rect 14275 20085 14361 20141
rect 14417 20085 14503 20141
rect 14559 20085 14645 20141
rect 14701 20085 14787 20141
rect 14843 20085 15000 20141
rect 0 19999 15000 20085
rect 0 19943 161 19999
rect 217 19943 303 19999
rect 359 19943 445 19999
rect 501 19943 587 19999
rect 643 19943 729 19999
rect 785 19943 871 19999
rect 927 19943 1013 19999
rect 1069 19943 1155 19999
rect 1211 19943 1297 19999
rect 1353 19943 1439 19999
rect 1495 19943 1581 19999
rect 1637 19943 1723 19999
rect 1779 19943 1865 19999
rect 1921 19943 2007 19999
rect 2063 19943 2149 19999
rect 2205 19943 2291 19999
rect 2347 19943 2433 19999
rect 2489 19943 2575 19999
rect 2631 19943 2717 19999
rect 2773 19943 2859 19999
rect 2915 19943 3001 19999
rect 3057 19943 3143 19999
rect 3199 19943 3285 19999
rect 3341 19943 3427 19999
rect 3483 19943 3569 19999
rect 3625 19943 3711 19999
rect 3767 19943 3853 19999
rect 3909 19943 3995 19999
rect 4051 19943 4137 19999
rect 4193 19943 4279 19999
rect 4335 19943 4421 19999
rect 4477 19943 4563 19999
rect 4619 19943 4705 19999
rect 4761 19943 4847 19999
rect 4903 19943 4989 19999
rect 5045 19943 5131 19999
rect 5187 19943 5273 19999
rect 5329 19943 5415 19999
rect 5471 19943 5557 19999
rect 5613 19943 5699 19999
rect 5755 19943 5841 19999
rect 5897 19943 5983 19999
rect 6039 19943 6125 19999
rect 6181 19943 6267 19999
rect 6323 19943 6409 19999
rect 6465 19943 6551 19999
rect 6607 19943 6693 19999
rect 6749 19943 6835 19999
rect 6891 19943 6977 19999
rect 7033 19943 7119 19999
rect 7175 19943 7261 19999
rect 7317 19943 7403 19999
rect 7459 19943 7545 19999
rect 7601 19943 7687 19999
rect 7743 19943 7829 19999
rect 7885 19943 7971 19999
rect 8027 19943 8113 19999
rect 8169 19943 8255 19999
rect 8311 19943 8397 19999
rect 8453 19943 8539 19999
rect 8595 19943 8681 19999
rect 8737 19943 8823 19999
rect 8879 19943 8965 19999
rect 9021 19943 9107 19999
rect 9163 19943 9249 19999
rect 9305 19943 9391 19999
rect 9447 19943 9533 19999
rect 9589 19943 9675 19999
rect 9731 19943 9817 19999
rect 9873 19943 9959 19999
rect 10015 19943 10101 19999
rect 10157 19943 10243 19999
rect 10299 19943 10385 19999
rect 10441 19943 10527 19999
rect 10583 19943 10669 19999
rect 10725 19943 10811 19999
rect 10867 19943 10953 19999
rect 11009 19943 11095 19999
rect 11151 19943 11237 19999
rect 11293 19943 11379 19999
rect 11435 19943 11521 19999
rect 11577 19943 11663 19999
rect 11719 19943 11805 19999
rect 11861 19943 11947 19999
rect 12003 19943 12089 19999
rect 12145 19943 12231 19999
rect 12287 19943 12373 19999
rect 12429 19943 12515 19999
rect 12571 19943 12657 19999
rect 12713 19943 12799 19999
rect 12855 19943 12941 19999
rect 12997 19943 13083 19999
rect 13139 19943 13225 19999
rect 13281 19943 13367 19999
rect 13423 19943 13509 19999
rect 13565 19943 13651 19999
rect 13707 19943 13793 19999
rect 13849 19943 13935 19999
rect 13991 19943 14077 19999
rect 14133 19943 14219 19999
rect 14275 19943 14361 19999
rect 14417 19943 14503 19999
rect 14559 19943 14645 19999
rect 14701 19943 14787 19999
rect 14843 19943 15000 19999
rect 0 19857 15000 19943
rect 0 19801 161 19857
rect 217 19801 303 19857
rect 359 19801 445 19857
rect 501 19801 587 19857
rect 643 19801 729 19857
rect 785 19801 871 19857
rect 927 19801 1013 19857
rect 1069 19801 1155 19857
rect 1211 19801 1297 19857
rect 1353 19801 1439 19857
rect 1495 19801 1581 19857
rect 1637 19801 1723 19857
rect 1779 19801 1865 19857
rect 1921 19801 2007 19857
rect 2063 19801 2149 19857
rect 2205 19801 2291 19857
rect 2347 19801 2433 19857
rect 2489 19801 2575 19857
rect 2631 19801 2717 19857
rect 2773 19801 2859 19857
rect 2915 19801 3001 19857
rect 3057 19801 3143 19857
rect 3199 19801 3285 19857
rect 3341 19801 3427 19857
rect 3483 19801 3569 19857
rect 3625 19801 3711 19857
rect 3767 19801 3853 19857
rect 3909 19801 3995 19857
rect 4051 19801 4137 19857
rect 4193 19801 4279 19857
rect 4335 19801 4421 19857
rect 4477 19801 4563 19857
rect 4619 19801 4705 19857
rect 4761 19801 4847 19857
rect 4903 19801 4989 19857
rect 5045 19801 5131 19857
rect 5187 19801 5273 19857
rect 5329 19801 5415 19857
rect 5471 19801 5557 19857
rect 5613 19801 5699 19857
rect 5755 19801 5841 19857
rect 5897 19801 5983 19857
rect 6039 19801 6125 19857
rect 6181 19801 6267 19857
rect 6323 19801 6409 19857
rect 6465 19801 6551 19857
rect 6607 19801 6693 19857
rect 6749 19801 6835 19857
rect 6891 19801 6977 19857
rect 7033 19801 7119 19857
rect 7175 19801 7261 19857
rect 7317 19801 7403 19857
rect 7459 19801 7545 19857
rect 7601 19801 7687 19857
rect 7743 19801 7829 19857
rect 7885 19801 7971 19857
rect 8027 19801 8113 19857
rect 8169 19801 8255 19857
rect 8311 19801 8397 19857
rect 8453 19801 8539 19857
rect 8595 19801 8681 19857
rect 8737 19801 8823 19857
rect 8879 19801 8965 19857
rect 9021 19801 9107 19857
rect 9163 19801 9249 19857
rect 9305 19801 9391 19857
rect 9447 19801 9533 19857
rect 9589 19801 9675 19857
rect 9731 19801 9817 19857
rect 9873 19801 9959 19857
rect 10015 19801 10101 19857
rect 10157 19801 10243 19857
rect 10299 19801 10385 19857
rect 10441 19801 10527 19857
rect 10583 19801 10669 19857
rect 10725 19801 10811 19857
rect 10867 19801 10953 19857
rect 11009 19801 11095 19857
rect 11151 19801 11237 19857
rect 11293 19801 11379 19857
rect 11435 19801 11521 19857
rect 11577 19801 11663 19857
rect 11719 19801 11805 19857
rect 11861 19801 11947 19857
rect 12003 19801 12089 19857
rect 12145 19801 12231 19857
rect 12287 19801 12373 19857
rect 12429 19801 12515 19857
rect 12571 19801 12657 19857
rect 12713 19801 12799 19857
rect 12855 19801 12941 19857
rect 12997 19801 13083 19857
rect 13139 19801 13225 19857
rect 13281 19801 13367 19857
rect 13423 19801 13509 19857
rect 13565 19801 13651 19857
rect 13707 19801 13793 19857
rect 13849 19801 13935 19857
rect 13991 19801 14077 19857
rect 14133 19801 14219 19857
rect 14275 19801 14361 19857
rect 14417 19801 14503 19857
rect 14559 19801 14645 19857
rect 14701 19801 14787 19857
rect 14843 19801 15000 19857
rect 0 19715 15000 19801
rect 0 19659 161 19715
rect 217 19659 303 19715
rect 359 19659 445 19715
rect 501 19659 587 19715
rect 643 19659 729 19715
rect 785 19659 871 19715
rect 927 19659 1013 19715
rect 1069 19659 1155 19715
rect 1211 19659 1297 19715
rect 1353 19659 1439 19715
rect 1495 19659 1581 19715
rect 1637 19659 1723 19715
rect 1779 19659 1865 19715
rect 1921 19659 2007 19715
rect 2063 19659 2149 19715
rect 2205 19659 2291 19715
rect 2347 19659 2433 19715
rect 2489 19659 2575 19715
rect 2631 19659 2717 19715
rect 2773 19659 2859 19715
rect 2915 19659 3001 19715
rect 3057 19659 3143 19715
rect 3199 19659 3285 19715
rect 3341 19659 3427 19715
rect 3483 19659 3569 19715
rect 3625 19659 3711 19715
rect 3767 19659 3853 19715
rect 3909 19659 3995 19715
rect 4051 19659 4137 19715
rect 4193 19659 4279 19715
rect 4335 19659 4421 19715
rect 4477 19659 4563 19715
rect 4619 19659 4705 19715
rect 4761 19659 4847 19715
rect 4903 19659 4989 19715
rect 5045 19659 5131 19715
rect 5187 19659 5273 19715
rect 5329 19659 5415 19715
rect 5471 19659 5557 19715
rect 5613 19659 5699 19715
rect 5755 19659 5841 19715
rect 5897 19659 5983 19715
rect 6039 19659 6125 19715
rect 6181 19659 6267 19715
rect 6323 19659 6409 19715
rect 6465 19659 6551 19715
rect 6607 19659 6693 19715
rect 6749 19659 6835 19715
rect 6891 19659 6977 19715
rect 7033 19659 7119 19715
rect 7175 19659 7261 19715
rect 7317 19659 7403 19715
rect 7459 19659 7545 19715
rect 7601 19659 7687 19715
rect 7743 19659 7829 19715
rect 7885 19659 7971 19715
rect 8027 19659 8113 19715
rect 8169 19659 8255 19715
rect 8311 19659 8397 19715
rect 8453 19659 8539 19715
rect 8595 19659 8681 19715
rect 8737 19659 8823 19715
rect 8879 19659 8965 19715
rect 9021 19659 9107 19715
rect 9163 19659 9249 19715
rect 9305 19659 9391 19715
rect 9447 19659 9533 19715
rect 9589 19659 9675 19715
rect 9731 19659 9817 19715
rect 9873 19659 9959 19715
rect 10015 19659 10101 19715
rect 10157 19659 10243 19715
rect 10299 19659 10385 19715
rect 10441 19659 10527 19715
rect 10583 19659 10669 19715
rect 10725 19659 10811 19715
rect 10867 19659 10953 19715
rect 11009 19659 11095 19715
rect 11151 19659 11237 19715
rect 11293 19659 11379 19715
rect 11435 19659 11521 19715
rect 11577 19659 11663 19715
rect 11719 19659 11805 19715
rect 11861 19659 11947 19715
rect 12003 19659 12089 19715
rect 12145 19659 12231 19715
rect 12287 19659 12373 19715
rect 12429 19659 12515 19715
rect 12571 19659 12657 19715
rect 12713 19659 12799 19715
rect 12855 19659 12941 19715
rect 12997 19659 13083 19715
rect 13139 19659 13225 19715
rect 13281 19659 13367 19715
rect 13423 19659 13509 19715
rect 13565 19659 13651 19715
rect 13707 19659 13793 19715
rect 13849 19659 13935 19715
rect 13991 19659 14077 19715
rect 14133 19659 14219 19715
rect 14275 19659 14361 19715
rect 14417 19659 14503 19715
rect 14559 19659 14645 19715
rect 14701 19659 14787 19715
rect 14843 19659 15000 19715
rect 0 19573 15000 19659
rect 0 19517 161 19573
rect 217 19517 303 19573
rect 359 19517 445 19573
rect 501 19517 587 19573
rect 643 19517 729 19573
rect 785 19517 871 19573
rect 927 19517 1013 19573
rect 1069 19517 1155 19573
rect 1211 19517 1297 19573
rect 1353 19517 1439 19573
rect 1495 19517 1581 19573
rect 1637 19517 1723 19573
rect 1779 19517 1865 19573
rect 1921 19517 2007 19573
rect 2063 19517 2149 19573
rect 2205 19517 2291 19573
rect 2347 19517 2433 19573
rect 2489 19517 2575 19573
rect 2631 19517 2717 19573
rect 2773 19517 2859 19573
rect 2915 19517 3001 19573
rect 3057 19517 3143 19573
rect 3199 19517 3285 19573
rect 3341 19517 3427 19573
rect 3483 19517 3569 19573
rect 3625 19517 3711 19573
rect 3767 19517 3853 19573
rect 3909 19517 3995 19573
rect 4051 19517 4137 19573
rect 4193 19517 4279 19573
rect 4335 19517 4421 19573
rect 4477 19517 4563 19573
rect 4619 19517 4705 19573
rect 4761 19517 4847 19573
rect 4903 19517 4989 19573
rect 5045 19517 5131 19573
rect 5187 19517 5273 19573
rect 5329 19517 5415 19573
rect 5471 19517 5557 19573
rect 5613 19517 5699 19573
rect 5755 19517 5841 19573
rect 5897 19517 5983 19573
rect 6039 19517 6125 19573
rect 6181 19517 6267 19573
rect 6323 19517 6409 19573
rect 6465 19517 6551 19573
rect 6607 19517 6693 19573
rect 6749 19517 6835 19573
rect 6891 19517 6977 19573
rect 7033 19517 7119 19573
rect 7175 19517 7261 19573
rect 7317 19517 7403 19573
rect 7459 19517 7545 19573
rect 7601 19517 7687 19573
rect 7743 19517 7829 19573
rect 7885 19517 7971 19573
rect 8027 19517 8113 19573
rect 8169 19517 8255 19573
rect 8311 19517 8397 19573
rect 8453 19517 8539 19573
rect 8595 19517 8681 19573
rect 8737 19517 8823 19573
rect 8879 19517 8965 19573
rect 9021 19517 9107 19573
rect 9163 19517 9249 19573
rect 9305 19517 9391 19573
rect 9447 19517 9533 19573
rect 9589 19517 9675 19573
rect 9731 19517 9817 19573
rect 9873 19517 9959 19573
rect 10015 19517 10101 19573
rect 10157 19517 10243 19573
rect 10299 19517 10385 19573
rect 10441 19517 10527 19573
rect 10583 19517 10669 19573
rect 10725 19517 10811 19573
rect 10867 19517 10953 19573
rect 11009 19517 11095 19573
rect 11151 19517 11237 19573
rect 11293 19517 11379 19573
rect 11435 19517 11521 19573
rect 11577 19517 11663 19573
rect 11719 19517 11805 19573
rect 11861 19517 11947 19573
rect 12003 19517 12089 19573
rect 12145 19517 12231 19573
rect 12287 19517 12373 19573
rect 12429 19517 12515 19573
rect 12571 19517 12657 19573
rect 12713 19517 12799 19573
rect 12855 19517 12941 19573
rect 12997 19517 13083 19573
rect 13139 19517 13225 19573
rect 13281 19517 13367 19573
rect 13423 19517 13509 19573
rect 13565 19517 13651 19573
rect 13707 19517 13793 19573
rect 13849 19517 13935 19573
rect 13991 19517 14077 19573
rect 14133 19517 14219 19573
rect 14275 19517 14361 19573
rect 14417 19517 14503 19573
rect 14559 19517 14645 19573
rect 14701 19517 14787 19573
rect 14843 19517 15000 19573
rect 0 19431 15000 19517
rect 0 19375 161 19431
rect 217 19375 303 19431
rect 359 19375 445 19431
rect 501 19375 587 19431
rect 643 19375 729 19431
rect 785 19375 871 19431
rect 927 19375 1013 19431
rect 1069 19375 1155 19431
rect 1211 19375 1297 19431
rect 1353 19375 1439 19431
rect 1495 19375 1581 19431
rect 1637 19375 1723 19431
rect 1779 19375 1865 19431
rect 1921 19375 2007 19431
rect 2063 19375 2149 19431
rect 2205 19375 2291 19431
rect 2347 19375 2433 19431
rect 2489 19375 2575 19431
rect 2631 19375 2717 19431
rect 2773 19375 2859 19431
rect 2915 19375 3001 19431
rect 3057 19375 3143 19431
rect 3199 19375 3285 19431
rect 3341 19375 3427 19431
rect 3483 19375 3569 19431
rect 3625 19375 3711 19431
rect 3767 19375 3853 19431
rect 3909 19375 3995 19431
rect 4051 19375 4137 19431
rect 4193 19375 4279 19431
rect 4335 19375 4421 19431
rect 4477 19375 4563 19431
rect 4619 19375 4705 19431
rect 4761 19375 4847 19431
rect 4903 19375 4989 19431
rect 5045 19375 5131 19431
rect 5187 19375 5273 19431
rect 5329 19375 5415 19431
rect 5471 19375 5557 19431
rect 5613 19375 5699 19431
rect 5755 19375 5841 19431
rect 5897 19375 5983 19431
rect 6039 19375 6125 19431
rect 6181 19375 6267 19431
rect 6323 19375 6409 19431
rect 6465 19375 6551 19431
rect 6607 19375 6693 19431
rect 6749 19375 6835 19431
rect 6891 19375 6977 19431
rect 7033 19375 7119 19431
rect 7175 19375 7261 19431
rect 7317 19375 7403 19431
rect 7459 19375 7545 19431
rect 7601 19375 7687 19431
rect 7743 19375 7829 19431
rect 7885 19375 7971 19431
rect 8027 19375 8113 19431
rect 8169 19375 8255 19431
rect 8311 19375 8397 19431
rect 8453 19375 8539 19431
rect 8595 19375 8681 19431
rect 8737 19375 8823 19431
rect 8879 19375 8965 19431
rect 9021 19375 9107 19431
rect 9163 19375 9249 19431
rect 9305 19375 9391 19431
rect 9447 19375 9533 19431
rect 9589 19375 9675 19431
rect 9731 19375 9817 19431
rect 9873 19375 9959 19431
rect 10015 19375 10101 19431
rect 10157 19375 10243 19431
rect 10299 19375 10385 19431
rect 10441 19375 10527 19431
rect 10583 19375 10669 19431
rect 10725 19375 10811 19431
rect 10867 19375 10953 19431
rect 11009 19375 11095 19431
rect 11151 19375 11237 19431
rect 11293 19375 11379 19431
rect 11435 19375 11521 19431
rect 11577 19375 11663 19431
rect 11719 19375 11805 19431
rect 11861 19375 11947 19431
rect 12003 19375 12089 19431
rect 12145 19375 12231 19431
rect 12287 19375 12373 19431
rect 12429 19375 12515 19431
rect 12571 19375 12657 19431
rect 12713 19375 12799 19431
rect 12855 19375 12941 19431
rect 12997 19375 13083 19431
rect 13139 19375 13225 19431
rect 13281 19375 13367 19431
rect 13423 19375 13509 19431
rect 13565 19375 13651 19431
rect 13707 19375 13793 19431
rect 13849 19375 13935 19431
rect 13991 19375 14077 19431
rect 14133 19375 14219 19431
rect 14275 19375 14361 19431
rect 14417 19375 14503 19431
rect 14559 19375 14645 19431
rect 14701 19375 14787 19431
rect 14843 19375 15000 19431
rect 0 19289 15000 19375
rect 0 19233 161 19289
rect 217 19233 303 19289
rect 359 19233 445 19289
rect 501 19233 587 19289
rect 643 19233 729 19289
rect 785 19233 871 19289
rect 927 19233 1013 19289
rect 1069 19233 1155 19289
rect 1211 19233 1297 19289
rect 1353 19233 1439 19289
rect 1495 19233 1581 19289
rect 1637 19233 1723 19289
rect 1779 19233 1865 19289
rect 1921 19233 2007 19289
rect 2063 19233 2149 19289
rect 2205 19233 2291 19289
rect 2347 19233 2433 19289
rect 2489 19233 2575 19289
rect 2631 19233 2717 19289
rect 2773 19233 2859 19289
rect 2915 19233 3001 19289
rect 3057 19233 3143 19289
rect 3199 19233 3285 19289
rect 3341 19233 3427 19289
rect 3483 19233 3569 19289
rect 3625 19233 3711 19289
rect 3767 19233 3853 19289
rect 3909 19233 3995 19289
rect 4051 19233 4137 19289
rect 4193 19233 4279 19289
rect 4335 19233 4421 19289
rect 4477 19233 4563 19289
rect 4619 19233 4705 19289
rect 4761 19233 4847 19289
rect 4903 19233 4989 19289
rect 5045 19233 5131 19289
rect 5187 19233 5273 19289
rect 5329 19233 5415 19289
rect 5471 19233 5557 19289
rect 5613 19233 5699 19289
rect 5755 19233 5841 19289
rect 5897 19233 5983 19289
rect 6039 19233 6125 19289
rect 6181 19233 6267 19289
rect 6323 19233 6409 19289
rect 6465 19233 6551 19289
rect 6607 19233 6693 19289
rect 6749 19233 6835 19289
rect 6891 19233 6977 19289
rect 7033 19233 7119 19289
rect 7175 19233 7261 19289
rect 7317 19233 7403 19289
rect 7459 19233 7545 19289
rect 7601 19233 7687 19289
rect 7743 19233 7829 19289
rect 7885 19233 7971 19289
rect 8027 19233 8113 19289
rect 8169 19233 8255 19289
rect 8311 19233 8397 19289
rect 8453 19233 8539 19289
rect 8595 19233 8681 19289
rect 8737 19233 8823 19289
rect 8879 19233 8965 19289
rect 9021 19233 9107 19289
rect 9163 19233 9249 19289
rect 9305 19233 9391 19289
rect 9447 19233 9533 19289
rect 9589 19233 9675 19289
rect 9731 19233 9817 19289
rect 9873 19233 9959 19289
rect 10015 19233 10101 19289
rect 10157 19233 10243 19289
rect 10299 19233 10385 19289
rect 10441 19233 10527 19289
rect 10583 19233 10669 19289
rect 10725 19233 10811 19289
rect 10867 19233 10953 19289
rect 11009 19233 11095 19289
rect 11151 19233 11237 19289
rect 11293 19233 11379 19289
rect 11435 19233 11521 19289
rect 11577 19233 11663 19289
rect 11719 19233 11805 19289
rect 11861 19233 11947 19289
rect 12003 19233 12089 19289
rect 12145 19233 12231 19289
rect 12287 19233 12373 19289
rect 12429 19233 12515 19289
rect 12571 19233 12657 19289
rect 12713 19233 12799 19289
rect 12855 19233 12941 19289
rect 12997 19233 13083 19289
rect 13139 19233 13225 19289
rect 13281 19233 13367 19289
rect 13423 19233 13509 19289
rect 13565 19233 13651 19289
rect 13707 19233 13793 19289
rect 13849 19233 13935 19289
rect 13991 19233 14077 19289
rect 14133 19233 14219 19289
rect 14275 19233 14361 19289
rect 14417 19233 14503 19289
rect 14559 19233 14645 19289
rect 14701 19233 14787 19289
rect 14843 19233 15000 19289
rect 0 19147 15000 19233
rect 0 19091 161 19147
rect 217 19091 303 19147
rect 359 19091 445 19147
rect 501 19091 587 19147
rect 643 19091 729 19147
rect 785 19091 871 19147
rect 927 19091 1013 19147
rect 1069 19091 1155 19147
rect 1211 19091 1297 19147
rect 1353 19091 1439 19147
rect 1495 19091 1581 19147
rect 1637 19091 1723 19147
rect 1779 19091 1865 19147
rect 1921 19091 2007 19147
rect 2063 19091 2149 19147
rect 2205 19091 2291 19147
rect 2347 19091 2433 19147
rect 2489 19091 2575 19147
rect 2631 19091 2717 19147
rect 2773 19091 2859 19147
rect 2915 19091 3001 19147
rect 3057 19091 3143 19147
rect 3199 19091 3285 19147
rect 3341 19091 3427 19147
rect 3483 19091 3569 19147
rect 3625 19091 3711 19147
rect 3767 19091 3853 19147
rect 3909 19091 3995 19147
rect 4051 19091 4137 19147
rect 4193 19091 4279 19147
rect 4335 19091 4421 19147
rect 4477 19091 4563 19147
rect 4619 19091 4705 19147
rect 4761 19091 4847 19147
rect 4903 19091 4989 19147
rect 5045 19091 5131 19147
rect 5187 19091 5273 19147
rect 5329 19091 5415 19147
rect 5471 19091 5557 19147
rect 5613 19091 5699 19147
rect 5755 19091 5841 19147
rect 5897 19091 5983 19147
rect 6039 19091 6125 19147
rect 6181 19091 6267 19147
rect 6323 19091 6409 19147
rect 6465 19091 6551 19147
rect 6607 19091 6693 19147
rect 6749 19091 6835 19147
rect 6891 19091 6977 19147
rect 7033 19091 7119 19147
rect 7175 19091 7261 19147
rect 7317 19091 7403 19147
rect 7459 19091 7545 19147
rect 7601 19091 7687 19147
rect 7743 19091 7829 19147
rect 7885 19091 7971 19147
rect 8027 19091 8113 19147
rect 8169 19091 8255 19147
rect 8311 19091 8397 19147
rect 8453 19091 8539 19147
rect 8595 19091 8681 19147
rect 8737 19091 8823 19147
rect 8879 19091 8965 19147
rect 9021 19091 9107 19147
rect 9163 19091 9249 19147
rect 9305 19091 9391 19147
rect 9447 19091 9533 19147
rect 9589 19091 9675 19147
rect 9731 19091 9817 19147
rect 9873 19091 9959 19147
rect 10015 19091 10101 19147
rect 10157 19091 10243 19147
rect 10299 19091 10385 19147
rect 10441 19091 10527 19147
rect 10583 19091 10669 19147
rect 10725 19091 10811 19147
rect 10867 19091 10953 19147
rect 11009 19091 11095 19147
rect 11151 19091 11237 19147
rect 11293 19091 11379 19147
rect 11435 19091 11521 19147
rect 11577 19091 11663 19147
rect 11719 19091 11805 19147
rect 11861 19091 11947 19147
rect 12003 19091 12089 19147
rect 12145 19091 12231 19147
rect 12287 19091 12373 19147
rect 12429 19091 12515 19147
rect 12571 19091 12657 19147
rect 12713 19091 12799 19147
rect 12855 19091 12941 19147
rect 12997 19091 13083 19147
rect 13139 19091 13225 19147
rect 13281 19091 13367 19147
rect 13423 19091 13509 19147
rect 13565 19091 13651 19147
rect 13707 19091 13793 19147
rect 13849 19091 13935 19147
rect 13991 19091 14077 19147
rect 14133 19091 14219 19147
rect 14275 19091 14361 19147
rect 14417 19091 14503 19147
rect 14559 19091 14645 19147
rect 14701 19091 14787 19147
rect 14843 19091 15000 19147
rect 0 19005 15000 19091
rect 0 18949 161 19005
rect 217 18949 303 19005
rect 359 18949 445 19005
rect 501 18949 587 19005
rect 643 18949 729 19005
rect 785 18949 871 19005
rect 927 18949 1013 19005
rect 1069 18949 1155 19005
rect 1211 18949 1297 19005
rect 1353 18949 1439 19005
rect 1495 18949 1581 19005
rect 1637 18949 1723 19005
rect 1779 18949 1865 19005
rect 1921 18949 2007 19005
rect 2063 18949 2149 19005
rect 2205 18949 2291 19005
rect 2347 18949 2433 19005
rect 2489 18949 2575 19005
rect 2631 18949 2717 19005
rect 2773 18949 2859 19005
rect 2915 18949 3001 19005
rect 3057 18949 3143 19005
rect 3199 18949 3285 19005
rect 3341 18949 3427 19005
rect 3483 18949 3569 19005
rect 3625 18949 3711 19005
rect 3767 18949 3853 19005
rect 3909 18949 3995 19005
rect 4051 18949 4137 19005
rect 4193 18949 4279 19005
rect 4335 18949 4421 19005
rect 4477 18949 4563 19005
rect 4619 18949 4705 19005
rect 4761 18949 4847 19005
rect 4903 18949 4989 19005
rect 5045 18949 5131 19005
rect 5187 18949 5273 19005
rect 5329 18949 5415 19005
rect 5471 18949 5557 19005
rect 5613 18949 5699 19005
rect 5755 18949 5841 19005
rect 5897 18949 5983 19005
rect 6039 18949 6125 19005
rect 6181 18949 6267 19005
rect 6323 18949 6409 19005
rect 6465 18949 6551 19005
rect 6607 18949 6693 19005
rect 6749 18949 6835 19005
rect 6891 18949 6977 19005
rect 7033 18949 7119 19005
rect 7175 18949 7261 19005
rect 7317 18949 7403 19005
rect 7459 18949 7545 19005
rect 7601 18949 7687 19005
rect 7743 18949 7829 19005
rect 7885 18949 7971 19005
rect 8027 18949 8113 19005
rect 8169 18949 8255 19005
rect 8311 18949 8397 19005
rect 8453 18949 8539 19005
rect 8595 18949 8681 19005
rect 8737 18949 8823 19005
rect 8879 18949 8965 19005
rect 9021 18949 9107 19005
rect 9163 18949 9249 19005
rect 9305 18949 9391 19005
rect 9447 18949 9533 19005
rect 9589 18949 9675 19005
rect 9731 18949 9817 19005
rect 9873 18949 9959 19005
rect 10015 18949 10101 19005
rect 10157 18949 10243 19005
rect 10299 18949 10385 19005
rect 10441 18949 10527 19005
rect 10583 18949 10669 19005
rect 10725 18949 10811 19005
rect 10867 18949 10953 19005
rect 11009 18949 11095 19005
rect 11151 18949 11237 19005
rect 11293 18949 11379 19005
rect 11435 18949 11521 19005
rect 11577 18949 11663 19005
rect 11719 18949 11805 19005
rect 11861 18949 11947 19005
rect 12003 18949 12089 19005
rect 12145 18949 12231 19005
rect 12287 18949 12373 19005
rect 12429 18949 12515 19005
rect 12571 18949 12657 19005
rect 12713 18949 12799 19005
rect 12855 18949 12941 19005
rect 12997 18949 13083 19005
rect 13139 18949 13225 19005
rect 13281 18949 13367 19005
rect 13423 18949 13509 19005
rect 13565 18949 13651 19005
rect 13707 18949 13793 19005
rect 13849 18949 13935 19005
rect 13991 18949 14077 19005
rect 14133 18949 14219 19005
rect 14275 18949 14361 19005
rect 14417 18949 14503 19005
rect 14559 18949 14645 19005
rect 14701 18949 14787 19005
rect 14843 18949 15000 19005
rect 0 18863 15000 18949
rect 0 18807 161 18863
rect 217 18807 303 18863
rect 359 18807 445 18863
rect 501 18807 587 18863
rect 643 18807 729 18863
rect 785 18807 871 18863
rect 927 18807 1013 18863
rect 1069 18807 1155 18863
rect 1211 18807 1297 18863
rect 1353 18807 1439 18863
rect 1495 18807 1581 18863
rect 1637 18807 1723 18863
rect 1779 18807 1865 18863
rect 1921 18807 2007 18863
rect 2063 18807 2149 18863
rect 2205 18807 2291 18863
rect 2347 18807 2433 18863
rect 2489 18807 2575 18863
rect 2631 18807 2717 18863
rect 2773 18807 2859 18863
rect 2915 18807 3001 18863
rect 3057 18807 3143 18863
rect 3199 18807 3285 18863
rect 3341 18807 3427 18863
rect 3483 18807 3569 18863
rect 3625 18807 3711 18863
rect 3767 18807 3853 18863
rect 3909 18807 3995 18863
rect 4051 18807 4137 18863
rect 4193 18807 4279 18863
rect 4335 18807 4421 18863
rect 4477 18807 4563 18863
rect 4619 18807 4705 18863
rect 4761 18807 4847 18863
rect 4903 18807 4989 18863
rect 5045 18807 5131 18863
rect 5187 18807 5273 18863
rect 5329 18807 5415 18863
rect 5471 18807 5557 18863
rect 5613 18807 5699 18863
rect 5755 18807 5841 18863
rect 5897 18807 5983 18863
rect 6039 18807 6125 18863
rect 6181 18807 6267 18863
rect 6323 18807 6409 18863
rect 6465 18807 6551 18863
rect 6607 18807 6693 18863
rect 6749 18807 6835 18863
rect 6891 18807 6977 18863
rect 7033 18807 7119 18863
rect 7175 18807 7261 18863
rect 7317 18807 7403 18863
rect 7459 18807 7545 18863
rect 7601 18807 7687 18863
rect 7743 18807 7829 18863
rect 7885 18807 7971 18863
rect 8027 18807 8113 18863
rect 8169 18807 8255 18863
rect 8311 18807 8397 18863
rect 8453 18807 8539 18863
rect 8595 18807 8681 18863
rect 8737 18807 8823 18863
rect 8879 18807 8965 18863
rect 9021 18807 9107 18863
rect 9163 18807 9249 18863
rect 9305 18807 9391 18863
rect 9447 18807 9533 18863
rect 9589 18807 9675 18863
rect 9731 18807 9817 18863
rect 9873 18807 9959 18863
rect 10015 18807 10101 18863
rect 10157 18807 10243 18863
rect 10299 18807 10385 18863
rect 10441 18807 10527 18863
rect 10583 18807 10669 18863
rect 10725 18807 10811 18863
rect 10867 18807 10953 18863
rect 11009 18807 11095 18863
rect 11151 18807 11237 18863
rect 11293 18807 11379 18863
rect 11435 18807 11521 18863
rect 11577 18807 11663 18863
rect 11719 18807 11805 18863
rect 11861 18807 11947 18863
rect 12003 18807 12089 18863
rect 12145 18807 12231 18863
rect 12287 18807 12373 18863
rect 12429 18807 12515 18863
rect 12571 18807 12657 18863
rect 12713 18807 12799 18863
rect 12855 18807 12941 18863
rect 12997 18807 13083 18863
rect 13139 18807 13225 18863
rect 13281 18807 13367 18863
rect 13423 18807 13509 18863
rect 13565 18807 13651 18863
rect 13707 18807 13793 18863
rect 13849 18807 13935 18863
rect 13991 18807 14077 18863
rect 14133 18807 14219 18863
rect 14275 18807 14361 18863
rect 14417 18807 14503 18863
rect 14559 18807 14645 18863
rect 14701 18807 14787 18863
rect 14843 18807 15000 18863
rect 0 18721 15000 18807
rect 0 18665 161 18721
rect 217 18665 303 18721
rect 359 18665 445 18721
rect 501 18665 587 18721
rect 643 18665 729 18721
rect 785 18665 871 18721
rect 927 18665 1013 18721
rect 1069 18665 1155 18721
rect 1211 18665 1297 18721
rect 1353 18665 1439 18721
rect 1495 18665 1581 18721
rect 1637 18665 1723 18721
rect 1779 18665 1865 18721
rect 1921 18665 2007 18721
rect 2063 18665 2149 18721
rect 2205 18665 2291 18721
rect 2347 18665 2433 18721
rect 2489 18665 2575 18721
rect 2631 18665 2717 18721
rect 2773 18665 2859 18721
rect 2915 18665 3001 18721
rect 3057 18665 3143 18721
rect 3199 18665 3285 18721
rect 3341 18665 3427 18721
rect 3483 18665 3569 18721
rect 3625 18665 3711 18721
rect 3767 18665 3853 18721
rect 3909 18665 3995 18721
rect 4051 18665 4137 18721
rect 4193 18665 4279 18721
rect 4335 18665 4421 18721
rect 4477 18665 4563 18721
rect 4619 18665 4705 18721
rect 4761 18665 4847 18721
rect 4903 18665 4989 18721
rect 5045 18665 5131 18721
rect 5187 18665 5273 18721
rect 5329 18665 5415 18721
rect 5471 18665 5557 18721
rect 5613 18665 5699 18721
rect 5755 18665 5841 18721
rect 5897 18665 5983 18721
rect 6039 18665 6125 18721
rect 6181 18665 6267 18721
rect 6323 18665 6409 18721
rect 6465 18665 6551 18721
rect 6607 18665 6693 18721
rect 6749 18665 6835 18721
rect 6891 18665 6977 18721
rect 7033 18665 7119 18721
rect 7175 18665 7261 18721
rect 7317 18665 7403 18721
rect 7459 18665 7545 18721
rect 7601 18665 7687 18721
rect 7743 18665 7829 18721
rect 7885 18665 7971 18721
rect 8027 18665 8113 18721
rect 8169 18665 8255 18721
rect 8311 18665 8397 18721
rect 8453 18665 8539 18721
rect 8595 18665 8681 18721
rect 8737 18665 8823 18721
rect 8879 18665 8965 18721
rect 9021 18665 9107 18721
rect 9163 18665 9249 18721
rect 9305 18665 9391 18721
rect 9447 18665 9533 18721
rect 9589 18665 9675 18721
rect 9731 18665 9817 18721
rect 9873 18665 9959 18721
rect 10015 18665 10101 18721
rect 10157 18665 10243 18721
rect 10299 18665 10385 18721
rect 10441 18665 10527 18721
rect 10583 18665 10669 18721
rect 10725 18665 10811 18721
rect 10867 18665 10953 18721
rect 11009 18665 11095 18721
rect 11151 18665 11237 18721
rect 11293 18665 11379 18721
rect 11435 18665 11521 18721
rect 11577 18665 11663 18721
rect 11719 18665 11805 18721
rect 11861 18665 11947 18721
rect 12003 18665 12089 18721
rect 12145 18665 12231 18721
rect 12287 18665 12373 18721
rect 12429 18665 12515 18721
rect 12571 18665 12657 18721
rect 12713 18665 12799 18721
rect 12855 18665 12941 18721
rect 12997 18665 13083 18721
rect 13139 18665 13225 18721
rect 13281 18665 13367 18721
rect 13423 18665 13509 18721
rect 13565 18665 13651 18721
rect 13707 18665 13793 18721
rect 13849 18665 13935 18721
rect 13991 18665 14077 18721
rect 14133 18665 14219 18721
rect 14275 18665 14361 18721
rect 14417 18665 14503 18721
rect 14559 18665 14645 18721
rect 14701 18665 14787 18721
rect 14843 18665 15000 18721
rect 0 18579 15000 18665
rect 0 18523 161 18579
rect 217 18523 303 18579
rect 359 18523 445 18579
rect 501 18523 587 18579
rect 643 18523 729 18579
rect 785 18523 871 18579
rect 927 18523 1013 18579
rect 1069 18523 1155 18579
rect 1211 18523 1297 18579
rect 1353 18523 1439 18579
rect 1495 18523 1581 18579
rect 1637 18523 1723 18579
rect 1779 18523 1865 18579
rect 1921 18523 2007 18579
rect 2063 18523 2149 18579
rect 2205 18523 2291 18579
rect 2347 18523 2433 18579
rect 2489 18523 2575 18579
rect 2631 18523 2717 18579
rect 2773 18523 2859 18579
rect 2915 18523 3001 18579
rect 3057 18523 3143 18579
rect 3199 18523 3285 18579
rect 3341 18523 3427 18579
rect 3483 18523 3569 18579
rect 3625 18523 3711 18579
rect 3767 18523 3853 18579
rect 3909 18523 3995 18579
rect 4051 18523 4137 18579
rect 4193 18523 4279 18579
rect 4335 18523 4421 18579
rect 4477 18523 4563 18579
rect 4619 18523 4705 18579
rect 4761 18523 4847 18579
rect 4903 18523 4989 18579
rect 5045 18523 5131 18579
rect 5187 18523 5273 18579
rect 5329 18523 5415 18579
rect 5471 18523 5557 18579
rect 5613 18523 5699 18579
rect 5755 18523 5841 18579
rect 5897 18523 5983 18579
rect 6039 18523 6125 18579
rect 6181 18523 6267 18579
rect 6323 18523 6409 18579
rect 6465 18523 6551 18579
rect 6607 18523 6693 18579
rect 6749 18523 6835 18579
rect 6891 18523 6977 18579
rect 7033 18523 7119 18579
rect 7175 18523 7261 18579
rect 7317 18523 7403 18579
rect 7459 18523 7545 18579
rect 7601 18523 7687 18579
rect 7743 18523 7829 18579
rect 7885 18523 7971 18579
rect 8027 18523 8113 18579
rect 8169 18523 8255 18579
rect 8311 18523 8397 18579
rect 8453 18523 8539 18579
rect 8595 18523 8681 18579
rect 8737 18523 8823 18579
rect 8879 18523 8965 18579
rect 9021 18523 9107 18579
rect 9163 18523 9249 18579
rect 9305 18523 9391 18579
rect 9447 18523 9533 18579
rect 9589 18523 9675 18579
rect 9731 18523 9817 18579
rect 9873 18523 9959 18579
rect 10015 18523 10101 18579
rect 10157 18523 10243 18579
rect 10299 18523 10385 18579
rect 10441 18523 10527 18579
rect 10583 18523 10669 18579
rect 10725 18523 10811 18579
rect 10867 18523 10953 18579
rect 11009 18523 11095 18579
rect 11151 18523 11237 18579
rect 11293 18523 11379 18579
rect 11435 18523 11521 18579
rect 11577 18523 11663 18579
rect 11719 18523 11805 18579
rect 11861 18523 11947 18579
rect 12003 18523 12089 18579
rect 12145 18523 12231 18579
rect 12287 18523 12373 18579
rect 12429 18523 12515 18579
rect 12571 18523 12657 18579
rect 12713 18523 12799 18579
rect 12855 18523 12941 18579
rect 12997 18523 13083 18579
rect 13139 18523 13225 18579
rect 13281 18523 13367 18579
rect 13423 18523 13509 18579
rect 13565 18523 13651 18579
rect 13707 18523 13793 18579
rect 13849 18523 13935 18579
rect 13991 18523 14077 18579
rect 14133 18523 14219 18579
rect 14275 18523 14361 18579
rect 14417 18523 14503 18579
rect 14559 18523 14645 18579
rect 14701 18523 14787 18579
rect 14843 18523 15000 18579
rect 0 18437 15000 18523
rect 0 18381 161 18437
rect 217 18381 303 18437
rect 359 18381 445 18437
rect 501 18381 587 18437
rect 643 18381 729 18437
rect 785 18381 871 18437
rect 927 18381 1013 18437
rect 1069 18381 1155 18437
rect 1211 18381 1297 18437
rect 1353 18381 1439 18437
rect 1495 18381 1581 18437
rect 1637 18381 1723 18437
rect 1779 18381 1865 18437
rect 1921 18381 2007 18437
rect 2063 18381 2149 18437
rect 2205 18381 2291 18437
rect 2347 18381 2433 18437
rect 2489 18381 2575 18437
rect 2631 18381 2717 18437
rect 2773 18381 2859 18437
rect 2915 18381 3001 18437
rect 3057 18381 3143 18437
rect 3199 18381 3285 18437
rect 3341 18381 3427 18437
rect 3483 18381 3569 18437
rect 3625 18381 3711 18437
rect 3767 18381 3853 18437
rect 3909 18381 3995 18437
rect 4051 18381 4137 18437
rect 4193 18381 4279 18437
rect 4335 18381 4421 18437
rect 4477 18381 4563 18437
rect 4619 18381 4705 18437
rect 4761 18381 4847 18437
rect 4903 18381 4989 18437
rect 5045 18381 5131 18437
rect 5187 18381 5273 18437
rect 5329 18381 5415 18437
rect 5471 18381 5557 18437
rect 5613 18381 5699 18437
rect 5755 18381 5841 18437
rect 5897 18381 5983 18437
rect 6039 18381 6125 18437
rect 6181 18381 6267 18437
rect 6323 18381 6409 18437
rect 6465 18381 6551 18437
rect 6607 18381 6693 18437
rect 6749 18381 6835 18437
rect 6891 18381 6977 18437
rect 7033 18381 7119 18437
rect 7175 18381 7261 18437
rect 7317 18381 7403 18437
rect 7459 18381 7545 18437
rect 7601 18381 7687 18437
rect 7743 18381 7829 18437
rect 7885 18381 7971 18437
rect 8027 18381 8113 18437
rect 8169 18381 8255 18437
rect 8311 18381 8397 18437
rect 8453 18381 8539 18437
rect 8595 18381 8681 18437
rect 8737 18381 8823 18437
rect 8879 18381 8965 18437
rect 9021 18381 9107 18437
rect 9163 18381 9249 18437
rect 9305 18381 9391 18437
rect 9447 18381 9533 18437
rect 9589 18381 9675 18437
rect 9731 18381 9817 18437
rect 9873 18381 9959 18437
rect 10015 18381 10101 18437
rect 10157 18381 10243 18437
rect 10299 18381 10385 18437
rect 10441 18381 10527 18437
rect 10583 18381 10669 18437
rect 10725 18381 10811 18437
rect 10867 18381 10953 18437
rect 11009 18381 11095 18437
rect 11151 18381 11237 18437
rect 11293 18381 11379 18437
rect 11435 18381 11521 18437
rect 11577 18381 11663 18437
rect 11719 18381 11805 18437
rect 11861 18381 11947 18437
rect 12003 18381 12089 18437
rect 12145 18381 12231 18437
rect 12287 18381 12373 18437
rect 12429 18381 12515 18437
rect 12571 18381 12657 18437
rect 12713 18381 12799 18437
rect 12855 18381 12941 18437
rect 12997 18381 13083 18437
rect 13139 18381 13225 18437
rect 13281 18381 13367 18437
rect 13423 18381 13509 18437
rect 13565 18381 13651 18437
rect 13707 18381 13793 18437
rect 13849 18381 13935 18437
rect 13991 18381 14077 18437
rect 14133 18381 14219 18437
rect 14275 18381 14361 18437
rect 14417 18381 14503 18437
rect 14559 18381 14645 18437
rect 14701 18381 14787 18437
rect 14843 18381 15000 18437
rect 0 18295 15000 18381
rect 0 18239 161 18295
rect 217 18239 303 18295
rect 359 18239 445 18295
rect 501 18239 587 18295
rect 643 18239 729 18295
rect 785 18239 871 18295
rect 927 18239 1013 18295
rect 1069 18239 1155 18295
rect 1211 18239 1297 18295
rect 1353 18239 1439 18295
rect 1495 18239 1581 18295
rect 1637 18239 1723 18295
rect 1779 18239 1865 18295
rect 1921 18239 2007 18295
rect 2063 18239 2149 18295
rect 2205 18239 2291 18295
rect 2347 18239 2433 18295
rect 2489 18239 2575 18295
rect 2631 18239 2717 18295
rect 2773 18239 2859 18295
rect 2915 18239 3001 18295
rect 3057 18239 3143 18295
rect 3199 18239 3285 18295
rect 3341 18239 3427 18295
rect 3483 18239 3569 18295
rect 3625 18239 3711 18295
rect 3767 18239 3853 18295
rect 3909 18239 3995 18295
rect 4051 18239 4137 18295
rect 4193 18239 4279 18295
rect 4335 18239 4421 18295
rect 4477 18239 4563 18295
rect 4619 18239 4705 18295
rect 4761 18239 4847 18295
rect 4903 18239 4989 18295
rect 5045 18239 5131 18295
rect 5187 18239 5273 18295
rect 5329 18239 5415 18295
rect 5471 18239 5557 18295
rect 5613 18239 5699 18295
rect 5755 18239 5841 18295
rect 5897 18239 5983 18295
rect 6039 18239 6125 18295
rect 6181 18239 6267 18295
rect 6323 18239 6409 18295
rect 6465 18239 6551 18295
rect 6607 18239 6693 18295
rect 6749 18239 6835 18295
rect 6891 18239 6977 18295
rect 7033 18239 7119 18295
rect 7175 18239 7261 18295
rect 7317 18239 7403 18295
rect 7459 18239 7545 18295
rect 7601 18239 7687 18295
rect 7743 18239 7829 18295
rect 7885 18239 7971 18295
rect 8027 18239 8113 18295
rect 8169 18239 8255 18295
rect 8311 18239 8397 18295
rect 8453 18239 8539 18295
rect 8595 18239 8681 18295
rect 8737 18239 8823 18295
rect 8879 18239 8965 18295
rect 9021 18239 9107 18295
rect 9163 18239 9249 18295
rect 9305 18239 9391 18295
rect 9447 18239 9533 18295
rect 9589 18239 9675 18295
rect 9731 18239 9817 18295
rect 9873 18239 9959 18295
rect 10015 18239 10101 18295
rect 10157 18239 10243 18295
rect 10299 18239 10385 18295
rect 10441 18239 10527 18295
rect 10583 18239 10669 18295
rect 10725 18239 10811 18295
rect 10867 18239 10953 18295
rect 11009 18239 11095 18295
rect 11151 18239 11237 18295
rect 11293 18239 11379 18295
rect 11435 18239 11521 18295
rect 11577 18239 11663 18295
rect 11719 18239 11805 18295
rect 11861 18239 11947 18295
rect 12003 18239 12089 18295
rect 12145 18239 12231 18295
rect 12287 18239 12373 18295
rect 12429 18239 12515 18295
rect 12571 18239 12657 18295
rect 12713 18239 12799 18295
rect 12855 18239 12941 18295
rect 12997 18239 13083 18295
rect 13139 18239 13225 18295
rect 13281 18239 13367 18295
rect 13423 18239 13509 18295
rect 13565 18239 13651 18295
rect 13707 18239 13793 18295
rect 13849 18239 13935 18295
rect 13991 18239 14077 18295
rect 14133 18239 14219 18295
rect 14275 18239 14361 18295
rect 14417 18239 14503 18295
rect 14559 18239 14645 18295
rect 14701 18239 14787 18295
rect 14843 18239 15000 18295
rect 0 18153 15000 18239
rect 0 18097 161 18153
rect 217 18097 303 18153
rect 359 18097 445 18153
rect 501 18097 587 18153
rect 643 18097 729 18153
rect 785 18097 871 18153
rect 927 18097 1013 18153
rect 1069 18097 1155 18153
rect 1211 18097 1297 18153
rect 1353 18097 1439 18153
rect 1495 18097 1581 18153
rect 1637 18097 1723 18153
rect 1779 18097 1865 18153
rect 1921 18097 2007 18153
rect 2063 18097 2149 18153
rect 2205 18097 2291 18153
rect 2347 18097 2433 18153
rect 2489 18097 2575 18153
rect 2631 18097 2717 18153
rect 2773 18097 2859 18153
rect 2915 18097 3001 18153
rect 3057 18097 3143 18153
rect 3199 18097 3285 18153
rect 3341 18097 3427 18153
rect 3483 18097 3569 18153
rect 3625 18097 3711 18153
rect 3767 18097 3853 18153
rect 3909 18097 3995 18153
rect 4051 18097 4137 18153
rect 4193 18097 4279 18153
rect 4335 18097 4421 18153
rect 4477 18097 4563 18153
rect 4619 18097 4705 18153
rect 4761 18097 4847 18153
rect 4903 18097 4989 18153
rect 5045 18097 5131 18153
rect 5187 18097 5273 18153
rect 5329 18097 5415 18153
rect 5471 18097 5557 18153
rect 5613 18097 5699 18153
rect 5755 18097 5841 18153
rect 5897 18097 5983 18153
rect 6039 18097 6125 18153
rect 6181 18097 6267 18153
rect 6323 18097 6409 18153
rect 6465 18097 6551 18153
rect 6607 18097 6693 18153
rect 6749 18097 6835 18153
rect 6891 18097 6977 18153
rect 7033 18097 7119 18153
rect 7175 18097 7261 18153
rect 7317 18097 7403 18153
rect 7459 18097 7545 18153
rect 7601 18097 7687 18153
rect 7743 18097 7829 18153
rect 7885 18097 7971 18153
rect 8027 18097 8113 18153
rect 8169 18097 8255 18153
rect 8311 18097 8397 18153
rect 8453 18097 8539 18153
rect 8595 18097 8681 18153
rect 8737 18097 8823 18153
rect 8879 18097 8965 18153
rect 9021 18097 9107 18153
rect 9163 18097 9249 18153
rect 9305 18097 9391 18153
rect 9447 18097 9533 18153
rect 9589 18097 9675 18153
rect 9731 18097 9817 18153
rect 9873 18097 9959 18153
rect 10015 18097 10101 18153
rect 10157 18097 10243 18153
rect 10299 18097 10385 18153
rect 10441 18097 10527 18153
rect 10583 18097 10669 18153
rect 10725 18097 10811 18153
rect 10867 18097 10953 18153
rect 11009 18097 11095 18153
rect 11151 18097 11237 18153
rect 11293 18097 11379 18153
rect 11435 18097 11521 18153
rect 11577 18097 11663 18153
rect 11719 18097 11805 18153
rect 11861 18097 11947 18153
rect 12003 18097 12089 18153
rect 12145 18097 12231 18153
rect 12287 18097 12373 18153
rect 12429 18097 12515 18153
rect 12571 18097 12657 18153
rect 12713 18097 12799 18153
rect 12855 18097 12941 18153
rect 12997 18097 13083 18153
rect 13139 18097 13225 18153
rect 13281 18097 13367 18153
rect 13423 18097 13509 18153
rect 13565 18097 13651 18153
rect 13707 18097 13793 18153
rect 13849 18097 13935 18153
rect 13991 18097 14077 18153
rect 14133 18097 14219 18153
rect 14275 18097 14361 18153
rect 14417 18097 14503 18153
rect 14559 18097 14645 18153
rect 14701 18097 14787 18153
rect 14843 18097 15000 18153
rect 0 18011 15000 18097
rect 0 17955 161 18011
rect 217 17955 303 18011
rect 359 17955 445 18011
rect 501 17955 587 18011
rect 643 17955 729 18011
rect 785 17955 871 18011
rect 927 17955 1013 18011
rect 1069 17955 1155 18011
rect 1211 17955 1297 18011
rect 1353 17955 1439 18011
rect 1495 17955 1581 18011
rect 1637 17955 1723 18011
rect 1779 17955 1865 18011
rect 1921 17955 2007 18011
rect 2063 17955 2149 18011
rect 2205 17955 2291 18011
rect 2347 17955 2433 18011
rect 2489 17955 2575 18011
rect 2631 17955 2717 18011
rect 2773 17955 2859 18011
rect 2915 17955 3001 18011
rect 3057 17955 3143 18011
rect 3199 17955 3285 18011
rect 3341 17955 3427 18011
rect 3483 17955 3569 18011
rect 3625 17955 3711 18011
rect 3767 17955 3853 18011
rect 3909 17955 3995 18011
rect 4051 17955 4137 18011
rect 4193 17955 4279 18011
rect 4335 17955 4421 18011
rect 4477 17955 4563 18011
rect 4619 17955 4705 18011
rect 4761 17955 4847 18011
rect 4903 17955 4989 18011
rect 5045 17955 5131 18011
rect 5187 17955 5273 18011
rect 5329 17955 5415 18011
rect 5471 17955 5557 18011
rect 5613 17955 5699 18011
rect 5755 17955 5841 18011
rect 5897 17955 5983 18011
rect 6039 17955 6125 18011
rect 6181 17955 6267 18011
rect 6323 17955 6409 18011
rect 6465 17955 6551 18011
rect 6607 17955 6693 18011
rect 6749 17955 6835 18011
rect 6891 17955 6977 18011
rect 7033 17955 7119 18011
rect 7175 17955 7261 18011
rect 7317 17955 7403 18011
rect 7459 17955 7545 18011
rect 7601 17955 7687 18011
rect 7743 17955 7829 18011
rect 7885 17955 7971 18011
rect 8027 17955 8113 18011
rect 8169 17955 8255 18011
rect 8311 17955 8397 18011
rect 8453 17955 8539 18011
rect 8595 17955 8681 18011
rect 8737 17955 8823 18011
rect 8879 17955 8965 18011
rect 9021 17955 9107 18011
rect 9163 17955 9249 18011
rect 9305 17955 9391 18011
rect 9447 17955 9533 18011
rect 9589 17955 9675 18011
rect 9731 17955 9817 18011
rect 9873 17955 9959 18011
rect 10015 17955 10101 18011
rect 10157 17955 10243 18011
rect 10299 17955 10385 18011
rect 10441 17955 10527 18011
rect 10583 17955 10669 18011
rect 10725 17955 10811 18011
rect 10867 17955 10953 18011
rect 11009 17955 11095 18011
rect 11151 17955 11237 18011
rect 11293 17955 11379 18011
rect 11435 17955 11521 18011
rect 11577 17955 11663 18011
rect 11719 17955 11805 18011
rect 11861 17955 11947 18011
rect 12003 17955 12089 18011
rect 12145 17955 12231 18011
rect 12287 17955 12373 18011
rect 12429 17955 12515 18011
rect 12571 17955 12657 18011
rect 12713 17955 12799 18011
rect 12855 17955 12941 18011
rect 12997 17955 13083 18011
rect 13139 17955 13225 18011
rect 13281 17955 13367 18011
rect 13423 17955 13509 18011
rect 13565 17955 13651 18011
rect 13707 17955 13793 18011
rect 13849 17955 13935 18011
rect 13991 17955 14077 18011
rect 14133 17955 14219 18011
rect 14275 17955 14361 18011
rect 14417 17955 14503 18011
rect 14559 17955 14645 18011
rect 14701 17955 14787 18011
rect 14843 17955 15000 18011
rect 0 17869 15000 17955
rect 0 17813 161 17869
rect 217 17813 303 17869
rect 359 17813 445 17869
rect 501 17813 587 17869
rect 643 17813 729 17869
rect 785 17813 871 17869
rect 927 17813 1013 17869
rect 1069 17813 1155 17869
rect 1211 17813 1297 17869
rect 1353 17813 1439 17869
rect 1495 17813 1581 17869
rect 1637 17813 1723 17869
rect 1779 17813 1865 17869
rect 1921 17813 2007 17869
rect 2063 17813 2149 17869
rect 2205 17813 2291 17869
rect 2347 17813 2433 17869
rect 2489 17813 2575 17869
rect 2631 17813 2717 17869
rect 2773 17813 2859 17869
rect 2915 17813 3001 17869
rect 3057 17813 3143 17869
rect 3199 17813 3285 17869
rect 3341 17813 3427 17869
rect 3483 17813 3569 17869
rect 3625 17813 3711 17869
rect 3767 17813 3853 17869
rect 3909 17813 3995 17869
rect 4051 17813 4137 17869
rect 4193 17813 4279 17869
rect 4335 17813 4421 17869
rect 4477 17813 4563 17869
rect 4619 17813 4705 17869
rect 4761 17813 4847 17869
rect 4903 17813 4989 17869
rect 5045 17813 5131 17869
rect 5187 17813 5273 17869
rect 5329 17813 5415 17869
rect 5471 17813 5557 17869
rect 5613 17813 5699 17869
rect 5755 17813 5841 17869
rect 5897 17813 5983 17869
rect 6039 17813 6125 17869
rect 6181 17813 6267 17869
rect 6323 17813 6409 17869
rect 6465 17813 6551 17869
rect 6607 17813 6693 17869
rect 6749 17813 6835 17869
rect 6891 17813 6977 17869
rect 7033 17813 7119 17869
rect 7175 17813 7261 17869
rect 7317 17813 7403 17869
rect 7459 17813 7545 17869
rect 7601 17813 7687 17869
rect 7743 17813 7829 17869
rect 7885 17813 7971 17869
rect 8027 17813 8113 17869
rect 8169 17813 8255 17869
rect 8311 17813 8397 17869
rect 8453 17813 8539 17869
rect 8595 17813 8681 17869
rect 8737 17813 8823 17869
rect 8879 17813 8965 17869
rect 9021 17813 9107 17869
rect 9163 17813 9249 17869
rect 9305 17813 9391 17869
rect 9447 17813 9533 17869
rect 9589 17813 9675 17869
rect 9731 17813 9817 17869
rect 9873 17813 9959 17869
rect 10015 17813 10101 17869
rect 10157 17813 10243 17869
rect 10299 17813 10385 17869
rect 10441 17813 10527 17869
rect 10583 17813 10669 17869
rect 10725 17813 10811 17869
rect 10867 17813 10953 17869
rect 11009 17813 11095 17869
rect 11151 17813 11237 17869
rect 11293 17813 11379 17869
rect 11435 17813 11521 17869
rect 11577 17813 11663 17869
rect 11719 17813 11805 17869
rect 11861 17813 11947 17869
rect 12003 17813 12089 17869
rect 12145 17813 12231 17869
rect 12287 17813 12373 17869
rect 12429 17813 12515 17869
rect 12571 17813 12657 17869
rect 12713 17813 12799 17869
rect 12855 17813 12941 17869
rect 12997 17813 13083 17869
rect 13139 17813 13225 17869
rect 13281 17813 13367 17869
rect 13423 17813 13509 17869
rect 13565 17813 13651 17869
rect 13707 17813 13793 17869
rect 13849 17813 13935 17869
rect 13991 17813 14077 17869
rect 14133 17813 14219 17869
rect 14275 17813 14361 17869
rect 14417 17813 14503 17869
rect 14559 17813 14645 17869
rect 14701 17813 14787 17869
rect 14843 17813 15000 17869
rect 0 17727 15000 17813
rect 0 17671 161 17727
rect 217 17671 303 17727
rect 359 17671 445 17727
rect 501 17671 587 17727
rect 643 17671 729 17727
rect 785 17671 871 17727
rect 927 17671 1013 17727
rect 1069 17671 1155 17727
rect 1211 17671 1297 17727
rect 1353 17671 1439 17727
rect 1495 17671 1581 17727
rect 1637 17671 1723 17727
rect 1779 17671 1865 17727
rect 1921 17671 2007 17727
rect 2063 17671 2149 17727
rect 2205 17671 2291 17727
rect 2347 17671 2433 17727
rect 2489 17671 2575 17727
rect 2631 17671 2717 17727
rect 2773 17671 2859 17727
rect 2915 17671 3001 17727
rect 3057 17671 3143 17727
rect 3199 17671 3285 17727
rect 3341 17671 3427 17727
rect 3483 17671 3569 17727
rect 3625 17671 3711 17727
rect 3767 17671 3853 17727
rect 3909 17671 3995 17727
rect 4051 17671 4137 17727
rect 4193 17671 4279 17727
rect 4335 17671 4421 17727
rect 4477 17671 4563 17727
rect 4619 17671 4705 17727
rect 4761 17671 4847 17727
rect 4903 17671 4989 17727
rect 5045 17671 5131 17727
rect 5187 17671 5273 17727
rect 5329 17671 5415 17727
rect 5471 17671 5557 17727
rect 5613 17671 5699 17727
rect 5755 17671 5841 17727
rect 5897 17671 5983 17727
rect 6039 17671 6125 17727
rect 6181 17671 6267 17727
rect 6323 17671 6409 17727
rect 6465 17671 6551 17727
rect 6607 17671 6693 17727
rect 6749 17671 6835 17727
rect 6891 17671 6977 17727
rect 7033 17671 7119 17727
rect 7175 17671 7261 17727
rect 7317 17671 7403 17727
rect 7459 17671 7545 17727
rect 7601 17671 7687 17727
rect 7743 17671 7829 17727
rect 7885 17671 7971 17727
rect 8027 17671 8113 17727
rect 8169 17671 8255 17727
rect 8311 17671 8397 17727
rect 8453 17671 8539 17727
rect 8595 17671 8681 17727
rect 8737 17671 8823 17727
rect 8879 17671 8965 17727
rect 9021 17671 9107 17727
rect 9163 17671 9249 17727
rect 9305 17671 9391 17727
rect 9447 17671 9533 17727
rect 9589 17671 9675 17727
rect 9731 17671 9817 17727
rect 9873 17671 9959 17727
rect 10015 17671 10101 17727
rect 10157 17671 10243 17727
rect 10299 17671 10385 17727
rect 10441 17671 10527 17727
rect 10583 17671 10669 17727
rect 10725 17671 10811 17727
rect 10867 17671 10953 17727
rect 11009 17671 11095 17727
rect 11151 17671 11237 17727
rect 11293 17671 11379 17727
rect 11435 17671 11521 17727
rect 11577 17671 11663 17727
rect 11719 17671 11805 17727
rect 11861 17671 11947 17727
rect 12003 17671 12089 17727
rect 12145 17671 12231 17727
rect 12287 17671 12373 17727
rect 12429 17671 12515 17727
rect 12571 17671 12657 17727
rect 12713 17671 12799 17727
rect 12855 17671 12941 17727
rect 12997 17671 13083 17727
rect 13139 17671 13225 17727
rect 13281 17671 13367 17727
rect 13423 17671 13509 17727
rect 13565 17671 13651 17727
rect 13707 17671 13793 17727
rect 13849 17671 13935 17727
rect 13991 17671 14077 17727
rect 14133 17671 14219 17727
rect 14275 17671 14361 17727
rect 14417 17671 14503 17727
rect 14559 17671 14645 17727
rect 14701 17671 14787 17727
rect 14843 17671 15000 17727
rect 0 17585 15000 17671
rect 0 17529 161 17585
rect 217 17529 303 17585
rect 359 17529 445 17585
rect 501 17529 587 17585
rect 643 17529 729 17585
rect 785 17529 871 17585
rect 927 17529 1013 17585
rect 1069 17529 1155 17585
rect 1211 17529 1297 17585
rect 1353 17529 1439 17585
rect 1495 17529 1581 17585
rect 1637 17529 1723 17585
rect 1779 17529 1865 17585
rect 1921 17529 2007 17585
rect 2063 17529 2149 17585
rect 2205 17529 2291 17585
rect 2347 17529 2433 17585
rect 2489 17529 2575 17585
rect 2631 17529 2717 17585
rect 2773 17529 2859 17585
rect 2915 17529 3001 17585
rect 3057 17529 3143 17585
rect 3199 17529 3285 17585
rect 3341 17529 3427 17585
rect 3483 17529 3569 17585
rect 3625 17529 3711 17585
rect 3767 17529 3853 17585
rect 3909 17529 3995 17585
rect 4051 17529 4137 17585
rect 4193 17529 4279 17585
rect 4335 17529 4421 17585
rect 4477 17529 4563 17585
rect 4619 17529 4705 17585
rect 4761 17529 4847 17585
rect 4903 17529 4989 17585
rect 5045 17529 5131 17585
rect 5187 17529 5273 17585
rect 5329 17529 5415 17585
rect 5471 17529 5557 17585
rect 5613 17529 5699 17585
rect 5755 17529 5841 17585
rect 5897 17529 5983 17585
rect 6039 17529 6125 17585
rect 6181 17529 6267 17585
rect 6323 17529 6409 17585
rect 6465 17529 6551 17585
rect 6607 17529 6693 17585
rect 6749 17529 6835 17585
rect 6891 17529 6977 17585
rect 7033 17529 7119 17585
rect 7175 17529 7261 17585
rect 7317 17529 7403 17585
rect 7459 17529 7545 17585
rect 7601 17529 7687 17585
rect 7743 17529 7829 17585
rect 7885 17529 7971 17585
rect 8027 17529 8113 17585
rect 8169 17529 8255 17585
rect 8311 17529 8397 17585
rect 8453 17529 8539 17585
rect 8595 17529 8681 17585
rect 8737 17529 8823 17585
rect 8879 17529 8965 17585
rect 9021 17529 9107 17585
rect 9163 17529 9249 17585
rect 9305 17529 9391 17585
rect 9447 17529 9533 17585
rect 9589 17529 9675 17585
rect 9731 17529 9817 17585
rect 9873 17529 9959 17585
rect 10015 17529 10101 17585
rect 10157 17529 10243 17585
rect 10299 17529 10385 17585
rect 10441 17529 10527 17585
rect 10583 17529 10669 17585
rect 10725 17529 10811 17585
rect 10867 17529 10953 17585
rect 11009 17529 11095 17585
rect 11151 17529 11237 17585
rect 11293 17529 11379 17585
rect 11435 17529 11521 17585
rect 11577 17529 11663 17585
rect 11719 17529 11805 17585
rect 11861 17529 11947 17585
rect 12003 17529 12089 17585
rect 12145 17529 12231 17585
rect 12287 17529 12373 17585
rect 12429 17529 12515 17585
rect 12571 17529 12657 17585
rect 12713 17529 12799 17585
rect 12855 17529 12941 17585
rect 12997 17529 13083 17585
rect 13139 17529 13225 17585
rect 13281 17529 13367 17585
rect 13423 17529 13509 17585
rect 13565 17529 13651 17585
rect 13707 17529 13793 17585
rect 13849 17529 13935 17585
rect 13991 17529 14077 17585
rect 14133 17529 14219 17585
rect 14275 17529 14361 17585
rect 14417 17529 14503 17585
rect 14559 17529 14645 17585
rect 14701 17529 14787 17585
rect 14843 17529 15000 17585
rect 0 17443 15000 17529
rect 0 17387 161 17443
rect 217 17387 303 17443
rect 359 17387 445 17443
rect 501 17387 587 17443
rect 643 17387 729 17443
rect 785 17387 871 17443
rect 927 17387 1013 17443
rect 1069 17387 1155 17443
rect 1211 17387 1297 17443
rect 1353 17387 1439 17443
rect 1495 17387 1581 17443
rect 1637 17387 1723 17443
rect 1779 17387 1865 17443
rect 1921 17387 2007 17443
rect 2063 17387 2149 17443
rect 2205 17387 2291 17443
rect 2347 17387 2433 17443
rect 2489 17387 2575 17443
rect 2631 17387 2717 17443
rect 2773 17387 2859 17443
rect 2915 17387 3001 17443
rect 3057 17387 3143 17443
rect 3199 17387 3285 17443
rect 3341 17387 3427 17443
rect 3483 17387 3569 17443
rect 3625 17387 3711 17443
rect 3767 17387 3853 17443
rect 3909 17387 3995 17443
rect 4051 17387 4137 17443
rect 4193 17387 4279 17443
rect 4335 17387 4421 17443
rect 4477 17387 4563 17443
rect 4619 17387 4705 17443
rect 4761 17387 4847 17443
rect 4903 17387 4989 17443
rect 5045 17387 5131 17443
rect 5187 17387 5273 17443
rect 5329 17387 5415 17443
rect 5471 17387 5557 17443
rect 5613 17387 5699 17443
rect 5755 17387 5841 17443
rect 5897 17387 5983 17443
rect 6039 17387 6125 17443
rect 6181 17387 6267 17443
rect 6323 17387 6409 17443
rect 6465 17387 6551 17443
rect 6607 17387 6693 17443
rect 6749 17387 6835 17443
rect 6891 17387 6977 17443
rect 7033 17387 7119 17443
rect 7175 17387 7261 17443
rect 7317 17387 7403 17443
rect 7459 17387 7545 17443
rect 7601 17387 7687 17443
rect 7743 17387 7829 17443
rect 7885 17387 7971 17443
rect 8027 17387 8113 17443
rect 8169 17387 8255 17443
rect 8311 17387 8397 17443
rect 8453 17387 8539 17443
rect 8595 17387 8681 17443
rect 8737 17387 8823 17443
rect 8879 17387 8965 17443
rect 9021 17387 9107 17443
rect 9163 17387 9249 17443
rect 9305 17387 9391 17443
rect 9447 17387 9533 17443
rect 9589 17387 9675 17443
rect 9731 17387 9817 17443
rect 9873 17387 9959 17443
rect 10015 17387 10101 17443
rect 10157 17387 10243 17443
rect 10299 17387 10385 17443
rect 10441 17387 10527 17443
rect 10583 17387 10669 17443
rect 10725 17387 10811 17443
rect 10867 17387 10953 17443
rect 11009 17387 11095 17443
rect 11151 17387 11237 17443
rect 11293 17387 11379 17443
rect 11435 17387 11521 17443
rect 11577 17387 11663 17443
rect 11719 17387 11805 17443
rect 11861 17387 11947 17443
rect 12003 17387 12089 17443
rect 12145 17387 12231 17443
rect 12287 17387 12373 17443
rect 12429 17387 12515 17443
rect 12571 17387 12657 17443
rect 12713 17387 12799 17443
rect 12855 17387 12941 17443
rect 12997 17387 13083 17443
rect 13139 17387 13225 17443
rect 13281 17387 13367 17443
rect 13423 17387 13509 17443
rect 13565 17387 13651 17443
rect 13707 17387 13793 17443
rect 13849 17387 13935 17443
rect 13991 17387 14077 17443
rect 14133 17387 14219 17443
rect 14275 17387 14361 17443
rect 14417 17387 14503 17443
rect 14559 17387 14645 17443
rect 14701 17387 14787 17443
rect 14843 17387 15000 17443
rect 0 17301 15000 17387
rect 0 17245 161 17301
rect 217 17245 303 17301
rect 359 17245 445 17301
rect 501 17245 587 17301
rect 643 17245 729 17301
rect 785 17245 871 17301
rect 927 17245 1013 17301
rect 1069 17245 1155 17301
rect 1211 17245 1297 17301
rect 1353 17245 1439 17301
rect 1495 17245 1581 17301
rect 1637 17245 1723 17301
rect 1779 17245 1865 17301
rect 1921 17245 2007 17301
rect 2063 17245 2149 17301
rect 2205 17245 2291 17301
rect 2347 17245 2433 17301
rect 2489 17245 2575 17301
rect 2631 17245 2717 17301
rect 2773 17245 2859 17301
rect 2915 17245 3001 17301
rect 3057 17245 3143 17301
rect 3199 17245 3285 17301
rect 3341 17245 3427 17301
rect 3483 17245 3569 17301
rect 3625 17245 3711 17301
rect 3767 17245 3853 17301
rect 3909 17245 3995 17301
rect 4051 17245 4137 17301
rect 4193 17245 4279 17301
rect 4335 17245 4421 17301
rect 4477 17245 4563 17301
rect 4619 17245 4705 17301
rect 4761 17245 4847 17301
rect 4903 17245 4989 17301
rect 5045 17245 5131 17301
rect 5187 17245 5273 17301
rect 5329 17245 5415 17301
rect 5471 17245 5557 17301
rect 5613 17245 5699 17301
rect 5755 17245 5841 17301
rect 5897 17245 5983 17301
rect 6039 17245 6125 17301
rect 6181 17245 6267 17301
rect 6323 17245 6409 17301
rect 6465 17245 6551 17301
rect 6607 17245 6693 17301
rect 6749 17245 6835 17301
rect 6891 17245 6977 17301
rect 7033 17245 7119 17301
rect 7175 17245 7261 17301
rect 7317 17245 7403 17301
rect 7459 17245 7545 17301
rect 7601 17245 7687 17301
rect 7743 17245 7829 17301
rect 7885 17245 7971 17301
rect 8027 17245 8113 17301
rect 8169 17245 8255 17301
rect 8311 17245 8397 17301
rect 8453 17245 8539 17301
rect 8595 17245 8681 17301
rect 8737 17245 8823 17301
rect 8879 17245 8965 17301
rect 9021 17245 9107 17301
rect 9163 17245 9249 17301
rect 9305 17245 9391 17301
rect 9447 17245 9533 17301
rect 9589 17245 9675 17301
rect 9731 17245 9817 17301
rect 9873 17245 9959 17301
rect 10015 17245 10101 17301
rect 10157 17245 10243 17301
rect 10299 17245 10385 17301
rect 10441 17245 10527 17301
rect 10583 17245 10669 17301
rect 10725 17245 10811 17301
rect 10867 17245 10953 17301
rect 11009 17245 11095 17301
rect 11151 17245 11237 17301
rect 11293 17245 11379 17301
rect 11435 17245 11521 17301
rect 11577 17245 11663 17301
rect 11719 17245 11805 17301
rect 11861 17245 11947 17301
rect 12003 17245 12089 17301
rect 12145 17245 12231 17301
rect 12287 17245 12373 17301
rect 12429 17245 12515 17301
rect 12571 17245 12657 17301
rect 12713 17245 12799 17301
rect 12855 17245 12941 17301
rect 12997 17245 13083 17301
rect 13139 17245 13225 17301
rect 13281 17245 13367 17301
rect 13423 17245 13509 17301
rect 13565 17245 13651 17301
rect 13707 17245 13793 17301
rect 13849 17245 13935 17301
rect 13991 17245 14077 17301
rect 14133 17245 14219 17301
rect 14275 17245 14361 17301
rect 14417 17245 14503 17301
rect 14559 17245 14645 17301
rect 14701 17245 14787 17301
rect 14843 17245 15000 17301
rect 0 17200 15000 17245
rect 937 17000 3937 17200
rect 4337 17000 7337 17200
rect 7737 17000 10737 17200
rect 11137 17000 14137 17200
rect 0 16941 15000 17000
rect 0 16885 161 16941
rect 217 16885 303 16941
rect 359 16885 445 16941
rect 501 16885 587 16941
rect 643 16885 729 16941
rect 785 16885 871 16941
rect 927 16885 1013 16941
rect 1069 16885 1155 16941
rect 1211 16885 1297 16941
rect 1353 16885 1439 16941
rect 1495 16885 1581 16941
rect 1637 16885 1723 16941
rect 1779 16885 1865 16941
rect 1921 16885 2007 16941
rect 2063 16885 2149 16941
rect 2205 16885 2291 16941
rect 2347 16885 2433 16941
rect 2489 16885 2575 16941
rect 2631 16885 2717 16941
rect 2773 16885 2859 16941
rect 2915 16885 3001 16941
rect 3057 16885 3143 16941
rect 3199 16885 3285 16941
rect 3341 16885 3427 16941
rect 3483 16885 3569 16941
rect 3625 16885 3711 16941
rect 3767 16885 3853 16941
rect 3909 16885 3995 16941
rect 4051 16885 4137 16941
rect 4193 16885 4279 16941
rect 4335 16885 4421 16941
rect 4477 16885 4563 16941
rect 4619 16885 4705 16941
rect 4761 16885 4847 16941
rect 4903 16885 4989 16941
rect 5045 16885 5131 16941
rect 5187 16885 5273 16941
rect 5329 16885 5415 16941
rect 5471 16885 5557 16941
rect 5613 16885 5699 16941
rect 5755 16885 5841 16941
rect 5897 16885 5983 16941
rect 6039 16885 6125 16941
rect 6181 16885 6267 16941
rect 6323 16885 6409 16941
rect 6465 16885 6551 16941
rect 6607 16885 6693 16941
rect 6749 16885 6835 16941
rect 6891 16885 6977 16941
rect 7033 16885 7119 16941
rect 7175 16885 7261 16941
rect 7317 16885 7403 16941
rect 7459 16885 7545 16941
rect 7601 16885 7687 16941
rect 7743 16885 7829 16941
rect 7885 16885 7971 16941
rect 8027 16885 8113 16941
rect 8169 16885 8255 16941
rect 8311 16885 8397 16941
rect 8453 16885 8539 16941
rect 8595 16885 8681 16941
rect 8737 16885 8823 16941
rect 8879 16885 8965 16941
rect 9021 16885 9107 16941
rect 9163 16885 9249 16941
rect 9305 16885 9391 16941
rect 9447 16885 9533 16941
rect 9589 16885 9675 16941
rect 9731 16885 9817 16941
rect 9873 16885 9959 16941
rect 10015 16885 10101 16941
rect 10157 16885 10243 16941
rect 10299 16885 10385 16941
rect 10441 16885 10527 16941
rect 10583 16885 10669 16941
rect 10725 16885 10811 16941
rect 10867 16885 10953 16941
rect 11009 16885 11095 16941
rect 11151 16885 11237 16941
rect 11293 16885 11379 16941
rect 11435 16885 11521 16941
rect 11577 16885 11663 16941
rect 11719 16885 11805 16941
rect 11861 16885 11947 16941
rect 12003 16885 12089 16941
rect 12145 16885 12231 16941
rect 12287 16885 12373 16941
rect 12429 16885 12515 16941
rect 12571 16885 12657 16941
rect 12713 16885 12799 16941
rect 12855 16885 12941 16941
rect 12997 16885 13083 16941
rect 13139 16885 13225 16941
rect 13281 16885 13367 16941
rect 13423 16885 13509 16941
rect 13565 16885 13651 16941
rect 13707 16885 13793 16941
rect 13849 16885 13935 16941
rect 13991 16885 14077 16941
rect 14133 16885 14219 16941
rect 14275 16885 14361 16941
rect 14417 16885 14503 16941
rect 14559 16885 14645 16941
rect 14701 16885 14787 16941
rect 14843 16885 15000 16941
rect 0 16799 15000 16885
rect 0 16743 161 16799
rect 217 16743 303 16799
rect 359 16743 445 16799
rect 501 16743 587 16799
rect 643 16743 729 16799
rect 785 16743 871 16799
rect 927 16743 1013 16799
rect 1069 16743 1155 16799
rect 1211 16743 1297 16799
rect 1353 16743 1439 16799
rect 1495 16743 1581 16799
rect 1637 16743 1723 16799
rect 1779 16743 1865 16799
rect 1921 16743 2007 16799
rect 2063 16743 2149 16799
rect 2205 16743 2291 16799
rect 2347 16743 2433 16799
rect 2489 16743 2575 16799
rect 2631 16743 2717 16799
rect 2773 16743 2859 16799
rect 2915 16743 3001 16799
rect 3057 16743 3143 16799
rect 3199 16743 3285 16799
rect 3341 16743 3427 16799
rect 3483 16743 3569 16799
rect 3625 16743 3711 16799
rect 3767 16743 3853 16799
rect 3909 16743 3995 16799
rect 4051 16743 4137 16799
rect 4193 16743 4279 16799
rect 4335 16743 4421 16799
rect 4477 16743 4563 16799
rect 4619 16743 4705 16799
rect 4761 16743 4847 16799
rect 4903 16743 4989 16799
rect 5045 16743 5131 16799
rect 5187 16743 5273 16799
rect 5329 16743 5415 16799
rect 5471 16743 5557 16799
rect 5613 16743 5699 16799
rect 5755 16743 5841 16799
rect 5897 16743 5983 16799
rect 6039 16743 6125 16799
rect 6181 16743 6267 16799
rect 6323 16743 6409 16799
rect 6465 16743 6551 16799
rect 6607 16743 6693 16799
rect 6749 16743 6835 16799
rect 6891 16743 6977 16799
rect 7033 16743 7119 16799
rect 7175 16743 7261 16799
rect 7317 16743 7403 16799
rect 7459 16743 7545 16799
rect 7601 16743 7687 16799
rect 7743 16743 7829 16799
rect 7885 16743 7971 16799
rect 8027 16743 8113 16799
rect 8169 16743 8255 16799
rect 8311 16743 8397 16799
rect 8453 16743 8539 16799
rect 8595 16743 8681 16799
rect 8737 16743 8823 16799
rect 8879 16743 8965 16799
rect 9021 16743 9107 16799
rect 9163 16743 9249 16799
rect 9305 16743 9391 16799
rect 9447 16743 9533 16799
rect 9589 16743 9675 16799
rect 9731 16743 9817 16799
rect 9873 16743 9959 16799
rect 10015 16743 10101 16799
rect 10157 16743 10243 16799
rect 10299 16743 10385 16799
rect 10441 16743 10527 16799
rect 10583 16743 10669 16799
rect 10725 16743 10811 16799
rect 10867 16743 10953 16799
rect 11009 16743 11095 16799
rect 11151 16743 11237 16799
rect 11293 16743 11379 16799
rect 11435 16743 11521 16799
rect 11577 16743 11663 16799
rect 11719 16743 11805 16799
rect 11861 16743 11947 16799
rect 12003 16743 12089 16799
rect 12145 16743 12231 16799
rect 12287 16743 12373 16799
rect 12429 16743 12515 16799
rect 12571 16743 12657 16799
rect 12713 16743 12799 16799
rect 12855 16743 12941 16799
rect 12997 16743 13083 16799
rect 13139 16743 13225 16799
rect 13281 16743 13367 16799
rect 13423 16743 13509 16799
rect 13565 16743 13651 16799
rect 13707 16743 13793 16799
rect 13849 16743 13935 16799
rect 13991 16743 14077 16799
rect 14133 16743 14219 16799
rect 14275 16743 14361 16799
rect 14417 16743 14503 16799
rect 14559 16743 14645 16799
rect 14701 16743 14787 16799
rect 14843 16743 15000 16799
rect 0 16657 15000 16743
rect 0 16601 161 16657
rect 217 16601 303 16657
rect 359 16601 445 16657
rect 501 16601 587 16657
rect 643 16601 729 16657
rect 785 16601 871 16657
rect 927 16601 1013 16657
rect 1069 16601 1155 16657
rect 1211 16601 1297 16657
rect 1353 16601 1439 16657
rect 1495 16601 1581 16657
rect 1637 16601 1723 16657
rect 1779 16601 1865 16657
rect 1921 16601 2007 16657
rect 2063 16601 2149 16657
rect 2205 16601 2291 16657
rect 2347 16601 2433 16657
rect 2489 16601 2575 16657
rect 2631 16601 2717 16657
rect 2773 16601 2859 16657
rect 2915 16601 3001 16657
rect 3057 16601 3143 16657
rect 3199 16601 3285 16657
rect 3341 16601 3427 16657
rect 3483 16601 3569 16657
rect 3625 16601 3711 16657
rect 3767 16601 3853 16657
rect 3909 16601 3995 16657
rect 4051 16601 4137 16657
rect 4193 16601 4279 16657
rect 4335 16601 4421 16657
rect 4477 16601 4563 16657
rect 4619 16601 4705 16657
rect 4761 16601 4847 16657
rect 4903 16601 4989 16657
rect 5045 16601 5131 16657
rect 5187 16601 5273 16657
rect 5329 16601 5415 16657
rect 5471 16601 5557 16657
rect 5613 16601 5699 16657
rect 5755 16601 5841 16657
rect 5897 16601 5983 16657
rect 6039 16601 6125 16657
rect 6181 16601 6267 16657
rect 6323 16601 6409 16657
rect 6465 16601 6551 16657
rect 6607 16601 6693 16657
rect 6749 16601 6835 16657
rect 6891 16601 6977 16657
rect 7033 16601 7119 16657
rect 7175 16601 7261 16657
rect 7317 16601 7403 16657
rect 7459 16601 7545 16657
rect 7601 16601 7687 16657
rect 7743 16601 7829 16657
rect 7885 16601 7971 16657
rect 8027 16601 8113 16657
rect 8169 16601 8255 16657
rect 8311 16601 8397 16657
rect 8453 16601 8539 16657
rect 8595 16601 8681 16657
rect 8737 16601 8823 16657
rect 8879 16601 8965 16657
rect 9021 16601 9107 16657
rect 9163 16601 9249 16657
rect 9305 16601 9391 16657
rect 9447 16601 9533 16657
rect 9589 16601 9675 16657
rect 9731 16601 9817 16657
rect 9873 16601 9959 16657
rect 10015 16601 10101 16657
rect 10157 16601 10243 16657
rect 10299 16601 10385 16657
rect 10441 16601 10527 16657
rect 10583 16601 10669 16657
rect 10725 16601 10811 16657
rect 10867 16601 10953 16657
rect 11009 16601 11095 16657
rect 11151 16601 11237 16657
rect 11293 16601 11379 16657
rect 11435 16601 11521 16657
rect 11577 16601 11663 16657
rect 11719 16601 11805 16657
rect 11861 16601 11947 16657
rect 12003 16601 12089 16657
rect 12145 16601 12231 16657
rect 12287 16601 12373 16657
rect 12429 16601 12515 16657
rect 12571 16601 12657 16657
rect 12713 16601 12799 16657
rect 12855 16601 12941 16657
rect 12997 16601 13083 16657
rect 13139 16601 13225 16657
rect 13281 16601 13367 16657
rect 13423 16601 13509 16657
rect 13565 16601 13651 16657
rect 13707 16601 13793 16657
rect 13849 16601 13935 16657
rect 13991 16601 14077 16657
rect 14133 16601 14219 16657
rect 14275 16601 14361 16657
rect 14417 16601 14503 16657
rect 14559 16601 14645 16657
rect 14701 16601 14787 16657
rect 14843 16601 15000 16657
rect 0 16515 15000 16601
rect 0 16459 161 16515
rect 217 16459 303 16515
rect 359 16459 445 16515
rect 501 16459 587 16515
rect 643 16459 729 16515
rect 785 16459 871 16515
rect 927 16459 1013 16515
rect 1069 16459 1155 16515
rect 1211 16459 1297 16515
rect 1353 16459 1439 16515
rect 1495 16459 1581 16515
rect 1637 16459 1723 16515
rect 1779 16459 1865 16515
rect 1921 16459 2007 16515
rect 2063 16459 2149 16515
rect 2205 16459 2291 16515
rect 2347 16459 2433 16515
rect 2489 16459 2575 16515
rect 2631 16459 2717 16515
rect 2773 16459 2859 16515
rect 2915 16459 3001 16515
rect 3057 16459 3143 16515
rect 3199 16459 3285 16515
rect 3341 16459 3427 16515
rect 3483 16459 3569 16515
rect 3625 16459 3711 16515
rect 3767 16459 3853 16515
rect 3909 16459 3995 16515
rect 4051 16459 4137 16515
rect 4193 16459 4279 16515
rect 4335 16459 4421 16515
rect 4477 16459 4563 16515
rect 4619 16459 4705 16515
rect 4761 16459 4847 16515
rect 4903 16459 4989 16515
rect 5045 16459 5131 16515
rect 5187 16459 5273 16515
rect 5329 16459 5415 16515
rect 5471 16459 5557 16515
rect 5613 16459 5699 16515
rect 5755 16459 5841 16515
rect 5897 16459 5983 16515
rect 6039 16459 6125 16515
rect 6181 16459 6267 16515
rect 6323 16459 6409 16515
rect 6465 16459 6551 16515
rect 6607 16459 6693 16515
rect 6749 16459 6835 16515
rect 6891 16459 6977 16515
rect 7033 16459 7119 16515
rect 7175 16459 7261 16515
rect 7317 16459 7403 16515
rect 7459 16459 7545 16515
rect 7601 16459 7687 16515
rect 7743 16459 7829 16515
rect 7885 16459 7971 16515
rect 8027 16459 8113 16515
rect 8169 16459 8255 16515
rect 8311 16459 8397 16515
rect 8453 16459 8539 16515
rect 8595 16459 8681 16515
rect 8737 16459 8823 16515
rect 8879 16459 8965 16515
rect 9021 16459 9107 16515
rect 9163 16459 9249 16515
rect 9305 16459 9391 16515
rect 9447 16459 9533 16515
rect 9589 16459 9675 16515
rect 9731 16459 9817 16515
rect 9873 16459 9959 16515
rect 10015 16459 10101 16515
rect 10157 16459 10243 16515
rect 10299 16459 10385 16515
rect 10441 16459 10527 16515
rect 10583 16459 10669 16515
rect 10725 16459 10811 16515
rect 10867 16459 10953 16515
rect 11009 16459 11095 16515
rect 11151 16459 11237 16515
rect 11293 16459 11379 16515
rect 11435 16459 11521 16515
rect 11577 16459 11663 16515
rect 11719 16459 11805 16515
rect 11861 16459 11947 16515
rect 12003 16459 12089 16515
rect 12145 16459 12231 16515
rect 12287 16459 12373 16515
rect 12429 16459 12515 16515
rect 12571 16459 12657 16515
rect 12713 16459 12799 16515
rect 12855 16459 12941 16515
rect 12997 16459 13083 16515
rect 13139 16459 13225 16515
rect 13281 16459 13367 16515
rect 13423 16459 13509 16515
rect 13565 16459 13651 16515
rect 13707 16459 13793 16515
rect 13849 16459 13935 16515
rect 13991 16459 14077 16515
rect 14133 16459 14219 16515
rect 14275 16459 14361 16515
rect 14417 16459 14503 16515
rect 14559 16459 14645 16515
rect 14701 16459 14787 16515
rect 14843 16459 15000 16515
rect 0 16373 15000 16459
rect 0 16317 161 16373
rect 217 16317 303 16373
rect 359 16317 445 16373
rect 501 16317 587 16373
rect 643 16317 729 16373
rect 785 16317 871 16373
rect 927 16317 1013 16373
rect 1069 16317 1155 16373
rect 1211 16317 1297 16373
rect 1353 16317 1439 16373
rect 1495 16317 1581 16373
rect 1637 16317 1723 16373
rect 1779 16317 1865 16373
rect 1921 16317 2007 16373
rect 2063 16317 2149 16373
rect 2205 16317 2291 16373
rect 2347 16317 2433 16373
rect 2489 16317 2575 16373
rect 2631 16317 2717 16373
rect 2773 16317 2859 16373
rect 2915 16317 3001 16373
rect 3057 16317 3143 16373
rect 3199 16317 3285 16373
rect 3341 16317 3427 16373
rect 3483 16317 3569 16373
rect 3625 16317 3711 16373
rect 3767 16317 3853 16373
rect 3909 16317 3995 16373
rect 4051 16317 4137 16373
rect 4193 16317 4279 16373
rect 4335 16317 4421 16373
rect 4477 16317 4563 16373
rect 4619 16317 4705 16373
rect 4761 16317 4847 16373
rect 4903 16317 4989 16373
rect 5045 16317 5131 16373
rect 5187 16317 5273 16373
rect 5329 16317 5415 16373
rect 5471 16317 5557 16373
rect 5613 16317 5699 16373
rect 5755 16317 5841 16373
rect 5897 16317 5983 16373
rect 6039 16317 6125 16373
rect 6181 16317 6267 16373
rect 6323 16317 6409 16373
rect 6465 16317 6551 16373
rect 6607 16317 6693 16373
rect 6749 16317 6835 16373
rect 6891 16317 6977 16373
rect 7033 16317 7119 16373
rect 7175 16317 7261 16373
rect 7317 16317 7403 16373
rect 7459 16317 7545 16373
rect 7601 16317 7687 16373
rect 7743 16317 7829 16373
rect 7885 16317 7971 16373
rect 8027 16317 8113 16373
rect 8169 16317 8255 16373
rect 8311 16317 8397 16373
rect 8453 16317 8539 16373
rect 8595 16317 8681 16373
rect 8737 16317 8823 16373
rect 8879 16317 8965 16373
rect 9021 16317 9107 16373
rect 9163 16317 9249 16373
rect 9305 16317 9391 16373
rect 9447 16317 9533 16373
rect 9589 16317 9675 16373
rect 9731 16317 9817 16373
rect 9873 16317 9959 16373
rect 10015 16317 10101 16373
rect 10157 16317 10243 16373
rect 10299 16317 10385 16373
rect 10441 16317 10527 16373
rect 10583 16317 10669 16373
rect 10725 16317 10811 16373
rect 10867 16317 10953 16373
rect 11009 16317 11095 16373
rect 11151 16317 11237 16373
rect 11293 16317 11379 16373
rect 11435 16317 11521 16373
rect 11577 16317 11663 16373
rect 11719 16317 11805 16373
rect 11861 16317 11947 16373
rect 12003 16317 12089 16373
rect 12145 16317 12231 16373
rect 12287 16317 12373 16373
rect 12429 16317 12515 16373
rect 12571 16317 12657 16373
rect 12713 16317 12799 16373
rect 12855 16317 12941 16373
rect 12997 16317 13083 16373
rect 13139 16317 13225 16373
rect 13281 16317 13367 16373
rect 13423 16317 13509 16373
rect 13565 16317 13651 16373
rect 13707 16317 13793 16373
rect 13849 16317 13935 16373
rect 13991 16317 14077 16373
rect 14133 16317 14219 16373
rect 14275 16317 14361 16373
rect 14417 16317 14503 16373
rect 14559 16317 14645 16373
rect 14701 16317 14787 16373
rect 14843 16317 15000 16373
rect 0 16231 15000 16317
rect 0 16175 161 16231
rect 217 16175 303 16231
rect 359 16175 445 16231
rect 501 16175 587 16231
rect 643 16175 729 16231
rect 785 16175 871 16231
rect 927 16175 1013 16231
rect 1069 16175 1155 16231
rect 1211 16175 1297 16231
rect 1353 16175 1439 16231
rect 1495 16175 1581 16231
rect 1637 16175 1723 16231
rect 1779 16175 1865 16231
rect 1921 16175 2007 16231
rect 2063 16175 2149 16231
rect 2205 16175 2291 16231
rect 2347 16175 2433 16231
rect 2489 16175 2575 16231
rect 2631 16175 2717 16231
rect 2773 16175 2859 16231
rect 2915 16175 3001 16231
rect 3057 16175 3143 16231
rect 3199 16175 3285 16231
rect 3341 16175 3427 16231
rect 3483 16175 3569 16231
rect 3625 16175 3711 16231
rect 3767 16175 3853 16231
rect 3909 16175 3995 16231
rect 4051 16175 4137 16231
rect 4193 16175 4279 16231
rect 4335 16175 4421 16231
rect 4477 16175 4563 16231
rect 4619 16175 4705 16231
rect 4761 16175 4847 16231
rect 4903 16175 4989 16231
rect 5045 16175 5131 16231
rect 5187 16175 5273 16231
rect 5329 16175 5415 16231
rect 5471 16175 5557 16231
rect 5613 16175 5699 16231
rect 5755 16175 5841 16231
rect 5897 16175 5983 16231
rect 6039 16175 6125 16231
rect 6181 16175 6267 16231
rect 6323 16175 6409 16231
rect 6465 16175 6551 16231
rect 6607 16175 6693 16231
rect 6749 16175 6835 16231
rect 6891 16175 6977 16231
rect 7033 16175 7119 16231
rect 7175 16175 7261 16231
rect 7317 16175 7403 16231
rect 7459 16175 7545 16231
rect 7601 16175 7687 16231
rect 7743 16175 7829 16231
rect 7885 16175 7971 16231
rect 8027 16175 8113 16231
rect 8169 16175 8255 16231
rect 8311 16175 8397 16231
rect 8453 16175 8539 16231
rect 8595 16175 8681 16231
rect 8737 16175 8823 16231
rect 8879 16175 8965 16231
rect 9021 16175 9107 16231
rect 9163 16175 9249 16231
rect 9305 16175 9391 16231
rect 9447 16175 9533 16231
rect 9589 16175 9675 16231
rect 9731 16175 9817 16231
rect 9873 16175 9959 16231
rect 10015 16175 10101 16231
rect 10157 16175 10243 16231
rect 10299 16175 10385 16231
rect 10441 16175 10527 16231
rect 10583 16175 10669 16231
rect 10725 16175 10811 16231
rect 10867 16175 10953 16231
rect 11009 16175 11095 16231
rect 11151 16175 11237 16231
rect 11293 16175 11379 16231
rect 11435 16175 11521 16231
rect 11577 16175 11663 16231
rect 11719 16175 11805 16231
rect 11861 16175 11947 16231
rect 12003 16175 12089 16231
rect 12145 16175 12231 16231
rect 12287 16175 12373 16231
rect 12429 16175 12515 16231
rect 12571 16175 12657 16231
rect 12713 16175 12799 16231
rect 12855 16175 12941 16231
rect 12997 16175 13083 16231
rect 13139 16175 13225 16231
rect 13281 16175 13367 16231
rect 13423 16175 13509 16231
rect 13565 16175 13651 16231
rect 13707 16175 13793 16231
rect 13849 16175 13935 16231
rect 13991 16175 14077 16231
rect 14133 16175 14219 16231
rect 14275 16175 14361 16231
rect 14417 16175 14503 16231
rect 14559 16175 14645 16231
rect 14701 16175 14787 16231
rect 14843 16175 15000 16231
rect 0 16089 15000 16175
rect 0 16033 161 16089
rect 217 16033 303 16089
rect 359 16033 445 16089
rect 501 16033 587 16089
rect 643 16033 729 16089
rect 785 16033 871 16089
rect 927 16033 1013 16089
rect 1069 16033 1155 16089
rect 1211 16033 1297 16089
rect 1353 16033 1439 16089
rect 1495 16033 1581 16089
rect 1637 16033 1723 16089
rect 1779 16033 1865 16089
rect 1921 16033 2007 16089
rect 2063 16033 2149 16089
rect 2205 16033 2291 16089
rect 2347 16033 2433 16089
rect 2489 16033 2575 16089
rect 2631 16033 2717 16089
rect 2773 16033 2859 16089
rect 2915 16033 3001 16089
rect 3057 16033 3143 16089
rect 3199 16033 3285 16089
rect 3341 16033 3427 16089
rect 3483 16033 3569 16089
rect 3625 16033 3711 16089
rect 3767 16033 3853 16089
rect 3909 16033 3995 16089
rect 4051 16033 4137 16089
rect 4193 16033 4279 16089
rect 4335 16033 4421 16089
rect 4477 16033 4563 16089
rect 4619 16033 4705 16089
rect 4761 16033 4847 16089
rect 4903 16033 4989 16089
rect 5045 16033 5131 16089
rect 5187 16033 5273 16089
rect 5329 16033 5415 16089
rect 5471 16033 5557 16089
rect 5613 16033 5699 16089
rect 5755 16033 5841 16089
rect 5897 16033 5983 16089
rect 6039 16033 6125 16089
rect 6181 16033 6267 16089
rect 6323 16033 6409 16089
rect 6465 16033 6551 16089
rect 6607 16033 6693 16089
rect 6749 16033 6835 16089
rect 6891 16033 6977 16089
rect 7033 16033 7119 16089
rect 7175 16033 7261 16089
rect 7317 16033 7403 16089
rect 7459 16033 7545 16089
rect 7601 16033 7687 16089
rect 7743 16033 7829 16089
rect 7885 16033 7971 16089
rect 8027 16033 8113 16089
rect 8169 16033 8255 16089
rect 8311 16033 8397 16089
rect 8453 16033 8539 16089
rect 8595 16033 8681 16089
rect 8737 16033 8823 16089
rect 8879 16033 8965 16089
rect 9021 16033 9107 16089
rect 9163 16033 9249 16089
rect 9305 16033 9391 16089
rect 9447 16033 9533 16089
rect 9589 16033 9675 16089
rect 9731 16033 9817 16089
rect 9873 16033 9959 16089
rect 10015 16033 10101 16089
rect 10157 16033 10243 16089
rect 10299 16033 10385 16089
rect 10441 16033 10527 16089
rect 10583 16033 10669 16089
rect 10725 16033 10811 16089
rect 10867 16033 10953 16089
rect 11009 16033 11095 16089
rect 11151 16033 11237 16089
rect 11293 16033 11379 16089
rect 11435 16033 11521 16089
rect 11577 16033 11663 16089
rect 11719 16033 11805 16089
rect 11861 16033 11947 16089
rect 12003 16033 12089 16089
rect 12145 16033 12231 16089
rect 12287 16033 12373 16089
rect 12429 16033 12515 16089
rect 12571 16033 12657 16089
rect 12713 16033 12799 16089
rect 12855 16033 12941 16089
rect 12997 16033 13083 16089
rect 13139 16033 13225 16089
rect 13281 16033 13367 16089
rect 13423 16033 13509 16089
rect 13565 16033 13651 16089
rect 13707 16033 13793 16089
rect 13849 16033 13935 16089
rect 13991 16033 14077 16089
rect 14133 16033 14219 16089
rect 14275 16033 14361 16089
rect 14417 16033 14503 16089
rect 14559 16033 14645 16089
rect 14701 16033 14787 16089
rect 14843 16033 15000 16089
rect 0 15947 15000 16033
rect 0 15891 161 15947
rect 217 15891 303 15947
rect 359 15891 445 15947
rect 501 15891 587 15947
rect 643 15891 729 15947
rect 785 15891 871 15947
rect 927 15891 1013 15947
rect 1069 15891 1155 15947
rect 1211 15891 1297 15947
rect 1353 15891 1439 15947
rect 1495 15891 1581 15947
rect 1637 15891 1723 15947
rect 1779 15891 1865 15947
rect 1921 15891 2007 15947
rect 2063 15891 2149 15947
rect 2205 15891 2291 15947
rect 2347 15891 2433 15947
rect 2489 15891 2575 15947
rect 2631 15891 2717 15947
rect 2773 15891 2859 15947
rect 2915 15891 3001 15947
rect 3057 15891 3143 15947
rect 3199 15891 3285 15947
rect 3341 15891 3427 15947
rect 3483 15891 3569 15947
rect 3625 15891 3711 15947
rect 3767 15891 3853 15947
rect 3909 15891 3995 15947
rect 4051 15891 4137 15947
rect 4193 15891 4279 15947
rect 4335 15891 4421 15947
rect 4477 15891 4563 15947
rect 4619 15891 4705 15947
rect 4761 15891 4847 15947
rect 4903 15891 4989 15947
rect 5045 15891 5131 15947
rect 5187 15891 5273 15947
rect 5329 15891 5415 15947
rect 5471 15891 5557 15947
rect 5613 15891 5699 15947
rect 5755 15891 5841 15947
rect 5897 15891 5983 15947
rect 6039 15891 6125 15947
rect 6181 15891 6267 15947
rect 6323 15891 6409 15947
rect 6465 15891 6551 15947
rect 6607 15891 6693 15947
rect 6749 15891 6835 15947
rect 6891 15891 6977 15947
rect 7033 15891 7119 15947
rect 7175 15891 7261 15947
rect 7317 15891 7403 15947
rect 7459 15891 7545 15947
rect 7601 15891 7687 15947
rect 7743 15891 7829 15947
rect 7885 15891 7971 15947
rect 8027 15891 8113 15947
rect 8169 15891 8255 15947
rect 8311 15891 8397 15947
rect 8453 15891 8539 15947
rect 8595 15891 8681 15947
rect 8737 15891 8823 15947
rect 8879 15891 8965 15947
rect 9021 15891 9107 15947
rect 9163 15891 9249 15947
rect 9305 15891 9391 15947
rect 9447 15891 9533 15947
rect 9589 15891 9675 15947
rect 9731 15891 9817 15947
rect 9873 15891 9959 15947
rect 10015 15891 10101 15947
rect 10157 15891 10243 15947
rect 10299 15891 10385 15947
rect 10441 15891 10527 15947
rect 10583 15891 10669 15947
rect 10725 15891 10811 15947
rect 10867 15891 10953 15947
rect 11009 15891 11095 15947
rect 11151 15891 11237 15947
rect 11293 15891 11379 15947
rect 11435 15891 11521 15947
rect 11577 15891 11663 15947
rect 11719 15891 11805 15947
rect 11861 15891 11947 15947
rect 12003 15891 12089 15947
rect 12145 15891 12231 15947
rect 12287 15891 12373 15947
rect 12429 15891 12515 15947
rect 12571 15891 12657 15947
rect 12713 15891 12799 15947
rect 12855 15891 12941 15947
rect 12997 15891 13083 15947
rect 13139 15891 13225 15947
rect 13281 15891 13367 15947
rect 13423 15891 13509 15947
rect 13565 15891 13651 15947
rect 13707 15891 13793 15947
rect 13849 15891 13935 15947
rect 13991 15891 14077 15947
rect 14133 15891 14219 15947
rect 14275 15891 14361 15947
rect 14417 15891 14503 15947
rect 14559 15891 14645 15947
rect 14701 15891 14787 15947
rect 14843 15891 15000 15947
rect 0 15805 15000 15891
rect 0 15749 161 15805
rect 217 15749 303 15805
rect 359 15749 445 15805
rect 501 15749 587 15805
rect 643 15749 729 15805
rect 785 15749 871 15805
rect 927 15749 1013 15805
rect 1069 15749 1155 15805
rect 1211 15749 1297 15805
rect 1353 15749 1439 15805
rect 1495 15749 1581 15805
rect 1637 15749 1723 15805
rect 1779 15749 1865 15805
rect 1921 15749 2007 15805
rect 2063 15749 2149 15805
rect 2205 15749 2291 15805
rect 2347 15749 2433 15805
rect 2489 15749 2575 15805
rect 2631 15749 2717 15805
rect 2773 15749 2859 15805
rect 2915 15749 3001 15805
rect 3057 15749 3143 15805
rect 3199 15749 3285 15805
rect 3341 15749 3427 15805
rect 3483 15749 3569 15805
rect 3625 15749 3711 15805
rect 3767 15749 3853 15805
rect 3909 15749 3995 15805
rect 4051 15749 4137 15805
rect 4193 15749 4279 15805
rect 4335 15749 4421 15805
rect 4477 15749 4563 15805
rect 4619 15749 4705 15805
rect 4761 15749 4847 15805
rect 4903 15749 4989 15805
rect 5045 15749 5131 15805
rect 5187 15749 5273 15805
rect 5329 15749 5415 15805
rect 5471 15749 5557 15805
rect 5613 15749 5699 15805
rect 5755 15749 5841 15805
rect 5897 15749 5983 15805
rect 6039 15749 6125 15805
rect 6181 15749 6267 15805
rect 6323 15749 6409 15805
rect 6465 15749 6551 15805
rect 6607 15749 6693 15805
rect 6749 15749 6835 15805
rect 6891 15749 6977 15805
rect 7033 15749 7119 15805
rect 7175 15749 7261 15805
rect 7317 15749 7403 15805
rect 7459 15749 7545 15805
rect 7601 15749 7687 15805
rect 7743 15749 7829 15805
rect 7885 15749 7971 15805
rect 8027 15749 8113 15805
rect 8169 15749 8255 15805
rect 8311 15749 8397 15805
rect 8453 15749 8539 15805
rect 8595 15749 8681 15805
rect 8737 15749 8823 15805
rect 8879 15749 8965 15805
rect 9021 15749 9107 15805
rect 9163 15749 9249 15805
rect 9305 15749 9391 15805
rect 9447 15749 9533 15805
rect 9589 15749 9675 15805
rect 9731 15749 9817 15805
rect 9873 15749 9959 15805
rect 10015 15749 10101 15805
rect 10157 15749 10243 15805
rect 10299 15749 10385 15805
rect 10441 15749 10527 15805
rect 10583 15749 10669 15805
rect 10725 15749 10811 15805
rect 10867 15749 10953 15805
rect 11009 15749 11095 15805
rect 11151 15749 11237 15805
rect 11293 15749 11379 15805
rect 11435 15749 11521 15805
rect 11577 15749 11663 15805
rect 11719 15749 11805 15805
rect 11861 15749 11947 15805
rect 12003 15749 12089 15805
rect 12145 15749 12231 15805
rect 12287 15749 12373 15805
rect 12429 15749 12515 15805
rect 12571 15749 12657 15805
rect 12713 15749 12799 15805
rect 12855 15749 12941 15805
rect 12997 15749 13083 15805
rect 13139 15749 13225 15805
rect 13281 15749 13367 15805
rect 13423 15749 13509 15805
rect 13565 15749 13651 15805
rect 13707 15749 13793 15805
rect 13849 15749 13935 15805
rect 13991 15749 14077 15805
rect 14133 15749 14219 15805
rect 14275 15749 14361 15805
rect 14417 15749 14503 15805
rect 14559 15749 14645 15805
rect 14701 15749 14787 15805
rect 14843 15749 15000 15805
rect 0 15663 15000 15749
rect 0 15607 161 15663
rect 217 15607 303 15663
rect 359 15607 445 15663
rect 501 15607 587 15663
rect 643 15607 729 15663
rect 785 15607 871 15663
rect 927 15607 1013 15663
rect 1069 15607 1155 15663
rect 1211 15607 1297 15663
rect 1353 15607 1439 15663
rect 1495 15607 1581 15663
rect 1637 15607 1723 15663
rect 1779 15607 1865 15663
rect 1921 15607 2007 15663
rect 2063 15607 2149 15663
rect 2205 15607 2291 15663
rect 2347 15607 2433 15663
rect 2489 15607 2575 15663
rect 2631 15607 2717 15663
rect 2773 15607 2859 15663
rect 2915 15607 3001 15663
rect 3057 15607 3143 15663
rect 3199 15607 3285 15663
rect 3341 15607 3427 15663
rect 3483 15607 3569 15663
rect 3625 15607 3711 15663
rect 3767 15607 3853 15663
rect 3909 15607 3995 15663
rect 4051 15607 4137 15663
rect 4193 15607 4279 15663
rect 4335 15607 4421 15663
rect 4477 15607 4563 15663
rect 4619 15607 4705 15663
rect 4761 15607 4847 15663
rect 4903 15607 4989 15663
rect 5045 15607 5131 15663
rect 5187 15607 5273 15663
rect 5329 15607 5415 15663
rect 5471 15607 5557 15663
rect 5613 15607 5699 15663
rect 5755 15607 5841 15663
rect 5897 15607 5983 15663
rect 6039 15607 6125 15663
rect 6181 15607 6267 15663
rect 6323 15607 6409 15663
rect 6465 15607 6551 15663
rect 6607 15607 6693 15663
rect 6749 15607 6835 15663
rect 6891 15607 6977 15663
rect 7033 15607 7119 15663
rect 7175 15607 7261 15663
rect 7317 15607 7403 15663
rect 7459 15607 7545 15663
rect 7601 15607 7687 15663
rect 7743 15607 7829 15663
rect 7885 15607 7971 15663
rect 8027 15607 8113 15663
rect 8169 15607 8255 15663
rect 8311 15607 8397 15663
rect 8453 15607 8539 15663
rect 8595 15607 8681 15663
rect 8737 15607 8823 15663
rect 8879 15607 8965 15663
rect 9021 15607 9107 15663
rect 9163 15607 9249 15663
rect 9305 15607 9391 15663
rect 9447 15607 9533 15663
rect 9589 15607 9675 15663
rect 9731 15607 9817 15663
rect 9873 15607 9959 15663
rect 10015 15607 10101 15663
rect 10157 15607 10243 15663
rect 10299 15607 10385 15663
rect 10441 15607 10527 15663
rect 10583 15607 10669 15663
rect 10725 15607 10811 15663
rect 10867 15607 10953 15663
rect 11009 15607 11095 15663
rect 11151 15607 11237 15663
rect 11293 15607 11379 15663
rect 11435 15607 11521 15663
rect 11577 15607 11663 15663
rect 11719 15607 11805 15663
rect 11861 15607 11947 15663
rect 12003 15607 12089 15663
rect 12145 15607 12231 15663
rect 12287 15607 12373 15663
rect 12429 15607 12515 15663
rect 12571 15607 12657 15663
rect 12713 15607 12799 15663
rect 12855 15607 12941 15663
rect 12997 15607 13083 15663
rect 13139 15607 13225 15663
rect 13281 15607 13367 15663
rect 13423 15607 13509 15663
rect 13565 15607 13651 15663
rect 13707 15607 13793 15663
rect 13849 15607 13935 15663
rect 13991 15607 14077 15663
rect 14133 15607 14219 15663
rect 14275 15607 14361 15663
rect 14417 15607 14503 15663
rect 14559 15607 14645 15663
rect 14701 15607 14787 15663
rect 14843 15607 15000 15663
rect 0 15521 15000 15607
rect 0 15465 161 15521
rect 217 15465 303 15521
rect 359 15465 445 15521
rect 501 15465 587 15521
rect 643 15465 729 15521
rect 785 15465 871 15521
rect 927 15465 1013 15521
rect 1069 15465 1155 15521
rect 1211 15465 1297 15521
rect 1353 15465 1439 15521
rect 1495 15465 1581 15521
rect 1637 15465 1723 15521
rect 1779 15465 1865 15521
rect 1921 15465 2007 15521
rect 2063 15465 2149 15521
rect 2205 15465 2291 15521
rect 2347 15465 2433 15521
rect 2489 15465 2575 15521
rect 2631 15465 2717 15521
rect 2773 15465 2859 15521
rect 2915 15465 3001 15521
rect 3057 15465 3143 15521
rect 3199 15465 3285 15521
rect 3341 15465 3427 15521
rect 3483 15465 3569 15521
rect 3625 15465 3711 15521
rect 3767 15465 3853 15521
rect 3909 15465 3995 15521
rect 4051 15465 4137 15521
rect 4193 15465 4279 15521
rect 4335 15465 4421 15521
rect 4477 15465 4563 15521
rect 4619 15465 4705 15521
rect 4761 15465 4847 15521
rect 4903 15465 4989 15521
rect 5045 15465 5131 15521
rect 5187 15465 5273 15521
rect 5329 15465 5415 15521
rect 5471 15465 5557 15521
rect 5613 15465 5699 15521
rect 5755 15465 5841 15521
rect 5897 15465 5983 15521
rect 6039 15465 6125 15521
rect 6181 15465 6267 15521
rect 6323 15465 6409 15521
rect 6465 15465 6551 15521
rect 6607 15465 6693 15521
rect 6749 15465 6835 15521
rect 6891 15465 6977 15521
rect 7033 15465 7119 15521
rect 7175 15465 7261 15521
rect 7317 15465 7403 15521
rect 7459 15465 7545 15521
rect 7601 15465 7687 15521
rect 7743 15465 7829 15521
rect 7885 15465 7971 15521
rect 8027 15465 8113 15521
rect 8169 15465 8255 15521
rect 8311 15465 8397 15521
rect 8453 15465 8539 15521
rect 8595 15465 8681 15521
rect 8737 15465 8823 15521
rect 8879 15465 8965 15521
rect 9021 15465 9107 15521
rect 9163 15465 9249 15521
rect 9305 15465 9391 15521
rect 9447 15465 9533 15521
rect 9589 15465 9675 15521
rect 9731 15465 9817 15521
rect 9873 15465 9959 15521
rect 10015 15465 10101 15521
rect 10157 15465 10243 15521
rect 10299 15465 10385 15521
rect 10441 15465 10527 15521
rect 10583 15465 10669 15521
rect 10725 15465 10811 15521
rect 10867 15465 10953 15521
rect 11009 15465 11095 15521
rect 11151 15465 11237 15521
rect 11293 15465 11379 15521
rect 11435 15465 11521 15521
rect 11577 15465 11663 15521
rect 11719 15465 11805 15521
rect 11861 15465 11947 15521
rect 12003 15465 12089 15521
rect 12145 15465 12231 15521
rect 12287 15465 12373 15521
rect 12429 15465 12515 15521
rect 12571 15465 12657 15521
rect 12713 15465 12799 15521
rect 12855 15465 12941 15521
rect 12997 15465 13083 15521
rect 13139 15465 13225 15521
rect 13281 15465 13367 15521
rect 13423 15465 13509 15521
rect 13565 15465 13651 15521
rect 13707 15465 13793 15521
rect 13849 15465 13935 15521
rect 13991 15465 14077 15521
rect 14133 15465 14219 15521
rect 14275 15465 14361 15521
rect 14417 15465 14503 15521
rect 14559 15465 14645 15521
rect 14701 15465 14787 15521
rect 14843 15465 15000 15521
rect 0 15379 15000 15465
rect 0 15323 161 15379
rect 217 15323 303 15379
rect 359 15323 445 15379
rect 501 15323 587 15379
rect 643 15323 729 15379
rect 785 15323 871 15379
rect 927 15323 1013 15379
rect 1069 15323 1155 15379
rect 1211 15323 1297 15379
rect 1353 15323 1439 15379
rect 1495 15323 1581 15379
rect 1637 15323 1723 15379
rect 1779 15323 1865 15379
rect 1921 15323 2007 15379
rect 2063 15323 2149 15379
rect 2205 15323 2291 15379
rect 2347 15323 2433 15379
rect 2489 15323 2575 15379
rect 2631 15323 2717 15379
rect 2773 15323 2859 15379
rect 2915 15323 3001 15379
rect 3057 15323 3143 15379
rect 3199 15323 3285 15379
rect 3341 15323 3427 15379
rect 3483 15323 3569 15379
rect 3625 15323 3711 15379
rect 3767 15323 3853 15379
rect 3909 15323 3995 15379
rect 4051 15323 4137 15379
rect 4193 15323 4279 15379
rect 4335 15323 4421 15379
rect 4477 15323 4563 15379
rect 4619 15323 4705 15379
rect 4761 15323 4847 15379
rect 4903 15323 4989 15379
rect 5045 15323 5131 15379
rect 5187 15323 5273 15379
rect 5329 15323 5415 15379
rect 5471 15323 5557 15379
rect 5613 15323 5699 15379
rect 5755 15323 5841 15379
rect 5897 15323 5983 15379
rect 6039 15323 6125 15379
rect 6181 15323 6267 15379
rect 6323 15323 6409 15379
rect 6465 15323 6551 15379
rect 6607 15323 6693 15379
rect 6749 15323 6835 15379
rect 6891 15323 6977 15379
rect 7033 15323 7119 15379
rect 7175 15323 7261 15379
rect 7317 15323 7403 15379
rect 7459 15323 7545 15379
rect 7601 15323 7687 15379
rect 7743 15323 7829 15379
rect 7885 15323 7971 15379
rect 8027 15323 8113 15379
rect 8169 15323 8255 15379
rect 8311 15323 8397 15379
rect 8453 15323 8539 15379
rect 8595 15323 8681 15379
rect 8737 15323 8823 15379
rect 8879 15323 8965 15379
rect 9021 15323 9107 15379
rect 9163 15323 9249 15379
rect 9305 15323 9391 15379
rect 9447 15323 9533 15379
rect 9589 15323 9675 15379
rect 9731 15323 9817 15379
rect 9873 15323 9959 15379
rect 10015 15323 10101 15379
rect 10157 15323 10243 15379
rect 10299 15323 10385 15379
rect 10441 15323 10527 15379
rect 10583 15323 10669 15379
rect 10725 15323 10811 15379
rect 10867 15323 10953 15379
rect 11009 15323 11095 15379
rect 11151 15323 11237 15379
rect 11293 15323 11379 15379
rect 11435 15323 11521 15379
rect 11577 15323 11663 15379
rect 11719 15323 11805 15379
rect 11861 15323 11947 15379
rect 12003 15323 12089 15379
rect 12145 15323 12231 15379
rect 12287 15323 12373 15379
rect 12429 15323 12515 15379
rect 12571 15323 12657 15379
rect 12713 15323 12799 15379
rect 12855 15323 12941 15379
rect 12997 15323 13083 15379
rect 13139 15323 13225 15379
rect 13281 15323 13367 15379
rect 13423 15323 13509 15379
rect 13565 15323 13651 15379
rect 13707 15323 13793 15379
rect 13849 15323 13935 15379
rect 13991 15323 14077 15379
rect 14133 15323 14219 15379
rect 14275 15323 14361 15379
rect 14417 15323 14503 15379
rect 14559 15323 14645 15379
rect 14701 15323 14787 15379
rect 14843 15323 15000 15379
rect 0 15237 15000 15323
rect 0 15181 161 15237
rect 217 15181 303 15237
rect 359 15181 445 15237
rect 501 15181 587 15237
rect 643 15181 729 15237
rect 785 15181 871 15237
rect 927 15181 1013 15237
rect 1069 15181 1155 15237
rect 1211 15181 1297 15237
rect 1353 15181 1439 15237
rect 1495 15181 1581 15237
rect 1637 15181 1723 15237
rect 1779 15181 1865 15237
rect 1921 15181 2007 15237
rect 2063 15181 2149 15237
rect 2205 15181 2291 15237
rect 2347 15181 2433 15237
rect 2489 15181 2575 15237
rect 2631 15181 2717 15237
rect 2773 15181 2859 15237
rect 2915 15181 3001 15237
rect 3057 15181 3143 15237
rect 3199 15181 3285 15237
rect 3341 15181 3427 15237
rect 3483 15181 3569 15237
rect 3625 15181 3711 15237
rect 3767 15181 3853 15237
rect 3909 15181 3995 15237
rect 4051 15181 4137 15237
rect 4193 15181 4279 15237
rect 4335 15181 4421 15237
rect 4477 15181 4563 15237
rect 4619 15181 4705 15237
rect 4761 15181 4847 15237
rect 4903 15181 4989 15237
rect 5045 15181 5131 15237
rect 5187 15181 5273 15237
rect 5329 15181 5415 15237
rect 5471 15181 5557 15237
rect 5613 15181 5699 15237
rect 5755 15181 5841 15237
rect 5897 15181 5983 15237
rect 6039 15181 6125 15237
rect 6181 15181 6267 15237
rect 6323 15181 6409 15237
rect 6465 15181 6551 15237
rect 6607 15181 6693 15237
rect 6749 15181 6835 15237
rect 6891 15181 6977 15237
rect 7033 15181 7119 15237
rect 7175 15181 7261 15237
rect 7317 15181 7403 15237
rect 7459 15181 7545 15237
rect 7601 15181 7687 15237
rect 7743 15181 7829 15237
rect 7885 15181 7971 15237
rect 8027 15181 8113 15237
rect 8169 15181 8255 15237
rect 8311 15181 8397 15237
rect 8453 15181 8539 15237
rect 8595 15181 8681 15237
rect 8737 15181 8823 15237
rect 8879 15181 8965 15237
rect 9021 15181 9107 15237
rect 9163 15181 9249 15237
rect 9305 15181 9391 15237
rect 9447 15181 9533 15237
rect 9589 15181 9675 15237
rect 9731 15181 9817 15237
rect 9873 15181 9959 15237
rect 10015 15181 10101 15237
rect 10157 15181 10243 15237
rect 10299 15181 10385 15237
rect 10441 15181 10527 15237
rect 10583 15181 10669 15237
rect 10725 15181 10811 15237
rect 10867 15181 10953 15237
rect 11009 15181 11095 15237
rect 11151 15181 11237 15237
rect 11293 15181 11379 15237
rect 11435 15181 11521 15237
rect 11577 15181 11663 15237
rect 11719 15181 11805 15237
rect 11861 15181 11947 15237
rect 12003 15181 12089 15237
rect 12145 15181 12231 15237
rect 12287 15181 12373 15237
rect 12429 15181 12515 15237
rect 12571 15181 12657 15237
rect 12713 15181 12799 15237
rect 12855 15181 12941 15237
rect 12997 15181 13083 15237
rect 13139 15181 13225 15237
rect 13281 15181 13367 15237
rect 13423 15181 13509 15237
rect 13565 15181 13651 15237
rect 13707 15181 13793 15237
rect 13849 15181 13935 15237
rect 13991 15181 14077 15237
rect 14133 15181 14219 15237
rect 14275 15181 14361 15237
rect 14417 15181 14503 15237
rect 14559 15181 14645 15237
rect 14701 15181 14787 15237
rect 14843 15181 15000 15237
rect 0 15095 15000 15181
rect 0 15039 161 15095
rect 217 15039 303 15095
rect 359 15039 445 15095
rect 501 15039 587 15095
rect 643 15039 729 15095
rect 785 15039 871 15095
rect 927 15039 1013 15095
rect 1069 15039 1155 15095
rect 1211 15039 1297 15095
rect 1353 15039 1439 15095
rect 1495 15039 1581 15095
rect 1637 15039 1723 15095
rect 1779 15039 1865 15095
rect 1921 15039 2007 15095
rect 2063 15039 2149 15095
rect 2205 15039 2291 15095
rect 2347 15039 2433 15095
rect 2489 15039 2575 15095
rect 2631 15039 2717 15095
rect 2773 15039 2859 15095
rect 2915 15039 3001 15095
rect 3057 15039 3143 15095
rect 3199 15039 3285 15095
rect 3341 15039 3427 15095
rect 3483 15039 3569 15095
rect 3625 15039 3711 15095
rect 3767 15039 3853 15095
rect 3909 15039 3995 15095
rect 4051 15039 4137 15095
rect 4193 15039 4279 15095
rect 4335 15039 4421 15095
rect 4477 15039 4563 15095
rect 4619 15039 4705 15095
rect 4761 15039 4847 15095
rect 4903 15039 4989 15095
rect 5045 15039 5131 15095
rect 5187 15039 5273 15095
rect 5329 15039 5415 15095
rect 5471 15039 5557 15095
rect 5613 15039 5699 15095
rect 5755 15039 5841 15095
rect 5897 15039 5983 15095
rect 6039 15039 6125 15095
rect 6181 15039 6267 15095
rect 6323 15039 6409 15095
rect 6465 15039 6551 15095
rect 6607 15039 6693 15095
rect 6749 15039 6835 15095
rect 6891 15039 6977 15095
rect 7033 15039 7119 15095
rect 7175 15039 7261 15095
rect 7317 15039 7403 15095
rect 7459 15039 7545 15095
rect 7601 15039 7687 15095
rect 7743 15039 7829 15095
rect 7885 15039 7971 15095
rect 8027 15039 8113 15095
rect 8169 15039 8255 15095
rect 8311 15039 8397 15095
rect 8453 15039 8539 15095
rect 8595 15039 8681 15095
rect 8737 15039 8823 15095
rect 8879 15039 8965 15095
rect 9021 15039 9107 15095
rect 9163 15039 9249 15095
rect 9305 15039 9391 15095
rect 9447 15039 9533 15095
rect 9589 15039 9675 15095
rect 9731 15039 9817 15095
rect 9873 15039 9959 15095
rect 10015 15039 10101 15095
rect 10157 15039 10243 15095
rect 10299 15039 10385 15095
rect 10441 15039 10527 15095
rect 10583 15039 10669 15095
rect 10725 15039 10811 15095
rect 10867 15039 10953 15095
rect 11009 15039 11095 15095
rect 11151 15039 11237 15095
rect 11293 15039 11379 15095
rect 11435 15039 11521 15095
rect 11577 15039 11663 15095
rect 11719 15039 11805 15095
rect 11861 15039 11947 15095
rect 12003 15039 12089 15095
rect 12145 15039 12231 15095
rect 12287 15039 12373 15095
rect 12429 15039 12515 15095
rect 12571 15039 12657 15095
rect 12713 15039 12799 15095
rect 12855 15039 12941 15095
rect 12997 15039 13083 15095
rect 13139 15039 13225 15095
rect 13281 15039 13367 15095
rect 13423 15039 13509 15095
rect 13565 15039 13651 15095
rect 13707 15039 13793 15095
rect 13849 15039 13935 15095
rect 13991 15039 14077 15095
rect 14133 15039 14219 15095
rect 14275 15039 14361 15095
rect 14417 15039 14503 15095
rect 14559 15039 14645 15095
rect 14701 15039 14787 15095
rect 14843 15039 15000 15095
rect 0 14953 15000 15039
rect 0 14897 161 14953
rect 217 14897 303 14953
rect 359 14897 445 14953
rect 501 14897 587 14953
rect 643 14897 729 14953
rect 785 14897 871 14953
rect 927 14897 1013 14953
rect 1069 14897 1155 14953
rect 1211 14897 1297 14953
rect 1353 14897 1439 14953
rect 1495 14897 1581 14953
rect 1637 14897 1723 14953
rect 1779 14897 1865 14953
rect 1921 14897 2007 14953
rect 2063 14897 2149 14953
rect 2205 14897 2291 14953
rect 2347 14897 2433 14953
rect 2489 14897 2575 14953
rect 2631 14897 2717 14953
rect 2773 14897 2859 14953
rect 2915 14897 3001 14953
rect 3057 14897 3143 14953
rect 3199 14897 3285 14953
rect 3341 14897 3427 14953
rect 3483 14897 3569 14953
rect 3625 14897 3711 14953
rect 3767 14897 3853 14953
rect 3909 14897 3995 14953
rect 4051 14897 4137 14953
rect 4193 14897 4279 14953
rect 4335 14897 4421 14953
rect 4477 14897 4563 14953
rect 4619 14897 4705 14953
rect 4761 14897 4847 14953
rect 4903 14897 4989 14953
rect 5045 14897 5131 14953
rect 5187 14897 5273 14953
rect 5329 14897 5415 14953
rect 5471 14897 5557 14953
rect 5613 14897 5699 14953
rect 5755 14897 5841 14953
rect 5897 14897 5983 14953
rect 6039 14897 6125 14953
rect 6181 14897 6267 14953
rect 6323 14897 6409 14953
rect 6465 14897 6551 14953
rect 6607 14897 6693 14953
rect 6749 14897 6835 14953
rect 6891 14897 6977 14953
rect 7033 14897 7119 14953
rect 7175 14897 7261 14953
rect 7317 14897 7403 14953
rect 7459 14897 7545 14953
rect 7601 14897 7687 14953
rect 7743 14897 7829 14953
rect 7885 14897 7971 14953
rect 8027 14897 8113 14953
rect 8169 14897 8255 14953
rect 8311 14897 8397 14953
rect 8453 14897 8539 14953
rect 8595 14897 8681 14953
rect 8737 14897 8823 14953
rect 8879 14897 8965 14953
rect 9021 14897 9107 14953
rect 9163 14897 9249 14953
rect 9305 14897 9391 14953
rect 9447 14897 9533 14953
rect 9589 14897 9675 14953
rect 9731 14897 9817 14953
rect 9873 14897 9959 14953
rect 10015 14897 10101 14953
rect 10157 14897 10243 14953
rect 10299 14897 10385 14953
rect 10441 14897 10527 14953
rect 10583 14897 10669 14953
rect 10725 14897 10811 14953
rect 10867 14897 10953 14953
rect 11009 14897 11095 14953
rect 11151 14897 11237 14953
rect 11293 14897 11379 14953
rect 11435 14897 11521 14953
rect 11577 14897 11663 14953
rect 11719 14897 11805 14953
rect 11861 14897 11947 14953
rect 12003 14897 12089 14953
rect 12145 14897 12231 14953
rect 12287 14897 12373 14953
rect 12429 14897 12515 14953
rect 12571 14897 12657 14953
rect 12713 14897 12799 14953
rect 12855 14897 12941 14953
rect 12997 14897 13083 14953
rect 13139 14897 13225 14953
rect 13281 14897 13367 14953
rect 13423 14897 13509 14953
rect 13565 14897 13651 14953
rect 13707 14897 13793 14953
rect 13849 14897 13935 14953
rect 13991 14897 14077 14953
rect 14133 14897 14219 14953
rect 14275 14897 14361 14953
rect 14417 14897 14503 14953
rect 14559 14897 14645 14953
rect 14701 14897 14787 14953
rect 14843 14897 15000 14953
rect 0 14811 15000 14897
rect 0 14755 161 14811
rect 217 14755 303 14811
rect 359 14755 445 14811
rect 501 14755 587 14811
rect 643 14755 729 14811
rect 785 14755 871 14811
rect 927 14755 1013 14811
rect 1069 14755 1155 14811
rect 1211 14755 1297 14811
rect 1353 14755 1439 14811
rect 1495 14755 1581 14811
rect 1637 14755 1723 14811
rect 1779 14755 1865 14811
rect 1921 14755 2007 14811
rect 2063 14755 2149 14811
rect 2205 14755 2291 14811
rect 2347 14755 2433 14811
rect 2489 14755 2575 14811
rect 2631 14755 2717 14811
rect 2773 14755 2859 14811
rect 2915 14755 3001 14811
rect 3057 14755 3143 14811
rect 3199 14755 3285 14811
rect 3341 14755 3427 14811
rect 3483 14755 3569 14811
rect 3625 14755 3711 14811
rect 3767 14755 3853 14811
rect 3909 14755 3995 14811
rect 4051 14755 4137 14811
rect 4193 14755 4279 14811
rect 4335 14755 4421 14811
rect 4477 14755 4563 14811
rect 4619 14755 4705 14811
rect 4761 14755 4847 14811
rect 4903 14755 4989 14811
rect 5045 14755 5131 14811
rect 5187 14755 5273 14811
rect 5329 14755 5415 14811
rect 5471 14755 5557 14811
rect 5613 14755 5699 14811
rect 5755 14755 5841 14811
rect 5897 14755 5983 14811
rect 6039 14755 6125 14811
rect 6181 14755 6267 14811
rect 6323 14755 6409 14811
rect 6465 14755 6551 14811
rect 6607 14755 6693 14811
rect 6749 14755 6835 14811
rect 6891 14755 6977 14811
rect 7033 14755 7119 14811
rect 7175 14755 7261 14811
rect 7317 14755 7403 14811
rect 7459 14755 7545 14811
rect 7601 14755 7687 14811
rect 7743 14755 7829 14811
rect 7885 14755 7971 14811
rect 8027 14755 8113 14811
rect 8169 14755 8255 14811
rect 8311 14755 8397 14811
rect 8453 14755 8539 14811
rect 8595 14755 8681 14811
rect 8737 14755 8823 14811
rect 8879 14755 8965 14811
rect 9021 14755 9107 14811
rect 9163 14755 9249 14811
rect 9305 14755 9391 14811
rect 9447 14755 9533 14811
rect 9589 14755 9675 14811
rect 9731 14755 9817 14811
rect 9873 14755 9959 14811
rect 10015 14755 10101 14811
rect 10157 14755 10243 14811
rect 10299 14755 10385 14811
rect 10441 14755 10527 14811
rect 10583 14755 10669 14811
rect 10725 14755 10811 14811
rect 10867 14755 10953 14811
rect 11009 14755 11095 14811
rect 11151 14755 11237 14811
rect 11293 14755 11379 14811
rect 11435 14755 11521 14811
rect 11577 14755 11663 14811
rect 11719 14755 11805 14811
rect 11861 14755 11947 14811
rect 12003 14755 12089 14811
rect 12145 14755 12231 14811
rect 12287 14755 12373 14811
rect 12429 14755 12515 14811
rect 12571 14755 12657 14811
rect 12713 14755 12799 14811
rect 12855 14755 12941 14811
rect 12997 14755 13083 14811
rect 13139 14755 13225 14811
rect 13281 14755 13367 14811
rect 13423 14755 13509 14811
rect 13565 14755 13651 14811
rect 13707 14755 13793 14811
rect 13849 14755 13935 14811
rect 13991 14755 14077 14811
rect 14133 14755 14219 14811
rect 14275 14755 14361 14811
rect 14417 14755 14503 14811
rect 14559 14755 14645 14811
rect 14701 14755 14787 14811
rect 14843 14755 15000 14811
rect 0 14669 15000 14755
rect 0 14613 161 14669
rect 217 14613 303 14669
rect 359 14613 445 14669
rect 501 14613 587 14669
rect 643 14613 729 14669
rect 785 14613 871 14669
rect 927 14613 1013 14669
rect 1069 14613 1155 14669
rect 1211 14613 1297 14669
rect 1353 14613 1439 14669
rect 1495 14613 1581 14669
rect 1637 14613 1723 14669
rect 1779 14613 1865 14669
rect 1921 14613 2007 14669
rect 2063 14613 2149 14669
rect 2205 14613 2291 14669
rect 2347 14613 2433 14669
rect 2489 14613 2575 14669
rect 2631 14613 2717 14669
rect 2773 14613 2859 14669
rect 2915 14613 3001 14669
rect 3057 14613 3143 14669
rect 3199 14613 3285 14669
rect 3341 14613 3427 14669
rect 3483 14613 3569 14669
rect 3625 14613 3711 14669
rect 3767 14613 3853 14669
rect 3909 14613 3995 14669
rect 4051 14613 4137 14669
rect 4193 14613 4279 14669
rect 4335 14613 4421 14669
rect 4477 14613 4563 14669
rect 4619 14613 4705 14669
rect 4761 14613 4847 14669
rect 4903 14613 4989 14669
rect 5045 14613 5131 14669
rect 5187 14613 5273 14669
rect 5329 14613 5415 14669
rect 5471 14613 5557 14669
rect 5613 14613 5699 14669
rect 5755 14613 5841 14669
rect 5897 14613 5983 14669
rect 6039 14613 6125 14669
rect 6181 14613 6267 14669
rect 6323 14613 6409 14669
rect 6465 14613 6551 14669
rect 6607 14613 6693 14669
rect 6749 14613 6835 14669
rect 6891 14613 6977 14669
rect 7033 14613 7119 14669
rect 7175 14613 7261 14669
rect 7317 14613 7403 14669
rect 7459 14613 7545 14669
rect 7601 14613 7687 14669
rect 7743 14613 7829 14669
rect 7885 14613 7971 14669
rect 8027 14613 8113 14669
rect 8169 14613 8255 14669
rect 8311 14613 8397 14669
rect 8453 14613 8539 14669
rect 8595 14613 8681 14669
rect 8737 14613 8823 14669
rect 8879 14613 8965 14669
rect 9021 14613 9107 14669
rect 9163 14613 9249 14669
rect 9305 14613 9391 14669
rect 9447 14613 9533 14669
rect 9589 14613 9675 14669
rect 9731 14613 9817 14669
rect 9873 14613 9959 14669
rect 10015 14613 10101 14669
rect 10157 14613 10243 14669
rect 10299 14613 10385 14669
rect 10441 14613 10527 14669
rect 10583 14613 10669 14669
rect 10725 14613 10811 14669
rect 10867 14613 10953 14669
rect 11009 14613 11095 14669
rect 11151 14613 11237 14669
rect 11293 14613 11379 14669
rect 11435 14613 11521 14669
rect 11577 14613 11663 14669
rect 11719 14613 11805 14669
rect 11861 14613 11947 14669
rect 12003 14613 12089 14669
rect 12145 14613 12231 14669
rect 12287 14613 12373 14669
rect 12429 14613 12515 14669
rect 12571 14613 12657 14669
rect 12713 14613 12799 14669
rect 12855 14613 12941 14669
rect 12997 14613 13083 14669
rect 13139 14613 13225 14669
rect 13281 14613 13367 14669
rect 13423 14613 13509 14669
rect 13565 14613 13651 14669
rect 13707 14613 13793 14669
rect 13849 14613 13935 14669
rect 13991 14613 14077 14669
rect 14133 14613 14219 14669
rect 14275 14613 14361 14669
rect 14417 14613 14503 14669
rect 14559 14613 14645 14669
rect 14701 14613 14787 14669
rect 14843 14613 15000 14669
rect 0 14527 15000 14613
rect 0 14471 161 14527
rect 217 14471 303 14527
rect 359 14471 445 14527
rect 501 14471 587 14527
rect 643 14471 729 14527
rect 785 14471 871 14527
rect 927 14471 1013 14527
rect 1069 14471 1155 14527
rect 1211 14471 1297 14527
rect 1353 14471 1439 14527
rect 1495 14471 1581 14527
rect 1637 14471 1723 14527
rect 1779 14471 1865 14527
rect 1921 14471 2007 14527
rect 2063 14471 2149 14527
rect 2205 14471 2291 14527
rect 2347 14471 2433 14527
rect 2489 14471 2575 14527
rect 2631 14471 2717 14527
rect 2773 14471 2859 14527
rect 2915 14471 3001 14527
rect 3057 14471 3143 14527
rect 3199 14471 3285 14527
rect 3341 14471 3427 14527
rect 3483 14471 3569 14527
rect 3625 14471 3711 14527
rect 3767 14471 3853 14527
rect 3909 14471 3995 14527
rect 4051 14471 4137 14527
rect 4193 14471 4279 14527
rect 4335 14471 4421 14527
rect 4477 14471 4563 14527
rect 4619 14471 4705 14527
rect 4761 14471 4847 14527
rect 4903 14471 4989 14527
rect 5045 14471 5131 14527
rect 5187 14471 5273 14527
rect 5329 14471 5415 14527
rect 5471 14471 5557 14527
rect 5613 14471 5699 14527
rect 5755 14471 5841 14527
rect 5897 14471 5983 14527
rect 6039 14471 6125 14527
rect 6181 14471 6267 14527
rect 6323 14471 6409 14527
rect 6465 14471 6551 14527
rect 6607 14471 6693 14527
rect 6749 14471 6835 14527
rect 6891 14471 6977 14527
rect 7033 14471 7119 14527
rect 7175 14471 7261 14527
rect 7317 14471 7403 14527
rect 7459 14471 7545 14527
rect 7601 14471 7687 14527
rect 7743 14471 7829 14527
rect 7885 14471 7971 14527
rect 8027 14471 8113 14527
rect 8169 14471 8255 14527
rect 8311 14471 8397 14527
rect 8453 14471 8539 14527
rect 8595 14471 8681 14527
rect 8737 14471 8823 14527
rect 8879 14471 8965 14527
rect 9021 14471 9107 14527
rect 9163 14471 9249 14527
rect 9305 14471 9391 14527
rect 9447 14471 9533 14527
rect 9589 14471 9675 14527
rect 9731 14471 9817 14527
rect 9873 14471 9959 14527
rect 10015 14471 10101 14527
rect 10157 14471 10243 14527
rect 10299 14471 10385 14527
rect 10441 14471 10527 14527
rect 10583 14471 10669 14527
rect 10725 14471 10811 14527
rect 10867 14471 10953 14527
rect 11009 14471 11095 14527
rect 11151 14471 11237 14527
rect 11293 14471 11379 14527
rect 11435 14471 11521 14527
rect 11577 14471 11663 14527
rect 11719 14471 11805 14527
rect 11861 14471 11947 14527
rect 12003 14471 12089 14527
rect 12145 14471 12231 14527
rect 12287 14471 12373 14527
rect 12429 14471 12515 14527
rect 12571 14471 12657 14527
rect 12713 14471 12799 14527
rect 12855 14471 12941 14527
rect 12997 14471 13083 14527
rect 13139 14471 13225 14527
rect 13281 14471 13367 14527
rect 13423 14471 13509 14527
rect 13565 14471 13651 14527
rect 13707 14471 13793 14527
rect 13849 14471 13935 14527
rect 13991 14471 14077 14527
rect 14133 14471 14219 14527
rect 14275 14471 14361 14527
rect 14417 14471 14503 14527
rect 14559 14471 14645 14527
rect 14701 14471 14787 14527
rect 14843 14471 15000 14527
rect 0 14385 15000 14471
rect 0 14329 161 14385
rect 217 14329 303 14385
rect 359 14329 445 14385
rect 501 14329 587 14385
rect 643 14329 729 14385
rect 785 14329 871 14385
rect 927 14329 1013 14385
rect 1069 14329 1155 14385
rect 1211 14329 1297 14385
rect 1353 14329 1439 14385
rect 1495 14329 1581 14385
rect 1637 14329 1723 14385
rect 1779 14329 1865 14385
rect 1921 14329 2007 14385
rect 2063 14329 2149 14385
rect 2205 14329 2291 14385
rect 2347 14329 2433 14385
rect 2489 14329 2575 14385
rect 2631 14329 2717 14385
rect 2773 14329 2859 14385
rect 2915 14329 3001 14385
rect 3057 14329 3143 14385
rect 3199 14329 3285 14385
rect 3341 14329 3427 14385
rect 3483 14329 3569 14385
rect 3625 14329 3711 14385
rect 3767 14329 3853 14385
rect 3909 14329 3995 14385
rect 4051 14329 4137 14385
rect 4193 14329 4279 14385
rect 4335 14329 4421 14385
rect 4477 14329 4563 14385
rect 4619 14329 4705 14385
rect 4761 14329 4847 14385
rect 4903 14329 4989 14385
rect 5045 14329 5131 14385
rect 5187 14329 5273 14385
rect 5329 14329 5415 14385
rect 5471 14329 5557 14385
rect 5613 14329 5699 14385
rect 5755 14329 5841 14385
rect 5897 14329 5983 14385
rect 6039 14329 6125 14385
rect 6181 14329 6267 14385
rect 6323 14329 6409 14385
rect 6465 14329 6551 14385
rect 6607 14329 6693 14385
rect 6749 14329 6835 14385
rect 6891 14329 6977 14385
rect 7033 14329 7119 14385
rect 7175 14329 7261 14385
rect 7317 14329 7403 14385
rect 7459 14329 7545 14385
rect 7601 14329 7687 14385
rect 7743 14329 7829 14385
rect 7885 14329 7971 14385
rect 8027 14329 8113 14385
rect 8169 14329 8255 14385
rect 8311 14329 8397 14385
rect 8453 14329 8539 14385
rect 8595 14329 8681 14385
rect 8737 14329 8823 14385
rect 8879 14329 8965 14385
rect 9021 14329 9107 14385
rect 9163 14329 9249 14385
rect 9305 14329 9391 14385
rect 9447 14329 9533 14385
rect 9589 14329 9675 14385
rect 9731 14329 9817 14385
rect 9873 14329 9959 14385
rect 10015 14329 10101 14385
rect 10157 14329 10243 14385
rect 10299 14329 10385 14385
rect 10441 14329 10527 14385
rect 10583 14329 10669 14385
rect 10725 14329 10811 14385
rect 10867 14329 10953 14385
rect 11009 14329 11095 14385
rect 11151 14329 11237 14385
rect 11293 14329 11379 14385
rect 11435 14329 11521 14385
rect 11577 14329 11663 14385
rect 11719 14329 11805 14385
rect 11861 14329 11947 14385
rect 12003 14329 12089 14385
rect 12145 14329 12231 14385
rect 12287 14329 12373 14385
rect 12429 14329 12515 14385
rect 12571 14329 12657 14385
rect 12713 14329 12799 14385
rect 12855 14329 12941 14385
rect 12997 14329 13083 14385
rect 13139 14329 13225 14385
rect 13281 14329 13367 14385
rect 13423 14329 13509 14385
rect 13565 14329 13651 14385
rect 13707 14329 13793 14385
rect 13849 14329 13935 14385
rect 13991 14329 14077 14385
rect 14133 14329 14219 14385
rect 14275 14329 14361 14385
rect 14417 14329 14503 14385
rect 14559 14329 14645 14385
rect 14701 14329 14787 14385
rect 14843 14329 15000 14385
rect 0 14243 15000 14329
rect 0 14187 161 14243
rect 217 14187 303 14243
rect 359 14187 445 14243
rect 501 14187 587 14243
rect 643 14187 729 14243
rect 785 14187 871 14243
rect 927 14187 1013 14243
rect 1069 14187 1155 14243
rect 1211 14187 1297 14243
rect 1353 14187 1439 14243
rect 1495 14187 1581 14243
rect 1637 14187 1723 14243
rect 1779 14187 1865 14243
rect 1921 14187 2007 14243
rect 2063 14187 2149 14243
rect 2205 14187 2291 14243
rect 2347 14187 2433 14243
rect 2489 14187 2575 14243
rect 2631 14187 2717 14243
rect 2773 14187 2859 14243
rect 2915 14187 3001 14243
rect 3057 14187 3143 14243
rect 3199 14187 3285 14243
rect 3341 14187 3427 14243
rect 3483 14187 3569 14243
rect 3625 14187 3711 14243
rect 3767 14187 3853 14243
rect 3909 14187 3995 14243
rect 4051 14187 4137 14243
rect 4193 14187 4279 14243
rect 4335 14187 4421 14243
rect 4477 14187 4563 14243
rect 4619 14187 4705 14243
rect 4761 14187 4847 14243
rect 4903 14187 4989 14243
rect 5045 14187 5131 14243
rect 5187 14187 5273 14243
rect 5329 14187 5415 14243
rect 5471 14187 5557 14243
rect 5613 14187 5699 14243
rect 5755 14187 5841 14243
rect 5897 14187 5983 14243
rect 6039 14187 6125 14243
rect 6181 14187 6267 14243
rect 6323 14187 6409 14243
rect 6465 14187 6551 14243
rect 6607 14187 6693 14243
rect 6749 14187 6835 14243
rect 6891 14187 6977 14243
rect 7033 14187 7119 14243
rect 7175 14187 7261 14243
rect 7317 14187 7403 14243
rect 7459 14187 7545 14243
rect 7601 14187 7687 14243
rect 7743 14187 7829 14243
rect 7885 14187 7971 14243
rect 8027 14187 8113 14243
rect 8169 14187 8255 14243
rect 8311 14187 8397 14243
rect 8453 14187 8539 14243
rect 8595 14187 8681 14243
rect 8737 14187 8823 14243
rect 8879 14187 8965 14243
rect 9021 14187 9107 14243
rect 9163 14187 9249 14243
rect 9305 14187 9391 14243
rect 9447 14187 9533 14243
rect 9589 14187 9675 14243
rect 9731 14187 9817 14243
rect 9873 14187 9959 14243
rect 10015 14187 10101 14243
rect 10157 14187 10243 14243
rect 10299 14187 10385 14243
rect 10441 14187 10527 14243
rect 10583 14187 10669 14243
rect 10725 14187 10811 14243
rect 10867 14187 10953 14243
rect 11009 14187 11095 14243
rect 11151 14187 11237 14243
rect 11293 14187 11379 14243
rect 11435 14187 11521 14243
rect 11577 14187 11663 14243
rect 11719 14187 11805 14243
rect 11861 14187 11947 14243
rect 12003 14187 12089 14243
rect 12145 14187 12231 14243
rect 12287 14187 12373 14243
rect 12429 14187 12515 14243
rect 12571 14187 12657 14243
rect 12713 14187 12799 14243
rect 12855 14187 12941 14243
rect 12997 14187 13083 14243
rect 13139 14187 13225 14243
rect 13281 14187 13367 14243
rect 13423 14187 13509 14243
rect 13565 14187 13651 14243
rect 13707 14187 13793 14243
rect 13849 14187 13935 14243
rect 13991 14187 14077 14243
rect 14133 14187 14219 14243
rect 14275 14187 14361 14243
rect 14417 14187 14503 14243
rect 14559 14187 14645 14243
rect 14701 14187 14787 14243
rect 14843 14187 15000 14243
rect 0 14101 15000 14187
rect 0 14045 161 14101
rect 217 14045 303 14101
rect 359 14045 445 14101
rect 501 14045 587 14101
rect 643 14045 729 14101
rect 785 14045 871 14101
rect 927 14045 1013 14101
rect 1069 14045 1155 14101
rect 1211 14045 1297 14101
rect 1353 14045 1439 14101
rect 1495 14045 1581 14101
rect 1637 14045 1723 14101
rect 1779 14045 1865 14101
rect 1921 14045 2007 14101
rect 2063 14045 2149 14101
rect 2205 14045 2291 14101
rect 2347 14045 2433 14101
rect 2489 14045 2575 14101
rect 2631 14045 2717 14101
rect 2773 14045 2859 14101
rect 2915 14045 3001 14101
rect 3057 14045 3143 14101
rect 3199 14045 3285 14101
rect 3341 14045 3427 14101
rect 3483 14045 3569 14101
rect 3625 14045 3711 14101
rect 3767 14045 3853 14101
rect 3909 14045 3995 14101
rect 4051 14045 4137 14101
rect 4193 14045 4279 14101
rect 4335 14045 4421 14101
rect 4477 14045 4563 14101
rect 4619 14045 4705 14101
rect 4761 14045 4847 14101
rect 4903 14045 4989 14101
rect 5045 14045 5131 14101
rect 5187 14045 5273 14101
rect 5329 14045 5415 14101
rect 5471 14045 5557 14101
rect 5613 14045 5699 14101
rect 5755 14045 5841 14101
rect 5897 14045 5983 14101
rect 6039 14045 6125 14101
rect 6181 14045 6267 14101
rect 6323 14045 6409 14101
rect 6465 14045 6551 14101
rect 6607 14045 6693 14101
rect 6749 14045 6835 14101
rect 6891 14045 6977 14101
rect 7033 14045 7119 14101
rect 7175 14045 7261 14101
rect 7317 14045 7403 14101
rect 7459 14045 7545 14101
rect 7601 14045 7687 14101
rect 7743 14045 7829 14101
rect 7885 14045 7971 14101
rect 8027 14045 8113 14101
rect 8169 14045 8255 14101
rect 8311 14045 8397 14101
rect 8453 14045 8539 14101
rect 8595 14045 8681 14101
rect 8737 14045 8823 14101
rect 8879 14045 8965 14101
rect 9021 14045 9107 14101
rect 9163 14045 9249 14101
rect 9305 14045 9391 14101
rect 9447 14045 9533 14101
rect 9589 14045 9675 14101
rect 9731 14045 9817 14101
rect 9873 14045 9959 14101
rect 10015 14045 10101 14101
rect 10157 14045 10243 14101
rect 10299 14045 10385 14101
rect 10441 14045 10527 14101
rect 10583 14045 10669 14101
rect 10725 14045 10811 14101
rect 10867 14045 10953 14101
rect 11009 14045 11095 14101
rect 11151 14045 11237 14101
rect 11293 14045 11379 14101
rect 11435 14045 11521 14101
rect 11577 14045 11663 14101
rect 11719 14045 11805 14101
rect 11861 14045 11947 14101
rect 12003 14045 12089 14101
rect 12145 14045 12231 14101
rect 12287 14045 12373 14101
rect 12429 14045 12515 14101
rect 12571 14045 12657 14101
rect 12713 14045 12799 14101
rect 12855 14045 12941 14101
rect 12997 14045 13083 14101
rect 13139 14045 13225 14101
rect 13281 14045 13367 14101
rect 13423 14045 13509 14101
rect 13565 14045 13651 14101
rect 13707 14045 13793 14101
rect 13849 14045 13935 14101
rect 13991 14045 14077 14101
rect 14133 14045 14219 14101
rect 14275 14045 14361 14101
rect 14417 14045 14503 14101
rect 14559 14045 14645 14101
rect 14701 14045 14787 14101
rect 14843 14045 15000 14101
rect 0 14000 15000 14045
use 3LM_METAL_RAIL  3LM_METAL_RAIL_0
timestamp 1586916644
transform 1 0 0 0 1 0
box -32 13097 15032 69968
<< labels >>
rlabel metal4 s 763 15661 763 15661 4 DVSS
port 1 nsew
rlabel metal4 s 716 18832 716 18832 4 DVSS
port 1 nsew
rlabel metal4 s 785 21818 785 21818 4 DVSS
port 1 nsew
rlabel metal4 s 785 24195 785 24195 4 DVDD
port 2 nsew
rlabel metal4 s 785 26011 785 26011 4 DVSS
port 1 nsew
rlabel metal4 s 785 28305 785 28305 4 DVDD
port 2 nsew
rlabel metal4 s 785 31520 785 31520 4 DVDD
port 2 nsew
rlabel metal4 s 785 34634 785 34634 4 DVDD
port 2 nsew
rlabel metal4 s 785 37870 785 37870 4 DVDD
port 2 nsew
rlabel metal4 s 785 40253 785 40253 4 DVSS
port 1 nsew
rlabel metal4 s 785 41888 785 41888 4 DVDD
port 2 nsew
rlabel metal4 s 785 44279 785 44279 4 DVDD
port 2 nsew
rlabel metal4 s 785 47506 785 47506 4 DVSS
port 1 nsew
rlabel metal4 s 785 49934 785 49934 4 VSS
port 3 nsew
rlabel metal4 s 785 51369 785 51369 4 VDD
port 4 nsew
rlabel metal4 s 785 53134 785 53134 4 DVDD
port 2 nsew
rlabel metal4 s 785 54569 785 54569 4 DVDD
port 2 nsew
rlabel metal4 s 785 56334 785 56334 4 DVDD
port 2 nsew
rlabel metal4 s 785 57769 785 57769 4 DVSS
port 1 nsew
rlabel metal4 s 785 59534 785 59534 4 DVDD
port 2 nsew
rlabel metal4 s 785 60969 785 60969 4 DVSS
port 1 nsew
rlabel metal4 s 785 62734 785 62734 4 VDD
port 4 nsew
rlabel metal4 s 785 64169 785 64169 4 VSS
port 3 nsew
rlabel metal4 s 785 65934 785 65934 4 DVSS
port 1 nsew
rlabel metal4 s 785 67369 785 67369 4 DVDD
port 2 nsew
rlabel metal4 s 785 68960 785 68960 4 DVSS
port 1 nsew
<< end >>
