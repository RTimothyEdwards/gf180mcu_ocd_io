VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_ocd_io__cor
  CLASS PAD SPACER ;
  FOREIGN gf180mcu_ocd_io__cor ;
  ORIGIN 0.000 0.000 ;
  SIZE 355.000 BY 355.000 ;
  SYMMETRY X Y R90 ;
  SITE GF_IO_Site ;
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 350.000 166.000 355.000 181.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 350.000 150.000 355.000 165.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 350.000 134.000 355.000 149.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 350.000 118.000 355.000 125.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 350.000 206.000 355.000 213.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 350.000 182.000 355.000 197.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 182.000 350.000 197.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 166.000 350.000 181.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 150.000 350.000 165.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 134.000 350.000 149.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 118.000 350.000 125.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 206.000 350.000 213.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 294.000 350.000 301.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 278.000 350.000 285.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 270.000 350.000 277.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 262.000 350.000 269.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 214.000 350.000 229.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 350.000 334.000 355.000 341.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 350.000 294.000 355.000 301.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 350.000 278.000 355.000 285.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 350.000 270.000 355.000 277.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 350.000 262.000 355.000 269.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 350.000 214.000 355.000 228.995 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 334.000 350.000 341.000 355.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 350.000 198.000 355.000 205.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 350.000 126.000 355.000 133.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 350.000 102.000 355.000 117.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 350.000 70.000 355.000 85.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 350.000 86.000 355.000 101.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 126.000 350.000 133.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 102.000 350.000 117.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 86.000 350.000 101.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 70.000 350.000 85.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 198.000 350.000 205.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 326.000 350.000 333.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 302.000 350.000 309.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 286.000 350.000 293.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 230.000 350.000 245.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 350.000 342.000 355.000 348.390 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 350.000 326.000 355.000 333.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 350.000 302.000 355.000 309.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 350.000 286.000 355.000 293.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 350.000 230.000 355.000 245.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 342.000 350.000 348.390 355.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 310.000 350.000 317.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 254.000 350.000 261.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 350.000 310.000 355.000 317.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 350.000 254.000 355.000 261.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 318.000 350.000 325.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 246.000 350.000 253.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 350.000 246.000 355.000 253.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 350.000 318.000 355.000 325.000 ;
    END
  END VSS
  OBS
      LAYER Nwell ;
        RECT 67.560 67.500 350.445 352.170 ;
      LAYER Metal1 ;
        RECT 65.540 65.540 355.000 355.000 ;
      LAYER Metal2 ;
        RECT 68.030 67.970 354.505 354.450 ;
      LAYER Metal3 ;
        RECT 70.000 70.000 355.000 355.000 ;
      LAYER Metal4 ;
        RECT 348.990 349.400 350.000 350.000 ;
        RECT 70.000 348.990 350.000 349.400 ;
        RECT 70.000 70.000 349.400 348.990 ;
  END
END gf180mcu_ocd_io__cor
END LIBRARY

