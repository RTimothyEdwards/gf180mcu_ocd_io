magic
tech gf180mcuD
magscale 1 10
timestamp 1758746585
<< isosubstrate >>
rect 251 53100 14727 57210
rect 2457 47163 12521 53100
rect 601 42936 14377 47163
rect 957 26552 12844 42936
rect 957 1096 14021 26552
<< nwell >>
rect 2457 52160 12521 52716
rect 2457 48116 3013 52160
rect 11965 48116 12521 52160
rect 2457 47560 12521 48116
<< pwell >>
rect 747 53655 3923 56655
rect 4183 53655 7359 56655
rect 7619 53655 10795 56655
rect 11055 53655 14231 56655
<< mvndiff >>
rect 747 56618 835 56655
rect 747 53692 760 56618
rect 806 53692 835 56618
rect 747 53655 835 53692
rect 3835 56618 3923 56655
rect 3835 53692 3864 56618
rect 3910 53692 3923 56618
rect 3835 53655 3923 53692
rect 4183 56618 4271 56655
rect 4183 53692 4196 56618
rect 4242 53692 4271 56618
rect 4183 53655 4271 53692
rect 7271 56618 7359 56655
rect 7271 53692 7300 56618
rect 7346 53692 7359 56618
rect 7271 53655 7359 53692
rect 7619 56618 7707 56655
rect 7619 53692 7632 56618
rect 7678 53692 7707 56618
rect 7619 53655 7707 53692
rect 10707 56618 10795 56655
rect 10707 53692 10736 56618
rect 10782 53692 10795 56618
rect 10707 53655 10795 53692
rect 11055 56618 11143 56655
rect 11055 53692 11068 56618
rect 11114 53692 11143 56618
rect 11055 53655 11143 53692
rect 14143 56618 14231 56655
rect 14143 53692 14172 56618
rect 14218 53692 14231 56618
rect 14143 53655 14231 53692
<< mvndiffc >>
rect 760 53692 806 56618
rect 3864 53692 3910 56618
rect 4196 53692 4242 56618
rect 7300 53692 7346 56618
rect 7632 53692 7678 56618
rect 10736 53692 10782 56618
rect 11068 53692 11114 56618
rect 14172 53692 14218 56618
<< psubdiff >>
rect 334 57105 14644 57127
rect 334 53205 356 57105
rect 402 57059 510 57105
rect 14468 57059 14576 57105
rect 402 57037 14576 57059
rect 402 53273 424 57037
rect 14554 53273 14576 57037
rect 402 53251 14576 53273
rect 402 53205 510 53251
rect 14468 53205 14576 53251
rect 14622 53205 14644 57105
rect 334 53183 14644 53205
rect 246 52611 2236 52633
rect 246 47665 268 52611
rect 2214 47665 2236 52611
rect 246 47643 2236 47665
rect 3094 52029 11884 52051
rect 3094 51983 3142 52029
rect 11836 51983 11884 52029
rect 3094 51900 11884 51983
rect 3094 48376 3116 51900
rect 3162 51875 11816 51900
rect 3162 51844 3424 51875
rect 3162 51234 3270 51844
rect 3316 51829 3424 51844
rect 11554 51844 11816 51875
rect 11554 51829 11662 51844
rect 3316 51807 11662 51829
rect 3316 51271 3338 51807
rect 11640 51271 11662 51807
rect 3316 51249 11662 51271
rect 3316 51234 3424 51249
rect 3162 51203 3424 51234
rect 11554 51234 11662 51249
rect 11708 51234 11816 51844
rect 11554 51203 11816 51234
rect 3162 51095 11816 51203
rect 3162 51049 3330 51095
rect 11648 51049 11816 51095
rect 3162 50941 11816 51049
rect 3162 50910 3424 50941
rect 3162 50300 3270 50910
rect 3316 50895 3424 50910
rect 11554 50910 11816 50941
rect 11554 50895 11662 50910
rect 3316 50873 11662 50895
rect 3316 50337 3338 50873
rect 11640 50337 11662 50873
rect 3316 50315 11662 50337
rect 3316 50300 3424 50315
rect 3162 50269 3424 50300
rect 11554 50300 11662 50315
rect 11708 50300 11816 50910
rect 11554 50269 11816 50300
rect 3162 50161 11816 50269
rect 3162 50115 3330 50161
rect 11648 50115 11816 50161
rect 3162 50007 11816 50115
rect 3162 49976 3424 50007
rect 3162 49366 3270 49976
rect 3316 49961 3424 49976
rect 11554 49976 11816 50007
rect 11554 49961 11662 49976
rect 3316 49939 11662 49961
rect 3316 49403 3338 49939
rect 11640 49403 11662 49939
rect 3316 49381 11662 49403
rect 3316 49366 3424 49381
rect 3162 49335 3424 49366
rect 11554 49366 11662 49381
rect 11708 49366 11816 49976
rect 11554 49335 11816 49366
rect 3162 49227 11816 49335
rect 3162 49181 3330 49227
rect 11648 49181 11816 49227
rect 3162 49073 11816 49181
rect 3162 49042 3424 49073
rect 3162 48432 3270 49042
rect 3316 49027 3424 49042
rect 11554 49042 11816 49073
rect 11554 49027 11662 49042
rect 3316 49005 11662 49027
rect 3316 48469 3338 49005
rect 11640 48469 11662 49005
rect 3316 48447 11662 48469
rect 3316 48432 3424 48447
rect 3162 48401 3424 48432
rect 11554 48432 11662 48447
rect 11708 48432 11816 49042
rect 11554 48401 11816 48432
rect 3162 48376 11816 48401
rect 11862 48376 11884 51900
rect 3094 48293 11884 48376
rect 3094 48247 3142 48293
rect 11836 48247 11884 48293
rect 3094 48225 11884 48247
rect 12742 52611 14732 52633
rect 12742 47665 12764 52611
rect 14710 47665 14732 52611
rect 12742 47643 14732 47665
rect 246 42647 736 42669
rect 246 1201 268 42647
rect 714 1201 736 42647
rect 13001 42647 13991 42669
rect 13001 27201 13023 42647
rect 13969 27201 13991 42647
rect 13001 27179 13991 27201
rect 14242 42647 14732 42669
rect 246 1179 736 1201
rect 14242 1201 14264 42647
rect 14710 1201 14732 42647
rect 14242 1179 14732 1201
<< nsubdiff >>
rect 2540 52611 12438 52633
rect 2540 47665 2562 52611
rect 2908 52265 3016 52611
rect 11962 52265 12070 52611
rect 2908 52243 12070 52265
rect 2908 48033 2930 52243
rect 12048 48033 12070 52243
rect 2908 48011 12070 48033
rect 2908 47665 3016 48011
rect 11962 47665 12070 48011
rect 12416 47665 12438 52611
rect 2540 47643 12438 47665
<< psubdiffcont >>
rect 356 53205 402 57105
rect 510 57059 14468 57105
rect 510 53205 14468 53251
rect 14576 53205 14622 57105
rect 268 47665 2214 52611
rect 3142 51983 11836 52029
rect 3116 48376 3162 51900
rect 3270 51234 3316 51844
rect 3424 51829 11554 51875
rect 3424 51203 11554 51249
rect 11662 51234 11708 51844
rect 3330 51049 11648 51095
rect 3270 50300 3316 50910
rect 3424 50895 11554 50941
rect 3424 50269 11554 50315
rect 11662 50300 11708 50910
rect 3330 50115 11648 50161
rect 3270 49366 3316 49976
rect 3424 49961 11554 50007
rect 3424 49335 11554 49381
rect 11662 49366 11708 49976
rect 3330 49181 11648 49227
rect 3270 48432 3316 49042
rect 3424 49027 11554 49073
rect 3424 48401 11554 48447
rect 11662 48432 11708 49042
rect 11816 48376 11862 51900
rect 3142 48247 11836 48293
rect 12764 47665 14710 52611
rect 268 1201 714 42647
rect 13023 27201 13969 42647
rect 14264 1201 14710 42647
<< nsubdiffcont >>
rect 2562 47665 2908 52611
rect 3016 52265 11962 52611
rect 3016 47665 11962 48011
rect 12070 47665 12416 52611
<< mvnmoscap >>
rect 835 53655 3835 56655
rect 4271 53655 7271 56655
rect 7707 53655 10707 56655
rect 11143 53655 14143 56655
<< polysilicon >>
rect 835 56734 3835 56747
rect 835 56688 888 56734
rect 3782 56688 3835 56734
rect 835 56655 3835 56688
rect 4271 56734 7271 56747
rect 4271 56688 4324 56734
rect 7218 56688 7271 56734
rect 4271 56655 7271 56688
rect 7707 56734 10707 56747
rect 7707 56688 7760 56734
rect 10654 56688 10707 56734
rect 7707 56655 10707 56688
rect 11143 56734 14143 56747
rect 11143 56688 11196 56734
rect 14090 56688 14143 56734
rect 11143 56655 14143 56688
rect 835 53622 3835 53655
rect 835 53576 888 53622
rect 3782 53576 3835 53622
rect 835 53563 3835 53576
rect 4271 53622 7271 53655
rect 4271 53576 4324 53622
rect 7218 53576 7271 53622
rect 4271 53563 7271 53576
rect 7707 53622 10707 53655
rect 7707 53576 7760 53622
rect 10654 53576 10707 53622
rect 7707 53563 10707 53576
rect 11143 53622 14143 53655
rect 11143 53576 11196 53622
rect 14090 53576 14143 53622
rect 11143 53563 14143 53576
<< polycontact >>
rect 888 56688 3782 56734
rect 4324 56688 7218 56734
rect 7760 56688 10654 56734
rect 11196 56688 14090 56734
rect 888 53576 3782 53622
rect 4324 53576 7218 53622
rect 7760 53576 10654 53622
rect 11196 53576 14090 53622
<< mvndiode >>
rect 3489 51626 11489 51639
rect 3489 51580 3502 51626
rect 11476 51580 11489 51626
rect 3489 51498 11489 51580
rect 3489 51452 3502 51498
rect 11476 51452 11489 51498
rect 3489 51439 11489 51452
rect 3489 50692 11489 50705
rect 3489 50646 3502 50692
rect 11476 50646 11489 50692
rect 3489 50564 11489 50646
rect 3489 50518 3502 50564
rect 11476 50518 11489 50564
rect 3489 50505 11489 50518
rect 3489 49758 11489 49771
rect 3489 49712 3502 49758
rect 11476 49712 11489 49758
rect 3489 49630 11489 49712
rect 3489 49584 3502 49630
rect 11476 49584 11489 49630
rect 3489 49571 11489 49584
rect 3489 48824 11489 48837
rect 3489 48778 3502 48824
rect 11476 48778 11489 48824
rect 3489 48696 11489 48778
rect 3489 48650 3502 48696
rect 11476 48650 11489 48696
rect 3489 48637 11489 48650
<< mvndiodec >>
rect 3502 51580 11476 51626
rect 3502 51452 11476 51498
rect 3502 50646 11476 50692
rect 3502 50518 11476 50564
rect 3502 49712 11476 49758
rect 3502 49584 11476 49630
rect 3502 48778 11476 48824
rect 3502 48650 11476 48696
<< metal1 >>
rect 2489 57116 2673 57120
rect 4859 57116 5043 57120
rect 7235 57116 7743 57120
rect 9935 57116 10119 57120
rect 12305 57116 12489 57120
rect 345 57108 14633 57116
rect 345 57105 2501 57108
rect 2553 57105 2609 57108
rect 2661 57105 4871 57108
rect 4923 57105 4979 57108
rect 5031 57105 7247 57108
rect 7299 57105 7355 57108
rect 7407 57105 7463 57108
rect 7515 57105 7571 57108
rect 7623 57105 7679 57108
rect 7731 57105 9947 57108
rect 9999 57105 10055 57108
rect 10107 57105 12317 57108
rect 12369 57105 12425 57108
rect 12477 57105 14633 57108
rect 345 53205 356 57105
rect 402 57059 510 57105
rect 14468 57059 14576 57105
rect 402 57056 2501 57059
rect 2553 57056 2609 57059
rect 2661 57056 4871 57059
rect 4923 57056 4979 57059
rect 5031 57056 7247 57059
rect 7299 57056 7355 57059
rect 7407 57056 7463 57059
rect 7515 57056 7571 57059
rect 7623 57056 7679 57059
rect 7731 57056 9947 57059
rect 9999 57056 10055 57059
rect 10107 57056 12317 57059
rect 12369 57056 12425 57059
rect 12477 57056 14576 57059
rect 402 57048 14576 57056
rect 402 56655 413 57048
rect 2489 57044 2673 57048
rect 4859 57044 5043 57048
rect 7235 57044 7743 57048
rect 9935 57044 10119 57048
rect 12305 57044 12489 57048
rect 877 56734 3793 56745
rect 877 56688 888 56734
rect 3782 56688 3793 56734
rect 877 56677 3793 56688
rect 877 56669 1877 56677
rect 402 56618 817 56655
rect 402 53692 760 56618
rect 806 53692 817 56618
rect 402 53505 817 53692
rect 877 56617 917 56669
rect 969 56617 1041 56669
rect 1093 56617 1165 56669
rect 1217 56617 1289 56669
rect 1341 56617 1413 56669
rect 1465 56617 1537 56669
rect 1589 56617 1661 56669
rect 1713 56617 1785 56669
rect 1837 56617 1877 56669
rect 877 56545 1877 56617
rect 877 56493 917 56545
rect 969 56493 1041 56545
rect 1093 56493 1165 56545
rect 1217 56493 1289 56545
rect 1341 56493 1413 56545
rect 1465 56493 1537 56545
rect 1589 56493 1661 56545
rect 1713 56493 1785 56545
rect 1837 56493 1877 56545
rect 877 56421 1877 56493
rect 877 56369 917 56421
rect 969 56369 1041 56421
rect 1093 56369 1165 56421
rect 1217 56369 1289 56421
rect 1341 56369 1413 56421
rect 1465 56369 1537 56421
rect 1589 56369 1661 56421
rect 1713 56369 1785 56421
rect 1837 56369 1877 56421
rect 877 56297 1877 56369
rect 877 56245 917 56297
rect 969 56245 1041 56297
rect 1093 56245 1165 56297
rect 1217 56245 1289 56297
rect 1341 56245 1413 56297
rect 1465 56245 1537 56297
rect 1589 56245 1661 56297
rect 1713 56245 1785 56297
rect 1837 56245 1877 56297
rect 877 56173 1877 56245
rect 877 56121 917 56173
rect 969 56121 1041 56173
rect 1093 56121 1165 56173
rect 1217 56121 1289 56173
rect 1341 56121 1413 56173
rect 1465 56121 1537 56173
rect 1589 56121 1661 56173
rect 1713 56121 1785 56173
rect 1837 56121 1877 56173
rect 877 56049 1877 56121
rect 877 55997 917 56049
rect 969 55997 1041 56049
rect 1093 55997 1165 56049
rect 1217 55997 1289 56049
rect 1341 55997 1413 56049
rect 1465 55997 1537 56049
rect 1589 55997 1661 56049
rect 1713 55997 1785 56049
rect 1837 55997 1877 56049
rect 877 55925 1877 55997
rect 877 55873 917 55925
rect 969 55873 1041 55925
rect 1093 55873 1165 55925
rect 1217 55873 1289 55925
rect 1341 55873 1413 55925
rect 1465 55873 1537 55925
rect 1589 55873 1661 55925
rect 1713 55873 1785 55925
rect 1837 55873 1877 55925
rect 877 55801 1877 55873
rect 877 55749 917 55801
rect 969 55749 1041 55801
rect 1093 55749 1165 55801
rect 1217 55749 1289 55801
rect 1341 55749 1413 55801
rect 1465 55749 1537 55801
rect 1589 55749 1661 55801
rect 1713 55749 1785 55801
rect 1837 55749 1877 55801
rect 877 55677 1877 55749
rect 877 55625 917 55677
rect 969 55625 1041 55677
rect 1093 55625 1165 55677
rect 1217 55625 1289 55677
rect 1341 55625 1413 55677
rect 1465 55625 1537 55677
rect 1589 55625 1661 55677
rect 1713 55625 1785 55677
rect 1837 55625 1877 55677
rect 877 55553 1877 55625
rect 877 55501 917 55553
rect 969 55501 1041 55553
rect 1093 55501 1165 55553
rect 1217 55501 1289 55553
rect 1341 55501 1413 55553
rect 1465 55501 1537 55553
rect 1589 55501 1661 55553
rect 1713 55501 1785 55553
rect 1837 55501 1877 55553
rect 877 55429 1877 55501
rect 877 55377 917 55429
rect 969 55377 1041 55429
rect 1093 55377 1165 55429
rect 1217 55377 1289 55429
rect 1341 55377 1413 55429
rect 1465 55377 1537 55429
rect 1589 55377 1661 55429
rect 1713 55377 1785 55429
rect 1837 55377 1877 55429
rect 877 55305 1877 55377
rect 877 55253 917 55305
rect 969 55253 1041 55305
rect 1093 55253 1165 55305
rect 1217 55253 1289 55305
rect 1341 55253 1413 55305
rect 1465 55253 1537 55305
rect 1589 55253 1661 55305
rect 1713 55253 1785 55305
rect 1837 55253 1877 55305
rect 877 55181 1877 55253
rect 877 55129 917 55181
rect 969 55129 1041 55181
rect 1093 55129 1165 55181
rect 1217 55129 1289 55181
rect 1341 55129 1413 55181
rect 1465 55129 1537 55181
rect 1589 55129 1661 55181
rect 1713 55129 1785 55181
rect 1837 55129 1877 55181
rect 877 55057 1877 55129
rect 877 55005 917 55057
rect 969 55005 1041 55057
rect 1093 55005 1165 55057
rect 1217 55005 1289 55057
rect 1341 55005 1413 55057
rect 1465 55005 1537 55057
rect 1589 55005 1661 55057
rect 1713 55005 1785 55057
rect 1837 55005 1877 55057
rect 877 54933 1877 55005
rect 877 54881 917 54933
rect 969 54881 1041 54933
rect 1093 54881 1165 54933
rect 1217 54881 1289 54933
rect 1341 54881 1413 54933
rect 1465 54881 1537 54933
rect 1589 54881 1661 54933
rect 1713 54881 1785 54933
rect 1837 54881 1877 54933
rect 877 54809 1877 54881
rect 877 54757 917 54809
rect 969 54757 1041 54809
rect 1093 54757 1165 54809
rect 1217 54757 1289 54809
rect 1341 54757 1413 54809
rect 1465 54757 1537 54809
rect 1589 54757 1661 54809
rect 1713 54757 1785 54809
rect 1837 54757 1877 54809
rect 877 54685 1877 54757
rect 877 54633 917 54685
rect 969 54633 1041 54685
rect 1093 54633 1165 54685
rect 1217 54633 1289 54685
rect 1341 54633 1413 54685
rect 1465 54633 1537 54685
rect 1589 54633 1661 54685
rect 1713 54633 1785 54685
rect 1837 54633 1877 54685
rect 877 54561 1877 54633
rect 877 54509 917 54561
rect 969 54509 1041 54561
rect 1093 54509 1165 54561
rect 1217 54509 1289 54561
rect 1341 54509 1413 54561
rect 1465 54509 1537 54561
rect 1589 54509 1661 54561
rect 1713 54509 1785 54561
rect 1837 54509 1877 54561
rect 877 54437 1877 54509
rect 877 54385 917 54437
rect 969 54385 1041 54437
rect 1093 54385 1165 54437
rect 1217 54385 1289 54437
rect 1341 54385 1413 54437
rect 1465 54385 1537 54437
rect 1589 54385 1661 54437
rect 1713 54385 1785 54437
rect 1837 54385 1877 54437
rect 877 54313 1877 54385
rect 877 54261 917 54313
rect 969 54261 1041 54313
rect 1093 54261 1165 54313
rect 1217 54261 1289 54313
rect 1341 54261 1413 54313
rect 1465 54261 1537 54313
rect 1589 54261 1661 54313
rect 1713 54261 1785 54313
rect 1837 54261 1877 54313
rect 877 54189 1877 54261
rect 877 54137 917 54189
rect 969 54137 1041 54189
rect 1093 54137 1165 54189
rect 1217 54137 1289 54189
rect 1341 54137 1413 54189
rect 1465 54137 1537 54189
rect 1589 54137 1661 54189
rect 1713 54137 1785 54189
rect 1837 54137 1877 54189
rect 877 54065 1877 54137
rect 877 54013 917 54065
rect 969 54013 1041 54065
rect 1093 54013 1165 54065
rect 1217 54013 1289 54065
rect 1341 54013 1413 54065
rect 1465 54013 1537 54065
rect 1589 54013 1661 54065
rect 1713 54013 1785 54065
rect 1837 54013 1877 54065
rect 877 53941 1877 54013
rect 877 53889 917 53941
rect 969 53889 1041 53941
rect 1093 53889 1165 53941
rect 1217 53889 1289 53941
rect 1341 53889 1413 53941
rect 1465 53889 1537 53941
rect 1589 53889 1661 53941
rect 1713 53889 1785 53941
rect 1837 53889 1877 53941
rect 877 53817 1877 53889
rect 877 53765 917 53817
rect 969 53765 1041 53817
rect 1093 53765 1165 53817
rect 1217 53765 1289 53817
rect 1341 53765 1413 53817
rect 1465 53765 1537 53817
rect 1589 53765 1661 53817
rect 1713 53765 1785 53817
rect 1837 53765 1877 53817
rect 877 53693 1877 53765
rect 877 53641 917 53693
rect 969 53641 1041 53693
rect 1093 53641 1165 53693
rect 1217 53641 1289 53693
rect 1341 53641 1413 53693
rect 1465 53641 1537 53693
rect 1589 53641 1661 53693
rect 1713 53641 1785 53693
rect 1837 53641 1877 53693
rect 877 53633 1877 53641
rect 2793 56669 3793 56677
rect 2793 56617 2833 56669
rect 2885 56617 2957 56669
rect 3009 56617 3081 56669
rect 3133 56617 3205 56669
rect 3257 56617 3329 56669
rect 3381 56617 3453 56669
rect 3505 56617 3577 56669
rect 3629 56617 3701 56669
rect 3753 56617 3793 56669
rect 4313 56734 7229 56745
rect 4313 56688 4324 56734
rect 7218 56688 7229 56734
rect 4313 56677 7229 56688
rect 4313 56669 5313 56677
rect 2793 56545 3793 56617
rect 2793 56493 2833 56545
rect 2885 56493 2957 56545
rect 3009 56493 3081 56545
rect 3133 56493 3205 56545
rect 3257 56493 3329 56545
rect 3381 56493 3453 56545
rect 3505 56493 3577 56545
rect 3629 56493 3701 56545
rect 3753 56493 3793 56545
rect 2793 56421 3793 56493
rect 2793 56369 2833 56421
rect 2885 56369 2957 56421
rect 3009 56369 3081 56421
rect 3133 56369 3205 56421
rect 3257 56369 3329 56421
rect 3381 56369 3453 56421
rect 3505 56369 3577 56421
rect 3629 56369 3701 56421
rect 3753 56369 3793 56421
rect 2793 56297 3793 56369
rect 2793 56245 2833 56297
rect 2885 56245 2957 56297
rect 3009 56245 3081 56297
rect 3133 56245 3205 56297
rect 3257 56245 3329 56297
rect 3381 56245 3453 56297
rect 3505 56245 3577 56297
rect 3629 56245 3701 56297
rect 3753 56245 3793 56297
rect 2793 56173 3793 56245
rect 2793 56121 2833 56173
rect 2885 56121 2957 56173
rect 3009 56121 3081 56173
rect 3133 56121 3205 56173
rect 3257 56121 3329 56173
rect 3381 56121 3453 56173
rect 3505 56121 3577 56173
rect 3629 56121 3701 56173
rect 3753 56121 3793 56173
rect 2793 56049 3793 56121
rect 2793 55997 2833 56049
rect 2885 55997 2957 56049
rect 3009 55997 3081 56049
rect 3133 55997 3205 56049
rect 3257 55997 3329 56049
rect 3381 55997 3453 56049
rect 3505 55997 3577 56049
rect 3629 55997 3701 56049
rect 3753 55997 3793 56049
rect 2793 55925 3793 55997
rect 2793 55873 2833 55925
rect 2885 55873 2957 55925
rect 3009 55873 3081 55925
rect 3133 55873 3205 55925
rect 3257 55873 3329 55925
rect 3381 55873 3453 55925
rect 3505 55873 3577 55925
rect 3629 55873 3701 55925
rect 3753 55873 3793 55925
rect 2793 55801 3793 55873
rect 2793 55749 2833 55801
rect 2885 55749 2957 55801
rect 3009 55749 3081 55801
rect 3133 55749 3205 55801
rect 3257 55749 3329 55801
rect 3381 55749 3453 55801
rect 3505 55749 3577 55801
rect 3629 55749 3701 55801
rect 3753 55749 3793 55801
rect 2793 55677 3793 55749
rect 2793 55625 2833 55677
rect 2885 55625 2957 55677
rect 3009 55625 3081 55677
rect 3133 55625 3205 55677
rect 3257 55625 3329 55677
rect 3381 55625 3453 55677
rect 3505 55625 3577 55677
rect 3629 55625 3701 55677
rect 3753 55625 3793 55677
rect 2793 55553 3793 55625
rect 2793 55501 2833 55553
rect 2885 55501 2957 55553
rect 3009 55501 3081 55553
rect 3133 55501 3205 55553
rect 3257 55501 3329 55553
rect 3381 55501 3453 55553
rect 3505 55501 3577 55553
rect 3629 55501 3701 55553
rect 3753 55501 3793 55553
rect 2793 55429 3793 55501
rect 2793 55377 2833 55429
rect 2885 55377 2957 55429
rect 3009 55377 3081 55429
rect 3133 55377 3205 55429
rect 3257 55377 3329 55429
rect 3381 55377 3453 55429
rect 3505 55377 3577 55429
rect 3629 55377 3701 55429
rect 3753 55377 3793 55429
rect 2793 55305 3793 55377
rect 2793 55253 2833 55305
rect 2885 55253 2957 55305
rect 3009 55253 3081 55305
rect 3133 55253 3205 55305
rect 3257 55253 3329 55305
rect 3381 55253 3453 55305
rect 3505 55253 3577 55305
rect 3629 55253 3701 55305
rect 3753 55253 3793 55305
rect 2793 55181 3793 55253
rect 2793 55129 2833 55181
rect 2885 55129 2957 55181
rect 3009 55129 3081 55181
rect 3133 55129 3205 55181
rect 3257 55129 3329 55181
rect 3381 55129 3453 55181
rect 3505 55129 3577 55181
rect 3629 55129 3701 55181
rect 3753 55129 3793 55181
rect 2793 55057 3793 55129
rect 2793 55005 2833 55057
rect 2885 55005 2957 55057
rect 3009 55005 3081 55057
rect 3133 55005 3205 55057
rect 3257 55005 3329 55057
rect 3381 55005 3453 55057
rect 3505 55005 3577 55057
rect 3629 55005 3701 55057
rect 3753 55005 3793 55057
rect 2793 54933 3793 55005
rect 2793 54881 2833 54933
rect 2885 54881 2957 54933
rect 3009 54881 3081 54933
rect 3133 54881 3205 54933
rect 3257 54881 3329 54933
rect 3381 54881 3453 54933
rect 3505 54881 3577 54933
rect 3629 54881 3701 54933
rect 3753 54881 3793 54933
rect 2793 54809 3793 54881
rect 2793 54757 2833 54809
rect 2885 54757 2957 54809
rect 3009 54757 3081 54809
rect 3133 54757 3205 54809
rect 3257 54757 3329 54809
rect 3381 54757 3453 54809
rect 3505 54757 3577 54809
rect 3629 54757 3701 54809
rect 3753 54757 3793 54809
rect 2793 54685 3793 54757
rect 2793 54633 2833 54685
rect 2885 54633 2957 54685
rect 3009 54633 3081 54685
rect 3133 54633 3205 54685
rect 3257 54633 3329 54685
rect 3381 54633 3453 54685
rect 3505 54633 3577 54685
rect 3629 54633 3701 54685
rect 3753 54633 3793 54685
rect 2793 54561 3793 54633
rect 2793 54509 2833 54561
rect 2885 54509 2957 54561
rect 3009 54509 3081 54561
rect 3133 54509 3205 54561
rect 3257 54509 3329 54561
rect 3381 54509 3453 54561
rect 3505 54509 3577 54561
rect 3629 54509 3701 54561
rect 3753 54509 3793 54561
rect 2793 54437 3793 54509
rect 2793 54385 2833 54437
rect 2885 54385 2957 54437
rect 3009 54385 3081 54437
rect 3133 54385 3205 54437
rect 3257 54385 3329 54437
rect 3381 54385 3453 54437
rect 3505 54385 3577 54437
rect 3629 54385 3701 54437
rect 3753 54385 3793 54437
rect 2793 54313 3793 54385
rect 2793 54261 2833 54313
rect 2885 54261 2957 54313
rect 3009 54261 3081 54313
rect 3133 54261 3205 54313
rect 3257 54261 3329 54313
rect 3381 54261 3453 54313
rect 3505 54261 3577 54313
rect 3629 54261 3701 54313
rect 3753 54261 3793 54313
rect 2793 54189 3793 54261
rect 2793 54137 2833 54189
rect 2885 54137 2957 54189
rect 3009 54137 3081 54189
rect 3133 54137 3205 54189
rect 3257 54137 3329 54189
rect 3381 54137 3453 54189
rect 3505 54137 3577 54189
rect 3629 54137 3701 54189
rect 3753 54137 3793 54189
rect 2793 54065 3793 54137
rect 2793 54013 2833 54065
rect 2885 54013 2957 54065
rect 3009 54013 3081 54065
rect 3133 54013 3205 54065
rect 3257 54013 3329 54065
rect 3381 54013 3453 54065
rect 3505 54013 3577 54065
rect 3629 54013 3701 54065
rect 3753 54013 3793 54065
rect 2793 53941 3793 54013
rect 2793 53889 2833 53941
rect 2885 53889 2957 53941
rect 3009 53889 3081 53941
rect 3133 53889 3205 53941
rect 3257 53889 3329 53941
rect 3381 53889 3453 53941
rect 3505 53889 3577 53941
rect 3629 53889 3701 53941
rect 3753 53889 3793 53941
rect 2793 53817 3793 53889
rect 2793 53765 2833 53817
rect 2885 53765 2957 53817
rect 3009 53765 3081 53817
rect 3133 53765 3205 53817
rect 3257 53765 3329 53817
rect 3381 53765 3453 53817
rect 3505 53765 3577 53817
rect 3629 53765 3701 53817
rect 3753 53765 3793 53817
rect 2793 53693 3793 53765
rect 2793 53641 2833 53693
rect 2885 53641 2957 53693
rect 3009 53641 3081 53693
rect 3133 53641 3205 53693
rect 3257 53641 3329 53693
rect 3381 53641 3453 53693
rect 3505 53641 3577 53693
rect 3629 53641 3701 53693
rect 3753 53641 3793 53693
rect 2793 53633 3793 53641
rect 877 53622 3793 53633
rect 877 53576 888 53622
rect 3782 53576 3793 53622
rect 877 53565 3793 53576
rect 3853 56618 4253 56655
rect 3853 53692 3864 56618
rect 3910 53692 4196 56618
rect 4242 53692 4253 56618
rect 3853 53505 4253 53692
rect 4313 56617 4340 56669
rect 4392 56617 4464 56669
rect 4516 56617 4588 56669
rect 4640 56617 4712 56669
rect 4764 56617 5313 56669
rect 4313 56545 5313 56617
rect 4313 56493 4340 56545
rect 4392 56493 4464 56545
rect 4516 56493 4588 56545
rect 4640 56493 4712 56545
rect 4764 56493 5313 56545
rect 4313 56421 5313 56493
rect 4313 56369 4340 56421
rect 4392 56369 4464 56421
rect 4516 56369 4588 56421
rect 4640 56369 4712 56421
rect 4764 56369 5313 56421
rect 4313 56297 5313 56369
rect 4313 56245 4340 56297
rect 4392 56245 4464 56297
rect 4516 56245 4588 56297
rect 4640 56245 4712 56297
rect 4764 56245 5313 56297
rect 4313 56173 5313 56245
rect 4313 56121 4340 56173
rect 4392 56121 4464 56173
rect 4516 56121 4588 56173
rect 4640 56121 4712 56173
rect 4764 56121 5313 56173
rect 4313 56049 5313 56121
rect 4313 55997 4340 56049
rect 4392 55997 4464 56049
rect 4516 55997 4588 56049
rect 4640 55997 4712 56049
rect 4764 55997 5313 56049
rect 4313 55925 5313 55997
rect 4313 55873 4340 55925
rect 4392 55873 4464 55925
rect 4516 55873 4588 55925
rect 4640 55873 4712 55925
rect 4764 55873 5313 55925
rect 4313 55801 5313 55873
rect 4313 55749 4340 55801
rect 4392 55749 4464 55801
rect 4516 55749 4588 55801
rect 4640 55749 4712 55801
rect 4764 55749 5313 55801
rect 4313 55677 5313 55749
rect 4313 55625 4340 55677
rect 4392 55625 4464 55677
rect 4516 55625 4588 55677
rect 4640 55625 4712 55677
rect 4764 55625 5313 55677
rect 4313 55553 5313 55625
rect 4313 55501 4340 55553
rect 4392 55501 4464 55553
rect 4516 55501 4588 55553
rect 4640 55501 4712 55553
rect 4764 55501 5313 55553
rect 4313 55429 5313 55501
rect 4313 55377 4340 55429
rect 4392 55377 4464 55429
rect 4516 55377 4588 55429
rect 4640 55377 4712 55429
rect 4764 55377 5313 55429
rect 4313 55305 5313 55377
rect 4313 55253 4340 55305
rect 4392 55253 4464 55305
rect 4516 55253 4588 55305
rect 4640 55253 4712 55305
rect 4764 55253 5313 55305
rect 4313 55181 5313 55253
rect 4313 55129 4340 55181
rect 4392 55129 4464 55181
rect 4516 55129 4588 55181
rect 4640 55129 4712 55181
rect 4764 55129 5313 55181
rect 4313 55057 5313 55129
rect 4313 55005 4340 55057
rect 4392 55005 4464 55057
rect 4516 55005 4588 55057
rect 4640 55005 4712 55057
rect 4764 55005 5313 55057
rect 4313 54933 5313 55005
rect 4313 54881 4340 54933
rect 4392 54881 4464 54933
rect 4516 54881 4588 54933
rect 4640 54881 4712 54933
rect 4764 54881 5313 54933
rect 4313 54809 5313 54881
rect 4313 54757 4340 54809
rect 4392 54757 4464 54809
rect 4516 54757 4588 54809
rect 4640 54757 4712 54809
rect 4764 54757 5313 54809
rect 4313 54685 5313 54757
rect 4313 54633 4340 54685
rect 4392 54633 4464 54685
rect 4516 54633 4588 54685
rect 4640 54633 4712 54685
rect 4764 54633 5313 54685
rect 4313 54561 5313 54633
rect 4313 54509 4340 54561
rect 4392 54509 4464 54561
rect 4516 54509 4588 54561
rect 4640 54509 4712 54561
rect 4764 54509 5313 54561
rect 4313 54437 5313 54509
rect 4313 54385 4340 54437
rect 4392 54385 4464 54437
rect 4516 54385 4588 54437
rect 4640 54385 4712 54437
rect 4764 54385 5313 54437
rect 4313 54313 5313 54385
rect 4313 54261 4340 54313
rect 4392 54261 4464 54313
rect 4516 54261 4588 54313
rect 4640 54261 4712 54313
rect 4764 54261 5313 54313
rect 4313 54189 5313 54261
rect 4313 54137 4340 54189
rect 4392 54137 4464 54189
rect 4516 54137 4588 54189
rect 4640 54137 4712 54189
rect 4764 54137 5313 54189
rect 4313 54065 5313 54137
rect 4313 54013 4340 54065
rect 4392 54013 4464 54065
rect 4516 54013 4588 54065
rect 4640 54013 4712 54065
rect 4764 54013 5313 54065
rect 4313 53941 5313 54013
rect 4313 53889 4340 53941
rect 4392 53889 4464 53941
rect 4516 53889 4588 53941
rect 4640 53889 4712 53941
rect 4764 53889 5313 53941
rect 4313 53817 5313 53889
rect 4313 53765 4340 53817
rect 4392 53765 4464 53817
rect 4516 53765 4588 53817
rect 4640 53765 4712 53817
rect 4764 53765 5313 53817
rect 4313 53693 5313 53765
rect 4313 53641 4340 53693
rect 4392 53641 4464 53693
rect 4516 53641 4588 53693
rect 4640 53641 4712 53693
rect 4764 53641 5313 53693
rect 4313 53633 5313 53641
rect 6229 56669 7229 56677
rect 6229 56617 6297 56669
rect 6349 56617 6421 56669
rect 6473 56617 6545 56669
rect 6597 56617 6669 56669
rect 6721 56617 6793 56669
rect 6845 56617 6917 56669
rect 6969 56617 7041 56669
rect 7093 56617 7229 56669
rect 7749 56734 10665 56745
rect 7749 56688 7760 56734
rect 10654 56688 10665 56734
rect 7749 56677 10665 56688
rect 7749 56669 8749 56677
rect 6229 56545 7229 56617
rect 6229 56493 6297 56545
rect 6349 56493 6421 56545
rect 6473 56493 6545 56545
rect 6597 56493 6669 56545
rect 6721 56493 6793 56545
rect 6845 56493 6917 56545
rect 6969 56493 7041 56545
rect 7093 56493 7229 56545
rect 6229 56421 7229 56493
rect 6229 56369 6297 56421
rect 6349 56369 6421 56421
rect 6473 56369 6545 56421
rect 6597 56369 6669 56421
rect 6721 56369 6793 56421
rect 6845 56369 6917 56421
rect 6969 56369 7041 56421
rect 7093 56369 7229 56421
rect 6229 56297 7229 56369
rect 6229 56245 6297 56297
rect 6349 56245 6421 56297
rect 6473 56245 6545 56297
rect 6597 56245 6669 56297
rect 6721 56245 6793 56297
rect 6845 56245 6917 56297
rect 6969 56245 7041 56297
rect 7093 56245 7229 56297
rect 6229 56173 7229 56245
rect 6229 56121 6297 56173
rect 6349 56121 6421 56173
rect 6473 56121 6545 56173
rect 6597 56121 6669 56173
rect 6721 56121 6793 56173
rect 6845 56121 6917 56173
rect 6969 56121 7041 56173
rect 7093 56121 7229 56173
rect 6229 56049 7229 56121
rect 6229 55997 6297 56049
rect 6349 55997 6421 56049
rect 6473 55997 6545 56049
rect 6597 55997 6669 56049
rect 6721 55997 6793 56049
rect 6845 55997 6917 56049
rect 6969 55997 7041 56049
rect 7093 55997 7229 56049
rect 6229 55925 7229 55997
rect 6229 55873 6297 55925
rect 6349 55873 6421 55925
rect 6473 55873 6545 55925
rect 6597 55873 6669 55925
rect 6721 55873 6793 55925
rect 6845 55873 6917 55925
rect 6969 55873 7041 55925
rect 7093 55873 7229 55925
rect 6229 55801 7229 55873
rect 6229 55749 6297 55801
rect 6349 55749 6421 55801
rect 6473 55749 6545 55801
rect 6597 55749 6669 55801
rect 6721 55749 6793 55801
rect 6845 55749 6917 55801
rect 6969 55749 7041 55801
rect 7093 55749 7229 55801
rect 6229 55677 7229 55749
rect 6229 55625 6297 55677
rect 6349 55625 6421 55677
rect 6473 55625 6545 55677
rect 6597 55625 6669 55677
rect 6721 55625 6793 55677
rect 6845 55625 6917 55677
rect 6969 55625 7041 55677
rect 7093 55625 7229 55677
rect 6229 55553 7229 55625
rect 6229 55501 6297 55553
rect 6349 55501 6421 55553
rect 6473 55501 6545 55553
rect 6597 55501 6669 55553
rect 6721 55501 6793 55553
rect 6845 55501 6917 55553
rect 6969 55501 7041 55553
rect 7093 55501 7229 55553
rect 6229 55429 7229 55501
rect 6229 55377 6297 55429
rect 6349 55377 6421 55429
rect 6473 55377 6545 55429
rect 6597 55377 6669 55429
rect 6721 55377 6793 55429
rect 6845 55377 6917 55429
rect 6969 55377 7041 55429
rect 7093 55377 7229 55429
rect 6229 55305 7229 55377
rect 6229 55253 6297 55305
rect 6349 55253 6421 55305
rect 6473 55253 6545 55305
rect 6597 55253 6669 55305
rect 6721 55253 6793 55305
rect 6845 55253 6917 55305
rect 6969 55253 7041 55305
rect 7093 55253 7229 55305
rect 6229 55181 7229 55253
rect 6229 55129 6297 55181
rect 6349 55129 6421 55181
rect 6473 55129 6545 55181
rect 6597 55129 6669 55181
rect 6721 55129 6793 55181
rect 6845 55129 6917 55181
rect 6969 55129 7041 55181
rect 7093 55129 7229 55181
rect 6229 55057 7229 55129
rect 6229 55005 6297 55057
rect 6349 55005 6421 55057
rect 6473 55005 6545 55057
rect 6597 55005 6669 55057
rect 6721 55005 6793 55057
rect 6845 55005 6917 55057
rect 6969 55005 7041 55057
rect 7093 55005 7229 55057
rect 6229 54933 7229 55005
rect 6229 54881 6297 54933
rect 6349 54881 6421 54933
rect 6473 54881 6545 54933
rect 6597 54881 6669 54933
rect 6721 54881 6793 54933
rect 6845 54881 6917 54933
rect 6969 54881 7041 54933
rect 7093 54881 7229 54933
rect 6229 54809 7229 54881
rect 6229 54757 6297 54809
rect 6349 54757 6421 54809
rect 6473 54757 6545 54809
rect 6597 54757 6669 54809
rect 6721 54757 6793 54809
rect 6845 54757 6917 54809
rect 6969 54757 7041 54809
rect 7093 54757 7229 54809
rect 6229 54685 7229 54757
rect 6229 54633 6297 54685
rect 6349 54633 6421 54685
rect 6473 54633 6545 54685
rect 6597 54633 6669 54685
rect 6721 54633 6793 54685
rect 6845 54633 6917 54685
rect 6969 54633 7041 54685
rect 7093 54633 7229 54685
rect 6229 54561 7229 54633
rect 6229 54509 6297 54561
rect 6349 54509 6421 54561
rect 6473 54509 6545 54561
rect 6597 54509 6669 54561
rect 6721 54509 6793 54561
rect 6845 54509 6917 54561
rect 6969 54509 7041 54561
rect 7093 54509 7229 54561
rect 6229 54437 7229 54509
rect 6229 54385 6297 54437
rect 6349 54385 6421 54437
rect 6473 54385 6545 54437
rect 6597 54385 6669 54437
rect 6721 54385 6793 54437
rect 6845 54385 6917 54437
rect 6969 54385 7041 54437
rect 7093 54385 7229 54437
rect 6229 54313 7229 54385
rect 6229 54261 6297 54313
rect 6349 54261 6421 54313
rect 6473 54261 6545 54313
rect 6597 54261 6669 54313
rect 6721 54261 6793 54313
rect 6845 54261 6917 54313
rect 6969 54261 7041 54313
rect 7093 54261 7229 54313
rect 6229 54189 7229 54261
rect 6229 54137 6297 54189
rect 6349 54137 6421 54189
rect 6473 54137 6545 54189
rect 6597 54137 6669 54189
rect 6721 54137 6793 54189
rect 6845 54137 6917 54189
rect 6969 54137 7041 54189
rect 7093 54137 7229 54189
rect 6229 54065 7229 54137
rect 6229 54013 6297 54065
rect 6349 54013 6421 54065
rect 6473 54013 6545 54065
rect 6597 54013 6669 54065
rect 6721 54013 6793 54065
rect 6845 54013 6917 54065
rect 6969 54013 7041 54065
rect 7093 54013 7229 54065
rect 6229 53941 7229 54013
rect 6229 53889 6297 53941
rect 6349 53889 6421 53941
rect 6473 53889 6545 53941
rect 6597 53889 6669 53941
rect 6721 53889 6793 53941
rect 6845 53889 6917 53941
rect 6969 53889 7041 53941
rect 7093 53889 7229 53941
rect 6229 53817 7229 53889
rect 6229 53765 6297 53817
rect 6349 53765 6421 53817
rect 6473 53765 6545 53817
rect 6597 53765 6669 53817
rect 6721 53765 6793 53817
rect 6845 53765 6917 53817
rect 6969 53765 7041 53817
rect 7093 53765 7229 53817
rect 6229 53693 7229 53765
rect 6229 53641 6297 53693
rect 6349 53641 6421 53693
rect 6473 53641 6545 53693
rect 6597 53641 6669 53693
rect 6721 53641 6793 53693
rect 6845 53641 6917 53693
rect 6969 53641 7041 53693
rect 7093 53641 7229 53693
rect 6229 53633 7229 53641
rect 4313 53622 7229 53633
rect 4313 53576 4324 53622
rect 7218 53576 7229 53622
rect 4313 53565 7229 53576
rect 7289 56618 7689 56655
rect 7289 53692 7300 56618
rect 7346 53692 7632 56618
rect 7678 53692 7689 56618
rect 7289 53505 7689 53692
rect 7749 56617 7885 56669
rect 7937 56617 8009 56669
rect 8061 56617 8133 56669
rect 8185 56617 8257 56669
rect 8309 56617 8381 56669
rect 8433 56617 8505 56669
rect 8557 56617 8629 56669
rect 8681 56617 8749 56669
rect 7749 56545 8749 56617
rect 7749 56493 7885 56545
rect 7937 56493 8009 56545
rect 8061 56493 8133 56545
rect 8185 56493 8257 56545
rect 8309 56493 8381 56545
rect 8433 56493 8505 56545
rect 8557 56493 8629 56545
rect 8681 56493 8749 56545
rect 7749 56421 8749 56493
rect 7749 56369 7885 56421
rect 7937 56369 8009 56421
rect 8061 56369 8133 56421
rect 8185 56369 8257 56421
rect 8309 56369 8381 56421
rect 8433 56369 8505 56421
rect 8557 56369 8629 56421
rect 8681 56369 8749 56421
rect 7749 56297 8749 56369
rect 7749 56245 7885 56297
rect 7937 56245 8009 56297
rect 8061 56245 8133 56297
rect 8185 56245 8257 56297
rect 8309 56245 8381 56297
rect 8433 56245 8505 56297
rect 8557 56245 8629 56297
rect 8681 56245 8749 56297
rect 7749 56173 8749 56245
rect 7749 56121 7885 56173
rect 7937 56121 8009 56173
rect 8061 56121 8133 56173
rect 8185 56121 8257 56173
rect 8309 56121 8381 56173
rect 8433 56121 8505 56173
rect 8557 56121 8629 56173
rect 8681 56121 8749 56173
rect 7749 56049 8749 56121
rect 7749 55997 7885 56049
rect 7937 55997 8009 56049
rect 8061 55997 8133 56049
rect 8185 55997 8257 56049
rect 8309 55997 8381 56049
rect 8433 55997 8505 56049
rect 8557 55997 8629 56049
rect 8681 55997 8749 56049
rect 7749 55925 8749 55997
rect 7749 55873 7885 55925
rect 7937 55873 8009 55925
rect 8061 55873 8133 55925
rect 8185 55873 8257 55925
rect 8309 55873 8381 55925
rect 8433 55873 8505 55925
rect 8557 55873 8629 55925
rect 8681 55873 8749 55925
rect 7749 55801 8749 55873
rect 7749 55749 7885 55801
rect 7937 55749 8009 55801
rect 8061 55749 8133 55801
rect 8185 55749 8257 55801
rect 8309 55749 8381 55801
rect 8433 55749 8505 55801
rect 8557 55749 8629 55801
rect 8681 55749 8749 55801
rect 7749 55677 8749 55749
rect 7749 55625 7885 55677
rect 7937 55625 8009 55677
rect 8061 55625 8133 55677
rect 8185 55625 8257 55677
rect 8309 55625 8381 55677
rect 8433 55625 8505 55677
rect 8557 55625 8629 55677
rect 8681 55625 8749 55677
rect 7749 55553 8749 55625
rect 7749 55501 7885 55553
rect 7937 55501 8009 55553
rect 8061 55501 8133 55553
rect 8185 55501 8257 55553
rect 8309 55501 8381 55553
rect 8433 55501 8505 55553
rect 8557 55501 8629 55553
rect 8681 55501 8749 55553
rect 7749 55429 8749 55501
rect 7749 55377 7885 55429
rect 7937 55377 8009 55429
rect 8061 55377 8133 55429
rect 8185 55377 8257 55429
rect 8309 55377 8381 55429
rect 8433 55377 8505 55429
rect 8557 55377 8629 55429
rect 8681 55377 8749 55429
rect 7749 55305 8749 55377
rect 7749 55253 7885 55305
rect 7937 55253 8009 55305
rect 8061 55253 8133 55305
rect 8185 55253 8257 55305
rect 8309 55253 8381 55305
rect 8433 55253 8505 55305
rect 8557 55253 8629 55305
rect 8681 55253 8749 55305
rect 7749 55181 8749 55253
rect 7749 55129 7885 55181
rect 7937 55129 8009 55181
rect 8061 55129 8133 55181
rect 8185 55129 8257 55181
rect 8309 55129 8381 55181
rect 8433 55129 8505 55181
rect 8557 55129 8629 55181
rect 8681 55129 8749 55181
rect 7749 55057 8749 55129
rect 7749 55005 7885 55057
rect 7937 55005 8009 55057
rect 8061 55005 8133 55057
rect 8185 55005 8257 55057
rect 8309 55005 8381 55057
rect 8433 55005 8505 55057
rect 8557 55005 8629 55057
rect 8681 55005 8749 55057
rect 7749 54933 8749 55005
rect 7749 54881 7885 54933
rect 7937 54881 8009 54933
rect 8061 54881 8133 54933
rect 8185 54881 8257 54933
rect 8309 54881 8381 54933
rect 8433 54881 8505 54933
rect 8557 54881 8629 54933
rect 8681 54881 8749 54933
rect 7749 54809 8749 54881
rect 7749 54757 7885 54809
rect 7937 54757 8009 54809
rect 8061 54757 8133 54809
rect 8185 54757 8257 54809
rect 8309 54757 8381 54809
rect 8433 54757 8505 54809
rect 8557 54757 8629 54809
rect 8681 54757 8749 54809
rect 7749 54685 8749 54757
rect 7749 54633 7885 54685
rect 7937 54633 8009 54685
rect 8061 54633 8133 54685
rect 8185 54633 8257 54685
rect 8309 54633 8381 54685
rect 8433 54633 8505 54685
rect 8557 54633 8629 54685
rect 8681 54633 8749 54685
rect 7749 54561 8749 54633
rect 7749 54509 7885 54561
rect 7937 54509 8009 54561
rect 8061 54509 8133 54561
rect 8185 54509 8257 54561
rect 8309 54509 8381 54561
rect 8433 54509 8505 54561
rect 8557 54509 8629 54561
rect 8681 54509 8749 54561
rect 7749 54437 8749 54509
rect 7749 54385 7885 54437
rect 7937 54385 8009 54437
rect 8061 54385 8133 54437
rect 8185 54385 8257 54437
rect 8309 54385 8381 54437
rect 8433 54385 8505 54437
rect 8557 54385 8629 54437
rect 8681 54385 8749 54437
rect 7749 54313 8749 54385
rect 7749 54261 7885 54313
rect 7937 54261 8009 54313
rect 8061 54261 8133 54313
rect 8185 54261 8257 54313
rect 8309 54261 8381 54313
rect 8433 54261 8505 54313
rect 8557 54261 8629 54313
rect 8681 54261 8749 54313
rect 7749 54189 8749 54261
rect 7749 54137 7885 54189
rect 7937 54137 8009 54189
rect 8061 54137 8133 54189
rect 8185 54137 8257 54189
rect 8309 54137 8381 54189
rect 8433 54137 8505 54189
rect 8557 54137 8629 54189
rect 8681 54137 8749 54189
rect 7749 54065 8749 54137
rect 7749 54013 7885 54065
rect 7937 54013 8009 54065
rect 8061 54013 8133 54065
rect 8185 54013 8257 54065
rect 8309 54013 8381 54065
rect 8433 54013 8505 54065
rect 8557 54013 8629 54065
rect 8681 54013 8749 54065
rect 7749 53941 8749 54013
rect 7749 53889 7885 53941
rect 7937 53889 8009 53941
rect 8061 53889 8133 53941
rect 8185 53889 8257 53941
rect 8309 53889 8381 53941
rect 8433 53889 8505 53941
rect 8557 53889 8629 53941
rect 8681 53889 8749 53941
rect 7749 53817 8749 53889
rect 7749 53765 7885 53817
rect 7937 53765 8009 53817
rect 8061 53765 8133 53817
rect 8185 53765 8257 53817
rect 8309 53765 8381 53817
rect 8433 53765 8505 53817
rect 8557 53765 8629 53817
rect 8681 53765 8749 53817
rect 7749 53693 8749 53765
rect 7749 53641 7885 53693
rect 7937 53641 8009 53693
rect 8061 53641 8133 53693
rect 8185 53641 8257 53693
rect 8309 53641 8381 53693
rect 8433 53641 8505 53693
rect 8557 53641 8629 53693
rect 8681 53641 8749 53693
rect 7749 53633 8749 53641
rect 9665 56669 10665 56677
rect 9665 56617 10214 56669
rect 10266 56617 10338 56669
rect 10390 56617 10462 56669
rect 10514 56617 10586 56669
rect 10638 56617 10665 56669
rect 11185 56734 14101 56745
rect 11185 56688 11196 56734
rect 14090 56688 14101 56734
rect 11185 56677 14101 56688
rect 11185 56669 12185 56677
rect 9665 56545 10665 56617
rect 9665 56493 10214 56545
rect 10266 56493 10338 56545
rect 10390 56493 10462 56545
rect 10514 56493 10586 56545
rect 10638 56493 10665 56545
rect 9665 56421 10665 56493
rect 9665 56369 10214 56421
rect 10266 56369 10338 56421
rect 10390 56369 10462 56421
rect 10514 56369 10586 56421
rect 10638 56369 10665 56421
rect 9665 56297 10665 56369
rect 9665 56245 10214 56297
rect 10266 56245 10338 56297
rect 10390 56245 10462 56297
rect 10514 56245 10586 56297
rect 10638 56245 10665 56297
rect 9665 56173 10665 56245
rect 9665 56121 10214 56173
rect 10266 56121 10338 56173
rect 10390 56121 10462 56173
rect 10514 56121 10586 56173
rect 10638 56121 10665 56173
rect 9665 56049 10665 56121
rect 9665 55997 10214 56049
rect 10266 55997 10338 56049
rect 10390 55997 10462 56049
rect 10514 55997 10586 56049
rect 10638 55997 10665 56049
rect 9665 55925 10665 55997
rect 9665 55873 10214 55925
rect 10266 55873 10338 55925
rect 10390 55873 10462 55925
rect 10514 55873 10586 55925
rect 10638 55873 10665 55925
rect 9665 55801 10665 55873
rect 9665 55749 10214 55801
rect 10266 55749 10338 55801
rect 10390 55749 10462 55801
rect 10514 55749 10586 55801
rect 10638 55749 10665 55801
rect 9665 55677 10665 55749
rect 9665 55625 10214 55677
rect 10266 55625 10338 55677
rect 10390 55625 10462 55677
rect 10514 55625 10586 55677
rect 10638 55625 10665 55677
rect 9665 55553 10665 55625
rect 9665 55501 10214 55553
rect 10266 55501 10338 55553
rect 10390 55501 10462 55553
rect 10514 55501 10586 55553
rect 10638 55501 10665 55553
rect 9665 55429 10665 55501
rect 9665 55377 10214 55429
rect 10266 55377 10338 55429
rect 10390 55377 10462 55429
rect 10514 55377 10586 55429
rect 10638 55377 10665 55429
rect 9665 55305 10665 55377
rect 9665 55253 10214 55305
rect 10266 55253 10338 55305
rect 10390 55253 10462 55305
rect 10514 55253 10586 55305
rect 10638 55253 10665 55305
rect 9665 55181 10665 55253
rect 9665 55129 10214 55181
rect 10266 55129 10338 55181
rect 10390 55129 10462 55181
rect 10514 55129 10586 55181
rect 10638 55129 10665 55181
rect 9665 55057 10665 55129
rect 9665 55005 10214 55057
rect 10266 55005 10338 55057
rect 10390 55005 10462 55057
rect 10514 55005 10586 55057
rect 10638 55005 10665 55057
rect 9665 54933 10665 55005
rect 9665 54881 10214 54933
rect 10266 54881 10338 54933
rect 10390 54881 10462 54933
rect 10514 54881 10586 54933
rect 10638 54881 10665 54933
rect 9665 54809 10665 54881
rect 9665 54757 10214 54809
rect 10266 54757 10338 54809
rect 10390 54757 10462 54809
rect 10514 54757 10586 54809
rect 10638 54757 10665 54809
rect 9665 54685 10665 54757
rect 9665 54633 10214 54685
rect 10266 54633 10338 54685
rect 10390 54633 10462 54685
rect 10514 54633 10586 54685
rect 10638 54633 10665 54685
rect 9665 54561 10665 54633
rect 9665 54509 10214 54561
rect 10266 54509 10338 54561
rect 10390 54509 10462 54561
rect 10514 54509 10586 54561
rect 10638 54509 10665 54561
rect 9665 54437 10665 54509
rect 9665 54385 10214 54437
rect 10266 54385 10338 54437
rect 10390 54385 10462 54437
rect 10514 54385 10586 54437
rect 10638 54385 10665 54437
rect 9665 54313 10665 54385
rect 9665 54261 10214 54313
rect 10266 54261 10338 54313
rect 10390 54261 10462 54313
rect 10514 54261 10586 54313
rect 10638 54261 10665 54313
rect 9665 54189 10665 54261
rect 9665 54137 10214 54189
rect 10266 54137 10338 54189
rect 10390 54137 10462 54189
rect 10514 54137 10586 54189
rect 10638 54137 10665 54189
rect 9665 54065 10665 54137
rect 9665 54013 10214 54065
rect 10266 54013 10338 54065
rect 10390 54013 10462 54065
rect 10514 54013 10586 54065
rect 10638 54013 10665 54065
rect 9665 53941 10665 54013
rect 9665 53889 10214 53941
rect 10266 53889 10338 53941
rect 10390 53889 10462 53941
rect 10514 53889 10586 53941
rect 10638 53889 10665 53941
rect 9665 53817 10665 53889
rect 9665 53765 10214 53817
rect 10266 53765 10338 53817
rect 10390 53765 10462 53817
rect 10514 53765 10586 53817
rect 10638 53765 10665 53817
rect 9665 53693 10665 53765
rect 9665 53641 10214 53693
rect 10266 53641 10338 53693
rect 10390 53641 10462 53693
rect 10514 53641 10586 53693
rect 10638 53641 10665 53693
rect 9665 53633 10665 53641
rect 7749 53622 10665 53633
rect 7749 53576 7760 53622
rect 10654 53576 10665 53622
rect 7749 53565 10665 53576
rect 10725 56618 11125 56655
rect 10725 53692 10736 56618
rect 10782 53692 11068 56618
rect 11114 53692 11125 56618
rect 10725 53505 11125 53692
rect 11185 56617 11225 56669
rect 11277 56617 11349 56669
rect 11401 56617 11473 56669
rect 11525 56617 11597 56669
rect 11649 56617 11721 56669
rect 11773 56617 11845 56669
rect 11897 56617 11969 56669
rect 12021 56617 12093 56669
rect 12145 56617 12185 56669
rect 11185 56545 12185 56617
rect 11185 56493 11225 56545
rect 11277 56493 11349 56545
rect 11401 56493 11473 56545
rect 11525 56493 11597 56545
rect 11649 56493 11721 56545
rect 11773 56493 11845 56545
rect 11897 56493 11969 56545
rect 12021 56493 12093 56545
rect 12145 56493 12185 56545
rect 11185 56421 12185 56493
rect 11185 56369 11225 56421
rect 11277 56369 11349 56421
rect 11401 56369 11473 56421
rect 11525 56369 11597 56421
rect 11649 56369 11721 56421
rect 11773 56369 11845 56421
rect 11897 56369 11969 56421
rect 12021 56369 12093 56421
rect 12145 56369 12185 56421
rect 11185 56297 12185 56369
rect 11185 56245 11225 56297
rect 11277 56245 11349 56297
rect 11401 56245 11473 56297
rect 11525 56245 11597 56297
rect 11649 56245 11721 56297
rect 11773 56245 11845 56297
rect 11897 56245 11969 56297
rect 12021 56245 12093 56297
rect 12145 56245 12185 56297
rect 11185 56173 12185 56245
rect 11185 56121 11225 56173
rect 11277 56121 11349 56173
rect 11401 56121 11473 56173
rect 11525 56121 11597 56173
rect 11649 56121 11721 56173
rect 11773 56121 11845 56173
rect 11897 56121 11969 56173
rect 12021 56121 12093 56173
rect 12145 56121 12185 56173
rect 11185 56049 12185 56121
rect 11185 55997 11225 56049
rect 11277 55997 11349 56049
rect 11401 55997 11473 56049
rect 11525 55997 11597 56049
rect 11649 55997 11721 56049
rect 11773 55997 11845 56049
rect 11897 55997 11969 56049
rect 12021 55997 12093 56049
rect 12145 55997 12185 56049
rect 11185 55925 12185 55997
rect 11185 55873 11225 55925
rect 11277 55873 11349 55925
rect 11401 55873 11473 55925
rect 11525 55873 11597 55925
rect 11649 55873 11721 55925
rect 11773 55873 11845 55925
rect 11897 55873 11969 55925
rect 12021 55873 12093 55925
rect 12145 55873 12185 55925
rect 11185 55801 12185 55873
rect 11185 55749 11225 55801
rect 11277 55749 11349 55801
rect 11401 55749 11473 55801
rect 11525 55749 11597 55801
rect 11649 55749 11721 55801
rect 11773 55749 11845 55801
rect 11897 55749 11969 55801
rect 12021 55749 12093 55801
rect 12145 55749 12185 55801
rect 11185 55677 12185 55749
rect 11185 55625 11225 55677
rect 11277 55625 11349 55677
rect 11401 55625 11473 55677
rect 11525 55625 11597 55677
rect 11649 55625 11721 55677
rect 11773 55625 11845 55677
rect 11897 55625 11969 55677
rect 12021 55625 12093 55677
rect 12145 55625 12185 55677
rect 11185 55553 12185 55625
rect 11185 55501 11225 55553
rect 11277 55501 11349 55553
rect 11401 55501 11473 55553
rect 11525 55501 11597 55553
rect 11649 55501 11721 55553
rect 11773 55501 11845 55553
rect 11897 55501 11969 55553
rect 12021 55501 12093 55553
rect 12145 55501 12185 55553
rect 11185 55429 12185 55501
rect 11185 55377 11225 55429
rect 11277 55377 11349 55429
rect 11401 55377 11473 55429
rect 11525 55377 11597 55429
rect 11649 55377 11721 55429
rect 11773 55377 11845 55429
rect 11897 55377 11969 55429
rect 12021 55377 12093 55429
rect 12145 55377 12185 55429
rect 11185 55305 12185 55377
rect 11185 55253 11225 55305
rect 11277 55253 11349 55305
rect 11401 55253 11473 55305
rect 11525 55253 11597 55305
rect 11649 55253 11721 55305
rect 11773 55253 11845 55305
rect 11897 55253 11969 55305
rect 12021 55253 12093 55305
rect 12145 55253 12185 55305
rect 11185 55181 12185 55253
rect 11185 55129 11225 55181
rect 11277 55129 11349 55181
rect 11401 55129 11473 55181
rect 11525 55129 11597 55181
rect 11649 55129 11721 55181
rect 11773 55129 11845 55181
rect 11897 55129 11969 55181
rect 12021 55129 12093 55181
rect 12145 55129 12185 55181
rect 11185 55057 12185 55129
rect 11185 55005 11225 55057
rect 11277 55005 11349 55057
rect 11401 55005 11473 55057
rect 11525 55005 11597 55057
rect 11649 55005 11721 55057
rect 11773 55005 11845 55057
rect 11897 55005 11969 55057
rect 12021 55005 12093 55057
rect 12145 55005 12185 55057
rect 11185 54933 12185 55005
rect 11185 54881 11225 54933
rect 11277 54881 11349 54933
rect 11401 54881 11473 54933
rect 11525 54881 11597 54933
rect 11649 54881 11721 54933
rect 11773 54881 11845 54933
rect 11897 54881 11969 54933
rect 12021 54881 12093 54933
rect 12145 54881 12185 54933
rect 11185 54809 12185 54881
rect 11185 54757 11225 54809
rect 11277 54757 11349 54809
rect 11401 54757 11473 54809
rect 11525 54757 11597 54809
rect 11649 54757 11721 54809
rect 11773 54757 11845 54809
rect 11897 54757 11969 54809
rect 12021 54757 12093 54809
rect 12145 54757 12185 54809
rect 11185 54685 12185 54757
rect 11185 54633 11225 54685
rect 11277 54633 11349 54685
rect 11401 54633 11473 54685
rect 11525 54633 11597 54685
rect 11649 54633 11721 54685
rect 11773 54633 11845 54685
rect 11897 54633 11969 54685
rect 12021 54633 12093 54685
rect 12145 54633 12185 54685
rect 11185 54561 12185 54633
rect 11185 54509 11225 54561
rect 11277 54509 11349 54561
rect 11401 54509 11473 54561
rect 11525 54509 11597 54561
rect 11649 54509 11721 54561
rect 11773 54509 11845 54561
rect 11897 54509 11969 54561
rect 12021 54509 12093 54561
rect 12145 54509 12185 54561
rect 11185 54437 12185 54509
rect 11185 54385 11225 54437
rect 11277 54385 11349 54437
rect 11401 54385 11473 54437
rect 11525 54385 11597 54437
rect 11649 54385 11721 54437
rect 11773 54385 11845 54437
rect 11897 54385 11969 54437
rect 12021 54385 12093 54437
rect 12145 54385 12185 54437
rect 11185 54313 12185 54385
rect 11185 54261 11225 54313
rect 11277 54261 11349 54313
rect 11401 54261 11473 54313
rect 11525 54261 11597 54313
rect 11649 54261 11721 54313
rect 11773 54261 11845 54313
rect 11897 54261 11969 54313
rect 12021 54261 12093 54313
rect 12145 54261 12185 54313
rect 11185 54189 12185 54261
rect 11185 54137 11225 54189
rect 11277 54137 11349 54189
rect 11401 54137 11473 54189
rect 11525 54137 11597 54189
rect 11649 54137 11721 54189
rect 11773 54137 11845 54189
rect 11897 54137 11969 54189
rect 12021 54137 12093 54189
rect 12145 54137 12185 54189
rect 11185 54065 12185 54137
rect 11185 54013 11225 54065
rect 11277 54013 11349 54065
rect 11401 54013 11473 54065
rect 11525 54013 11597 54065
rect 11649 54013 11721 54065
rect 11773 54013 11845 54065
rect 11897 54013 11969 54065
rect 12021 54013 12093 54065
rect 12145 54013 12185 54065
rect 11185 53941 12185 54013
rect 11185 53889 11225 53941
rect 11277 53889 11349 53941
rect 11401 53889 11473 53941
rect 11525 53889 11597 53941
rect 11649 53889 11721 53941
rect 11773 53889 11845 53941
rect 11897 53889 11969 53941
rect 12021 53889 12093 53941
rect 12145 53889 12185 53941
rect 11185 53817 12185 53889
rect 11185 53765 11225 53817
rect 11277 53765 11349 53817
rect 11401 53765 11473 53817
rect 11525 53765 11597 53817
rect 11649 53765 11721 53817
rect 11773 53765 11845 53817
rect 11897 53765 11969 53817
rect 12021 53765 12093 53817
rect 12145 53765 12185 53817
rect 11185 53693 12185 53765
rect 11185 53641 11225 53693
rect 11277 53641 11349 53693
rect 11401 53641 11473 53693
rect 11525 53641 11597 53693
rect 11649 53641 11721 53693
rect 11773 53641 11845 53693
rect 11897 53641 11969 53693
rect 12021 53641 12093 53693
rect 12145 53641 12185 53693
rect 11185 53633 12185 53641
rect 13101 56669 14101 56677
rect 13101 56617 13141 56669
rect 13193 56617 13265 56669
rect 13317 56617 13389 56669
rect 13441 56617 13513 56669
rect 13565 56617 13637 56669
rect 13689 56617 13761 56669
rect 13813 56617 13885 56669
rect 13937 56617 14009 56669
rect 14061 56617 14101 56669
rect 14565 56655 14576 57048
rect 13101 56545 14101 56617
rect 13101 56493 13141 56545
rect 13193 56493 13265 56545
rect 13317 56493 13389 56545
rect 13441 56493 13513 56545
rect 13565 56493 13637 56545
rect 13689 56493 13761 56545
rect 13813 56493 13885 56545
rect 13937 56493 14009 56545
rect 14061 56493 14101 56545
rect 13101 56421 14101 56493
rect 13101 56369 13141 56421
rect 13193 56369 13265 56421
rect 13317 56369 13389 56421
rect 13441 56369 13513 56421
rect 13565 56369 13637 56421
rect 13689 56369 13761 56421
rect 13813 56369 13885 56421
rect 13937 56369 14009 56421
rect 14061 56369 14101 56421
rect 13101 56297 14101 56369
rect 13101 56245 13141 56297
rect 13193 56245 13265 56297
rect 13317 56245 13389 56297
rect 13441 56245 13513 56297
rect 13565 56245 13637 56297
rect 13689 56245 13761 56297
rect 13813 56245 13885 56297
rect 13937 56245 14009 56297
rect 14061 56245 14101 56297
rect 13101 56173 14101 56245
rect 13101 56121 13141 56173
rect 13193 56121 13265 56173
rect 13317 56121 13389 56173
rect 13441 56121 13513 56173
rect 13565 56121 13637 56173
rect 13689 56121 13761 56173
rect 13813 56121 13885 56173
rect 13937 56121 14009 56173
rect 14061 56121 14101 56173
rect 13101 56049 14101 56121
rect 13101 55997 13141 56049
rect 13193 55997 13265 56049
rect 13317 55997 13389 56049
rect 13441 55997 13513 56049
rect 13565 55997 13637 56049
rect 13689 55997 13761 56049
rect 13813 55997 13885 56049
rect 13937 55997 14009 56049
rect 14061 55997 14101 56049
rect 13101 55925 14101 55997
rect 13101 55873 13141 55925
rect 13193 55873 13265 55925
rect 13317 55873 13389 55925
rect 13441 55873 13513 55925
rect 13565 55873 13637 55925
rect 13689 55873 13761 55925
rect 13813 55873 13885 55925
rect 13937 55873 14009 55925
rect 14061 55873 14101 55925
rect 13101 55801 14101 55873
rect 13101 55749 13141 55801
rect 13193 55749 13265 55801
rect 13317 55749 13389 55801
rect 13441 55749 13513 55801
rect 13565 55749 13637 55801
rect 13689 55749 13761 55801
rect 13813 55749 13885 55801
rect 13937 55749 14009 55801
rect 14061 55749 14101 55801
rect 13101 55677 14101 55749
rect 13101 55625 13141 55677
rect 13193 55625 13265 55677
rect 13317 55625 13389 55677
rect 13441 55625 13513 55677
rect 13565 55625 13637 55677
rect 13689 55625 13761 55677
rect 13813 55625 13885 55677
rect 13937 55625 14009 55677
rect 14061 55625 14101 55677
rect 13101 55553 14101 55625
rect 13101 55501 13141 55553
rect 13193 55501 13265 55553
rect 13317 55501 13389 55553
rect 13441 55501 13513 55553
rect 13565 55501 13637 55553
rect 13689 55501 13761 55553
rect 13813 55501 13885 55553
rect 13937 55501 14009 55553
rect 14061 55501 14101 55553
rect 13101 55429 14101 55501
rect 13101 55377 13141 55429
rect 13193 55377 13265 55429
rect 13317 55377 13389 55429
rect 13441 55377 13513 55429
rect 13565 55377 13637 55429
rect 13689 55377 13761 55429
rect 13813 55377 13885 55429
rect 13937 55377 14009 55429
rect 14061 55377 14101 55429
rect 13101 55305 14101 55377
rect 13101 55253 13141 55305
rect 13193 55253 13265 55305
rect 13317 55253 13389 55305
rect 13441 55253 13513 55305
rect 13565 55253 13637 55305
rect 13689 55253 13761 55305
rect 13813 55253 13885 55305
rect 13937 55253 14009 55305
rect 14061 55253 14101 55305
rect 13101 55181 14101 55253
rect 13101 55129 13141 55181
rect 13193 55129 13265 55181
rect 13317 55129 13389 55181
rect 13441 55129 13513 55181
rect 13565 55129 13637 55181
rect 13689 55129 13761 55181
rect 13813 55129 13885 55181
rect 13937 55129 14009 55181
rect 14061 55129 14101 55181
rect 13101 55057 14101 55129
rect 13101 55005 13141 55057
rect 13193 55005 13265 55057
rect 13317 55005 13389 55057
rect 13441 55005 13513 55057
rect 13565 55005 13637 55057
rect 13689 55005 13761 55057
rect 13813 55005 13885 55057
rect 13937 55005 14009 55057
rect 14061 55005 14101 55057
rect 13101 54933 14101 55005
rect 13101 54881 13141 54933
rect 13193 54881 13265 54933
rect 13317 54881 13389 54933
rect 13441 54881 13513 54933
rect 13565 54881 13637 54933
rect 13689 54881 13761 54933
rect 13813 54881 13885 54933
rect 13937 54881 14009 54933
rect 14061 54881 14101 54933
rect 13101 54809 14101 54881
rect 13101 54757 13141 54809
rect 13193 54757 13265 54809
rect 13317 54757 13389 54809
rect 13441 54757 13513 54809
rect 13565 54757 13637 54809
rect 13689 54757 13761 54809
rect 13813 54757 13885 54809
rect 13937 54757 14009 54809
rect 14061 54757 14101 54809
rect 13101 54685 14101 54757
rect 13101 54633 13141 54685
rect 13193 54633 13265 54685
rect 13317 54633 13389 54685
rect 13441 54633 13513 54685
rect 13565 54633 13637 54685
rect 13689 54633 13761 54685
rect 13813 54633 13885 54685
rect 13937 54633 14009 54685
rect 14061 54633 14101 54685
rect 13101 54561 14101 54633
rect 13101 54509 13141 54561
rect 13193 54509 13265 54561
rect 13317 54509 13389 54561
rect 13441 54509 13513 54561
rect 13565 54509 13637 54561
rect 13689 54509 13761 54561
rect 13813 54509 13885 54561
rect 13937 54509 14009 54561
rect 14061 54509 14101 54561
rect 13101 54437 14101 54509
rect 13101 54385 13141 54437
rect 13193 54385 13265 54437
rect 13317 54385 13389 54437
rect 13441 54385 13513 54437
rect 13565 54385 13637 54437
rect 13689 54385 13761 54437
rect 13813 54385 13885 54437
rect 13937 54385 14009 54437
rect 14061 54385 14101 54437
rect 13101 54313 14101 54385
rect 13101 54261 13141 54313
rect 13193 54261 13265 54313
rect 13317 54261 13389 54313
rect 13441 54261 13513 54313
rect 13565 54261 13637 54313
rect 13689 54261 13761 54313
rect 13813 54261 13885 54313
rect 13937 54261 14009 54313
rect 14061 54261 14101 54313
rect 13101 54189 14101 54261
rect 13101 54137 13141 54189
rect 13193 54137 13265 54189
rect 13317 54137 13389 54189
rect 13441 54137 13513 54189
rect 13565 54137 13637 54189
rect 13689 54137 13761 54189
rect 13813 54137 13885 54189
rect 13937 54137 14009 54189
rect 14061 54137 14101 54189
rect 13101 54065 14101 54137
rect 13101 54013 13141 54065
rect 13193 54013 13265 54065
rect 13317 54013 13389 54065
rect 13441 54013 13513 54065
rect 13565 54013 13637 54065
rect 13689 54013 13761 54065
rect 13813 54013 13885 54065
rect 13937 54013 14009 54065
rect 14061 54013 14101 54065
rect 13101 53941 14101 54013
rect 13101 53889 13141 53941
rect 13193 53889 13265 53941
rect 13317 53889 13389 53941
rect 13441 53889 13513 53941
rect 13565 53889 13637 53941
rect 13689 53889 13761 53941
rect 13813 53889 13885 53941
rect 13937 53889 14009 53941
rect 14061 53889 14101 53941
rect 13101 53817 14101 53889
rect 13101 53765 13141 53817
rect 13193 53765 13265 53817
rect 13317 53765 13389 53817
rect 13441 53765 13513 53817
rect 13565 53765 13637 53817
rect 13689 53765 13761 53817
rect 13813 53765 13885 53817
rect 13937 53765 14009 53817
rect 14061 53765 14101 53817
rect 13101 53693 14101 53765
rect 13101 53641 13141 53693
rect 13193 53641 13265 53693
rect 13317 53641 13389 53693
rect 13441 53641 13513 53693
rect 13565 53641 13637 53693
rect 13689 53641 13761 53693
rect 13813 53641 13885 53693
rect 13937 53641 14009 53693
rect 14061 53641 14101 53693
rect 13101 53633 14101 53641
rect 11185 53622 14101 53633
rect 11185 53576 11196 53622
rect 14090 53576 14101 53622
rect 11185 53565 14101 53576
rect 14161 56618 14576 56655
rect 14161 53692 14172 56618
rect 14218 53692 14576 56618
rect 14161 53505 14576 53692
rect 402 53484 14576 53505
rect 402 53432 2501 53484
rect 2553 53432 2609 53484
rect 2661 53432 4871 53484
rect 4923 53432 4979 53484
rect 5031 53432 7247 53484
rect 7299 53432 7355 53484
rect 7407 53432 7463 53484
rect 7515 53432 7571 53484
rect 7623 53432 7679 53484
rect 7731 53432 9947 53484
rect 9999 53432 10055 53484
rect 10107 53432 12317 53484
rect 12369 53432 12425 53484
rect 12477 53432 14576 53484
rect 402 53376 14576 53432
rect 402 53324 2501 53376
rect 2553 53324 2609 53376
rect 2661 53324 4871 53376
rect 4923 53324 4979 53376
rect 5031 53324 7247 53376
rect 7299 53324 7355 53376
rect 7407 53324 7463 53376
rect 7515 53324 7571 53376
rect 7623 53324 7679 53376
rect 7731 53324 9947 53376
rect 9999 53324 10055 53376
rect 10107 53324 12317 53376
rect 12369 53324 12425 53376
rect 12477 53324 14576 53376
rect 402 53268 14576 53324
rect 402 53251 2501 53268
rect 2553 53251 2609 53268
rect 2661 53251 4871 53268
rect 4923 53251 4979 53268
rect 5031 53251 7247 53268
rect 7299 53251 7355 53268
rect 7407 53251 7463 53268
rect 7515 53251 7571 53268
rect 7623 53251 7679 53268
rect 7731 53251 9947 53268
rect 9999 53251 10055 53268
rect 10107 53251 12317 53268
rect 12369 53251 12425 53268
rect 12477 53251 14576 53268
rect 402 53205 510 53251
rect 14468 53205 14576 53251
rect 14622 53205 14633 57105
rect 345 53194 14633 53205
rect 71 52611 2225 52622
rect 71 52586 268 52611
rect 10 52574 268 52586
rect 10 52522 22 52574
rect 74 52522 268 52574
rect 10 52466 268 52522
rect 10 52414 22 52466
rect 74 52414 268 52466
rect 10 52358 268 52414
rect 10 52306 22 52358
rect 74 52306 268 52358
rect 10 52250 268 52306
rect 10 52198 22 52250
rect 74 52198 268 52250
rect 10 52142 268 52198
rect 10 52090 22 52142
rect 74 52090 268 52142
rect 10 52034 268 52090
rect 10 51982 22 52034
rect 74 51982 268 52034
rect 10 51926 268 51982
rect 10 51874 22 51926
rect 74 51874 268 51926
rect 10 51818 268 51874
rect 10 51766 22 51818
rect 74 51766 268 51818
rect 10 51710 268 51766
rect 10 51658 22 51710
rect 74 51658 268 51710
rect 10 51622 268 51658
rect 10 51602 86 51622
rect 10 51550 22 51602
rect 74 51550 86 51602
rect 10 51494 86 51550
rect 10 51442 22 51494
rect 74 51442 86 51494
rect 10 51422 86 51442
rect 257 51422 268 51622
rect 10 51386 268 51422
rect 10 51334 22 51386
rect 74 51334 268 51386
rect 10 51278 268 51334
rect 10 51226 22 51278
rect 74 51226 268 51278
rect 10 51214 268 51226
rect 71 50422 268 51214
rect 257 49854 268 50422
rect 71 48854 268 49854
rect 257 48654 268 48854
rect 71 47665 268 48654
rect 2214 47665 2225 52611
rect 71 47654 2225 47665
rect 2551 52611 12427 52622
rect 2551 47665 2562 52611
rect 2908 52588 3016 52611
rect 11962 52588 12070 52611
rect 2908 52536 2934 52588
rect 2986 52536 3016 52588
rect 11962 52536 11992 52588
rect 12044 52536 12070 52588
rect 2908 52464 3016 52536
rect 11962 52464 12070 52536
rect 2908 52412 2934 52464
rect 2986 52412 3016 52464
rect 11962 52412 11992 52464
rect 12044 52412 12070 52464
rect 2908 52340 3016 52412
rect 11962 52340 12070 52412
rect 2908 52288 2934 52340
rect 2986 52288 3016 52340
rect 11962 52288 11992 52340
rect 12044 52288 12070 52340
rect 2908 52265 3016 52288
rect 11962 52265 12070 52288
rect 2908 52254 12070 52265
rect 2908 48022 2919 52254
rect 3105 52029 11873 52040
rect 3105 51983 3142 52029
rect 11836 51983 11873 52029
rect 3105 51965 4863 51983
rect 4915 51965 4987 51983
rect 5039 51965 7277 51983
rect 7329 51965 7401 51983
rect 7453 51965 7525 51983
rect 7577 51965 7649 51983
rect 7701 51965 9939 51983
rect 9991 51965 10063 51983
rect 10115 51965 11873 51983
rect 3105 51900 11873 51965
rect 3105 48376 3116 51900
rect 3162 51893 11816 51900
rect 3162 51875 4863 51893
rect 4915 51875 4987 51893
rect 5039 51875 7277 51893
rect 7329 51875 7401 51893
rect 7453 51875 7525 51893
rect 7577 51875 7649 51893
rect 7701 51875 9939 51893
rect 9991 51875 10063 51893
rect 10115 51875 11816 51893
rect 3162 51844 3424 51875
rect 3162 51234 3270 51844
rect 3316 51829 3424 51844
rect 11554 51844 11816 51875
rect 11554 51829 11662 51844
rect 3316 51818 11662 51829
rect 3316 51260 3327 51818
rect 3489 51627 11489 51639
rect 3489 51626 3559 51627
rect 3611 51626 3683 51627
rect 3735 51626 3807 51627
rect 3859 51626 3931 51627
rect 3983 51626 4055 51627
rect 4107 51626 4179 51627
rect 4231 51626 4303 51627
rect 4355 51626 4427 51627
rect 4479 51626 4551 51627
rect 4603 51626 4675 51627
rect 4727 51626 5180 51627
rect 5232 51626 5304 51627
rect 5356 51626 5428 51627
rect 5480 51626 5552 51627
rect 5604 51626 5676 51627
rect 5728 51626 5800 51627
rect 5852 51626 5924 51627
rect 5976 51626 6048 51627
rect 6100 51626 6172 51627
rect 6224 51626 6296 51627
rect 6348 51626 6420 51627
rect 6472 51626 6544 51627
rect 6596 51626 6668 51627
rect 6720 51626 6792 51627
rect 6844 51626 6916 51627
rect 6968 51626 7040 51627
rect 7092 51626 7886 51627
rect 7938 51626 8010 51627
rect 8062 51626 8134 51627
rect 8186 51626 8258 51627
rect 8310 51626 8382 51627
rect 8434 51626 8506 51627
rect 8558 51626 8630 51627
rect 8682 51626 8754 51627
rect 8806 51626 8878 51627
rect 8930 51626 9002 51627
rect 9054 51626 9126 51627
rect 9178 51626 9250 51627
rect 9302 51626 9374 51627
rect 9426 51626 9498 51627
rect 9550 51626 9622 51627
rect 9674 51626 9746 51627
rect 9798 51626 10251 51627
rect 10303 51626 10375 51627
rect 10427 51626 10499 51627
rect 10551 51626 10623 51627
rect 10675 51626 10747 51627
rect 10799 51626 10871 51627
rect 10923 51626 10995 51627
rect 11047 51626 11119 51627
rect 11171 51626 11243 51627
rect 11295 51626 11367 51627
rect 11419 51626 11489 51627
rect 3489 51580 3502 51626
rect 11476 51580 11489 51626
rect 3489 51575 3559 51580
rect 3611 51575 3683 51580
rect 3735 51575 3807 51580
rect 3859 51575 3931 51580
rect 3983 51575 4055 51580
rect 4107 51575 4179 51580
rect 4231 51575 4303 51580
rect 4355 51575 4427 51580
rect 4479 51575 4551 51580
rect 4603 51575 4675 51580
rect 4727 51575 5180 51580
rect 5232 51575 5304 51580
rect 5356 51575 5428 51580
rect 5480 51575 5552 51580
rect 5604 51575 5676 51580
rect 5728 51575 5800 51580
rect 5852 51575 5924 51580
rect 5976 51575 6048 51580
rect 6100 51575 6172 51580
rect 6224 51575 6296 51580
rect 6348 51575 6420 51580
rect 6472 51575 6544 51580
rect 6596 51575 6668 51580
rect 6720 51575 6792 51580
rect 6844 51575 6916 51580
rect 6968 51575 7040 51580
rect 7092 51575 7886 51580
rect 7938 51575 8010 51580
rect 8062 51575 8134 51580
rect 8186 51575 8258 51580
rect 8310 51575 8382 51580
rect 8434 51575 8506 51580
rect 8558 51575 8630 51580
rect 8682 51575 8754 51580
rect 8806 51575 8878 51580
rect 8930 51575 9002 51580
rect 9054 51575 9126 51580
rect 9178 51575 9250 51580
rect 9302 51575 9374 51580
rect 9426 51575 9498 51580
rect 9550 51575 9622 51580
rect 9674 51575 9746 51580
rect 9798 51575 10251 51580
rect 10303 51575 10375 51580
rect 10427 51575 10499 51580
rect 10551 51575 10623 51580
rect 10675 51575 10747 51580
rect 10799 51575 10871 51580
rect 10923 51575 10995 51580
rect 11047 51575 11119 51580
rect 11171 51575 11243 51580
rect 11295 51575 11367 51580
rect 11419 51575 11489 51580
rect 3489 51503 11489 51575
rect 3489 51498 3559 51503
rect 3611 51498 3683 51503
rect 3735 51498 3807 51503
rect 3859 51498 3931 51503
rect 3983 51498 4055 51503
rect 4107 51498 4179 51503
rect 4231 51498 4303 51503
rect 4355 51498 4427 51503
rect 4479 51498 4551 51503
rect 4603 51498 4675 51503
rect 4727 51498 5180 51503
rect 5232 51498 5304 51503
rect 5356 51498 5428 51503
rect 5480 51498 5552 51503
rect 5604 51498 5676 51503
rect 5728 51498 5800 51503
rect 5852 51498 5924 51503
rect 5976 51498 6048 51503
rect 6100 51498 6172 51503
rect 6224 51498 6296 51503
rect 6348 51498 6420 51503
rect 6472 51498 6544 51503
rect 6596 51498 6668 51503
rect 6720 51498 6792 51503
rect 6844 51498 6916 51503
rect 6968 51498 7040 51503
rect 7092 51498 7886 51503
rect 7938 51498 8010 51503
rect 8062 51498 8134 51503
rect 8186 51498 8258 51503
rect 8310 51498 8382 51503
rect 8434 51498 8506 51503
rect 8558 51498 8630 51503
rect 8682 51498 8754 51503
rect 8806 51498 8878 51503
rect 8930 51498 9002 51503
rect 9054 51498 9126 51503
rect 9178 51498 9250 51503
rect 9302 51498 9374 51503
rect 9426 51498 9498 51503
rect 9550 51498 9622 51503
rect 9674 51498 9746 51503
rect 9798 51498 10251 51503
rect 10303 51498 10375 51503
rect 10427 51498 10499 51503
rect 10551 51498 10623 51503
rect 10675 51498 10747 51503
rect 10799 51498 10871 51503
rect 10923 51498 10995 51503
rect 11047 51498 11119 51503
rect 11171 51498 11243 51503
rect 11295 51498 11367 51503
rect 11419 51498 11489 51503
rect 3489 51452 3502 51498
rect 11476 51452 11489 51498
rect 3489 51451 3559 51452
rect 3611 51451 3683 51452
rect 3735 51451 3807 51452
rect 3859 51451 3931 51452
rect 3983 51451 4055 51452
rect 4107 51451 4179 51452
rect 4231 51451 4303 51452
rect 4355 51451 4427 51452
rect 4479 51451 4551 51452
rect 4603 51451 4675 51452
rect 4727 51451 5180 51452
rect 5232 51451 5304 51452
rect 5356 51451 5428 51452
rect 5480 51451 5552 51452
rect 5604 51451 5676 51452
rect 5728 51451 5800 51452
rect 5852 51451 5924 51452
rect 5976 51451 6048 51452
rect 6100 51451 6172 51452
rect 6224 51451 6296 51452
rect 6348 51451 6420 51452
rect 6472 51451 6544 51452
rect 6596 51451 6668 51452
rect 6720 51451 6792 51452
rect 6844 51451 6916 51452
rect 6968 51451 7040 51452
rect 7092 51451 7886 51452
rect 7938 51451 8010 51452
rect 8062 51451 8134 51452
rect 8186 51451 8258 51452
rect 8310 51451 8382 51452
rect 8434 51451 8506 51452
rect 8558 51451 8630 51452
rect 8682 51451 8754 51452
rect 8806 51451 8878 51452
rect 8930 51451 9002 51452
rect 9054 51451 9126 51452
rect 9178 51451 9250 51452
rect 9302 51451 9374 51452
rect 9426 51451 9498 51452
rect 9550 51451 9622 51452
rect 9674 51451 9746 51452
rect 9798 51451 10251 51452
rect 10303 51451 10375 51452
rect 10427 51451 10499 51452
rect 10551 51451 10623 51452
rect 10675 51451 10747 51452
rect 10799 51451 10871 51452
rect 10923 51451 10995 51452
rect 11047 51451 11119 51452
rect 11171 51451 11243 51452
rect 11295 51451 11367 51452
rect 11419 51451 11489 51452
rect 3489 51439 11489 51451
rect 11651 51260 11662 51818
rect 3316 51249 11662 51260
rect 3316 51234 3424 51249
rect 3162 51203 3424 51234
rect 11554 51234 11662 51249
rect 11708 51234 11816 51844
rect 11554 51203 11816 51234
rect 3162 51170 4863 51203
rect 4915 51170 4987 51203
rect 5039 51170 7277 51203
rect 7329 51170 7401 51203
rect 7453 51170 7525 51203
rect 7577 51170 7649 51203
rect 7701 51170 9939 51203
rect 9991 51170 10063 51203
rect 10115 51170 11816 51203
rect 3162 51098 11816 51170
rect 3162 51095 4863 51098
rect 4915 51095 4987 51098
rect 5039 51095 7277 51098
rect 7329 51095 7401 51098
rect 7453 51095 7525 51098
rect 7577 51095 7649 51098
rect 7701 51095 9939 51098
rect 9991 51095 10063 51098
rect 10115 51095 11816 51098
rect 3162 51049 3330 51095
rect 11648 51049 11816 51095
rect 3162 51046 4863 51049
rect 4915 51046 4987 51049
rect 5039 51046 7277 51049
rect 7329 51046 7401 51049
rect 7453 51046 7525 51049
rect 7577 51046 7649 51049
rect 7701 51046 9939 51049
rect 9991 51046 10063 51049
rect 10115 51046 11816 51049
rect 3162 50974 11816 51046
rect 3162 50941 4863 50974
rect 4915 50941 4987 50974
rect 5039 50941 7277 50974
rect 7329 50941 7401 50974
rect 7453 50941 7525 50974
rect 7577 50941 7649 50974
rect 7701 50941 9939 50974
rect 9991 50941 10063 50974
rect 10115 50941 11816 50974
rect 3162 50910 3424 50941
rect 3162 50300 3270 50910
rect 3316 50895 3424 50910
rect 11554 50910 11816 50941
rect 11554 50895 11662 50910
rect 3316 50884 11662 50895
rect 3316 50326 3327 50884
rect 3489 50693 11489 50705
rect 3489 50692 3559 50693
rect 3611 50692 3683 50693
rect 3735 50692 3807 50693
rect 3859 50692 3931 50693
rect 3983 50692 4055 50693
rect 4107 50692 4179 50693
rect 4231 50692 4303 50693
rect 4355 50692 4427 50693
rect 4479 50692 4551 50693
rect 4603 50692 4675 50693
rect 4727 50692 5180 50693
rect 5232 50692 5304 50693
rect 5356 50692 5428 50693
rect 5480 50692 5552 50693
rect 5604 50692 5676 50693
rect 5728 50692 5800 50693
rect 5852 50692 5924 50693
rect 5976 50692 6048 50693
rect 6100 50692 6172 50693
rect 6224 50692 6296 50693
rect 6348 50692 6420 50693
rect 6472 50692 6544 50693
rect 6596 50692 6668 50693
rect 6720 50692 6792 50693
rect 6844 50692 6916 50693
rect 6968 50692 7040 50693
rect 7092 50692 7886 50693
rect 7938 50692 8010 50693
rect 8062 50692 8134 50693
rect 8186 50692 8258 50693
rect 8310 50692 8382 50693
rect 8434 50692 8506 50693
rect 8558 50692 8630 50693
rect 8682 50692 8754 50693
rect 8806 50692 8878 50693
rect 8930 50692 9002 50693
rect 9054 50692 9126 50693
rect 9178 50692 9250 50693
rect 9302 50692 9374 50693
rect 9426 50692 9498 50693
rect 9550 50692 9622 50693
rect 9674 50692 9746 50693
rect 9798 50692 10251 50693
rect 10303 50692 10375 50693
rect 10427 50692 10499 50693
rect 10551 50692 10623 50693
rect 10675 50692 10747 50693
rect 10799 50692 10871 50693
rect 10923 50692 10995 50693
rect 11047 50692 11119 50693
rect 11171 50692 11243 50693
rect 11295 50692 11367 50693
rect 11419 50692 11489 50693
rect 3489 50646 3502 50692
rect 11476 50646 11489 50692
rect 3489 50641 3559 50646
rect 3611 50641 3683 50646
rect 3735 50641 3807 50646
rect 3859 50641 3931 50646
rect 3983 50641 4055 50646
rect 4107 50641 4179 50646
rect 4231 50641 4303 50646
rect 4355 50641 4427 50646
rect 4479 50641 4551 50646
rect 4603 50641 4675 50646
rect 4727 50641 5180 50646
rect 5232 50641 5304 50646
rect 5356 50641 5428 50646
rect 5480 50641 5552 50646
rect 5604 50641 5676 50646
rect 5728 50641 5800 50646
rect 5852 50641 5924 50646
rect 5976 50641 6048 50646
rect 6100 50641 6172 50646
rect 6224 50641 6296 50646
rect 6348 50641 6420 50646
rect 6472 50641 6544 50646
rect 6596 50641 6668 50646
rect 6720 50641 6792 50646
rect 6844 50641 6916 50646
rect 6968 50641 7040 50646
rect 7092 50641 7886 50646
rect 7938 50641 8010 50646
rect 8062 50641 8134 50646
rect 8186 50641 8258 50646
rect 8310 50641 8382 50646
rect 8434 50641 8506 50646
rect 8558 50641 8630 50646
rect 8682 50641 8754 50646
rect 8806 50641 8878 50646
rect 8930 50641 9002 50646
rect 9054 50641 9126 50646
rect 9178 50641 9250 50646
rect 9302 50641 9374 50646
rect 9426 50641 9498 50646
rect 9550 50641 9622 50646
rect 9674 50641 9746 50646
rect 9798 50641 10251 50646
rect 10303 50641 10375 50646
rect 10427 50641 10499 50646
rect 10551 50641 10623 50646
rect 10675 50641 10747 50646
rect 10799 50641 10871 50646
rect 10923 50641 10995 50646
rect 11047 50641 11119 50646
rect 11171 50641 11243 50646
rect 11295 50641 11367 50646
rect 11419 50641 11489 50646
rect 3489 50569 11489 50641
rect 3489 50564 3559 50569
rect 3611 50564 3683 50569
rect 3735 50564 3807 50569
rect 3859 50564 3931 50569
rect 3983 50564 4055 50569
rect 4107 50564 4179 50569
rect 4231 50564 4303 50569
rect 4355 50564 4427 50569
rect 4479 50564 4551 50569
rect 4603 50564 4675 50569
rect 4727 50564 5180 50569
rect 5232 50564 5304 50569
rect 5356 50564 5428 50569
rect 5480 50564 5552 50569
rect 5604 50564 5676 50569
rect 5728 50564 5800 50569
rect 5852 50564 5924 50569
rect 5976 50564 6048 50569
rect 6100 50564 6172 50569
rect 6224 50564 6296 50569
rect 6348 50564 6420 50569
rect 6472 50564 6544 50569
rect 6596 50564 6668 50569
rect 6720 50564 6792 50569
rect 6844 50564 6916 50569
rect 6968 50564 7040 50569
rect 7092 50564 7886 50569
rect 7938 50564 8010 50569
rect 8062 50564 8134 50569
rect 8186 50564 8258 50569
rect 8310 50564 8382 50569
rect 8434 50564 8506 50569
rect 8558 50564 8630 50569
rect 8682 50564 8754 50569
rect 8806 50564 8878 50569
rect 8930 50564 9002 50569
rect 9054 50564 9126 50569
rect 9178 50564 9250 50569
rect 9302 50564 9374 50569
rect 9426 50564 9498 50569
rect 9550 50564 9622 50569
rect 9674 50564 9746 50569
rect 9798 50564 10251 50569
rect 10303 50564 10375 50569
rect 10427 50564 10499 50569
rect 10551 50564 10623 50569
rect 10675 50564 10747 50569
rect 10799 50564 10871 50569
rect 10923 50564 10995 50569
rect 11047 50564 11119 50569
rect 11171 50564 11243 50569
rect 11295 50564 11367 50569
rect 11419 50564 11489 50569
rect 3489 50518 3502 50564
rect 11476 50518 11489 50564
rect 3489 50517 3559 50518
rect 3611 50517 3683 50518
rect 3735 50517 3807 50518
rect 3859 50517 3931 50518
rect 3983 50517 4055 50518
rect 4107 50517 4179 50518
rect 4231 50517 4303 50518
rect 4355 50517 4427 50518
rect 4479 50517 4551 50518
rect 4603 50517 4675 50518
rect 4727 50517 5180 50518
rect 5232 50517 5304 50518
rect 5356 50517 5428 50518
rect 5480 50517 5552 50518
rect 5604 50517 5676 50518
rect 5728 50517 5800 50518
rect 5852 50517 5924 50518
rect 5976 50517 6048 50518
rect 6100 50517 6172 50518
rect 6224 50517 6296 50518
rect 6348 50517 6420 50518
rect 6472 50517 6544 50518
rect 6596 50517 6668 50518
rect 6720 50517 6792 50518
rect 6844 50517 6916 50518
rect 6968 50517 7040 50518
rect 7092 50517 7886 50518
rect 7938 50517 8010 50518
rect 8062 50517 8134 50518
rect 8186 50517 8258 50518
rect 8310 50517 8382 50518
rect 8434 50517 8506 50518
rect 8558 50517 8630 50518
rect 8682 50517 8754 50518
rect 8806 50517 8878 50518
rect 8930 50517 9002 50518
rect 9054 50517 9126 50518
rect 9178 50517 9250 50518
rect 9302 50517 9374 50518
rect 9426 50517 9498 50518
rect 9550 50517 9622 50518
rect 9674 50517 9746 50518
rect 9798 50517 10251 50518
rect 10303 50517 10375 50518
rect 10427 50517 10499 50518
rect 10551 50517 10623 50518
rect 10675 50517 10747 50518
rect 10799 50517 10871 50518
rect 10923 50517 10995 50518
rect 11047 50517 11119 50518
rect 11171 50517 11243 50518
rect 11295 50517 11367 50518
rect 11419 50517 11489 50518
rect 3489 50505 11489 50517
rect 11651 50326 11662 50884
rect 3316 50315 11662 50326
rect 3316 50300 3424 50315
rect 3162 50269 3424 50300
rect 11554 50300 11662 50315
rect 11708 50300 11816 50910
rect 11554 50269 11816 50300
rect 3162 50236 4863 50269
rect 4915 50236 4987 50269
rect 5039 50236 7277 50269
rect 7329 50236 7401 50269
rect 7453 50236 7525 50269
rect 7577 50236 7649 50269
rect 7701 50236 9939 50269
rect 9991 50236 10063 50269
rect 10115 50236 11816 50269
rect 3162 50164 11816 50236
rect 3162 50161 4863 50164
rect 4915 50161 4987 50164
rect 5039 50161 7277 50164
rect 7329 50161 7401 50164
rect 7453 50161 7525 50164
rect 7577 50161 7649 50164
rect 7701 50161 9939 50164
rect 9991 50161 10063 50164
rect 10115 50161 11816 50164
rect 3162 50115 3330 50161
rect 11648 50115 11816 50161
rect 3162 50112 4863 50115
rect 4915 50112 4987 50115
rect 5039 50112 7277 50115
rect 7329 50112 7401 50115
rect 7453 50112 7525 50115
rect 7577 50112 7649 50115
rect 7701 50112 9939 50115
rect 9991 50112 10063 50115
rect 10115 50112 11816 50115
rect 3162 50040 11816 50112
rect 3162 50007 4863 50040
rect 4915 50007 4987 50040
rect 5039 50007 7277 50040
rect 7329 50007 7401 50040
rect 7453 50007 7525 50040
rect 7577 50007 7649 50040
rect 7701 50007 9939 50040
rect 9991 50007 10063 50040
rect 10115 50007 11816 50040
rect 3162 49976 3424 50007
rect 3162 49366 3270 49976
rect 3316 49961 3424 49976
rect 11554 49976 11816 50007
rect 11554 49961 11662 49976
rect 3316 49950 11662 49961
rect 3316 49392 3327 49950
rect 3489 49759 11489 49771
rect 3489 49758 3559 49759
rect 3611 49758 3683 49759
rect 3735 49758 3807 49759
rect 3859 49758 3931 49759
rect 3983 49758 4055 49759
rect 4107 49758 4179 49759
rect 4231 49758 4303 49759
rect 4355 49758 4427 49759
rect 4479 49758 4551 49759
rect 4603 49758 4675 49759
rect 4727 49758 5180 49759
rect 5232 49758 5304 49759
rect 5356 49758 5428 49759
rect 5480 49758 5552 49759
rect 5604 49758 5676 49759
rect 5728 49758 5800 49759
rect 5852 49758 5924 49759
rect 5976 49758 6048 49759
rect 6100 49758 6172 49759
rect 6224 49758 6296 49759
rect 6348 49758 6420 49759
rect 6472 49758 6544 49759
rect 6596 49758 6668 49759
rect 6720 49758 6792 49759
rect 6844 49758 6916 49759
rect 6968 49758 7040 49759
rect 7092 49758 7886 49759
rect 7938 49758 8010 49759
rect 8062 49758 8134 49759
rect 8186 49758 8258 49759
rect 8310 49758 8382 49759
rect 8434 49758 8506 49759
rect 8558 49758 8630 49759
rect 8682 49758 8754 49759
rect 8806 49758 8878 49759
rect 8930 49758 9002 49759
rect 9054 49758 9126 49759
rect 9178 49758 9250 49759
rect 9302 49758 9374 49759
rect 9426 49758 9498 49759
rect 9550 49758 9622 49759
rect 9674 49758 9746 49759
rect 9798 49758 10251 49759
rect 10303 49758 10375 49759
rect 10427 49758 10499 49759
rect 10551 49758 10623 49759
rect 10675 49758 10747 49759
rect 10799 49758 10871 49759
rect 10923 49758 10995 49759
rect 11047 49758 11119 49759
rect 11171 49758 11243 49759
rect 11295 49758 11367 49759
rect 11419 49758 11489 49759
rect 3489 49712 3502 49758
rect 11476 49712 11489 49758
rect 3489 49707 3559 49712
rect 3611 49707 3683 49712
rect 3735 49707 3807 49712
rect 3859 49707 3931 49712
rect 3983 49707 4055 49712
rect 4107 49707 4179 49712
rect 4231 49707 4303 49712
rect 4355 49707 4427 49712
rect 4479 49707 4551 49712
rect 4603 49707 4675 49712
rect 4727 49707 5180 49712
rect 5232 49707 5304 49712
rect 5356 49707 5428 49712
rect 5480 49707 5552 49712
rect 5604 49707 5676 49712
rect 5728 49707 5800 49712
rect 5852 49707 5924 49712
rect 5976 49707 6048 49712
rect 6100 49707 6172 49712
rect 6224 49707 6296 49712
rect 6348 49707 6420 49712
rect 6472 49707 6544 49712
rect 6596 49707 6668 49712
rect 6720 49707 6792 49712
rect 6844 49707 6916 49712
rect 6968 49707 7040 49712
rect 7092 49707 7886 49712
rect 7938 49707 8010 49712
rect 8062 49707 8134 49712
rect 8186 49707 8258 49712
rect 8310 49707 8382 49712
rect 8434 49707 8506 49712
rect 8558 49707 8630 49712
rect 8682 49707 8754 49712
rect 8806 49707 8878 49712
rect 8930 49707 9002 49712
rect 9054 49707 9126 49712
rect 9178 49707 9250 49712
rect 9302 49707 9374 49712
rect 9426 49707 9498 49712
rect 9550 49707 9622 49712
rect 9674 49707 9746 49712
rect 9798 49707 10251 49712
rect 10303 49707 10375 49712
rect 10427 49707 10499 49712
rect 10551 49707 10623 49712
rect 10675 49707 10747 49712
rect 10799 49707 10871 49712
rect 10923 49707 10995 49712
rect 11047 49707 11119 49712
rect 11171 49707 11243 49712
rect 11295 49707 11367 49712
rect 11419 49707 11489 49712
rect 3489 49635 11489 49707
rect 3489 49630 3559 49635
rect 3611 49630 3683 49635
rect 3735 49630 3807 49635
rect 3859 49630 3931 49635
rect 3983 49630 4055 49635
rect 4107 49630 4179 49635
rect 4231 49630 4303 49635
rect 4355 49630 4427 49635
rect 4479 49630 4551 49635
rect 4603 49630 4675 49635
rect 4727 49630 5180 49635
rect 5232 49630 5304 49635
rect 5356 49630 5428 49635
rect 5480 49630 5552 49635
rect 5604 49630 5676 49635
rect 5728 49630 5800 49635
rect 5852 49630 5924 49635
rect 5976 49630 6048 49635
rect 6100 49630 6172 49635
rect 6224 49630 6296 49635
rect 6348 49630 6420 49635
rect 6472 49630 6544 49635
rect 6596 49630 6668 49635
rect 6720 49630 6792 49635
rect 6844 49630 6916 49635
rect 6968 49630 7040 49635
rect 7092 49630 7886 49635
rect 7938 49630 8010 49635
rect 8062 49630 8134 49635
rect 8186 49630 8258 49635
rect 8310 49630 8382 49635
rect 8434 49630 8506 49635
rect 8558 49630 8630 49635
rect 8682 49630 8754 49635
rect 8806 49630 8878 49635
rect 8930 49630 9002 49635
rect 9054 49630 9126 49635
rect 9178 49630 9250 49635
rect 9302 49630 9374 49635
rect 9426 49630 9498 49635
rect 9550 49630 9622 49635
rect 9674 49630 9746 49635
rect 9798 49630 10251 49635
rect 10303 49630 10375 49635
rect 10427 49630 10499 49635
rect 10551 49630 10623 49635
rect 10675 49630 10747 49635
rect 10799 49630 10871 49635
rect 10923 49630 10995 49635
rect 11047 49630 11119 49635
rect 11171 49630 11243 49635
rect 11295 49630 11367 49635
rect 11419 49630 11489 49635
rect 3489 49584 3502 49630
rect 11476 49584 11489 49630
rect 3489 49583 3559 49584
rect 3611 49583 3683 49584
rect 3735 49583 3807 49584
rect 3859 49583 3931 49584
rect 3983 49583 4055 49584
rect 4107 49583 4179 49584
rect 4231 49583 4303 49584
rect 4355 49583 4427 49584
rect 4479 49583 4551 49584
rect 4603 49583 4675 49584
rect 4727 49583 5180 49584
rect 5232 49583 5304 49584
rect 5356 49583 5428 49584
rect 5480 49583 5552 49584
rect 5604 49583 5676 49584
rect 5728 49583 5800 49584
rect 5852 49583 5924 49584
rect 5976 49583 6048 49584
rect 6100 49583 6172 49584
rect 6224 49583 6296 49584
rect 6348 49583 6420 49584
rect 6472 49583 6544 49584
rect 6596 49583 6668 49584
rect 6720 49583 6792 49584
rect 6844 49583 6916 49584
rect 6968 49583 7040 49584
rect 7092 49583 7886 49584
rect 7938 49583 8010 49584
rect 8062 49583 8134 49584
rect 8186 49583 8258 49584
rect 8310 49583 8382 49584
rect 8434 49583 8506 49584
rect 8558 49583 8630 49584
rect 8682 49583 8754 49584
rect 8806 49583 8878 49584
rect 8930 49583 9002 49584
rect 9054 49583 9126 49584
rect 9178 49583 9250 49584
rect 9302 49583 9374 49584
rect 9426 49583 9498 49584
rect 9550 49583 9622 49584
rect 9674 49583 9746 49584
rect 9798 49583 10251 49584
rect 10303 49583 10375 49584
rect 10427 49583 10499 49584
rect 10551 49583 10623 49584
rect 10675 49583 10747 49584
rect 10799 49583 10871 49584
rect 10923 49583 10995 49584
rect 11047 49583 11119 49584
rect 11171 49583 11243 49584
rect 11295 49583 11367 49584
rect 11419 49583 11489 49584
rect 3489 49571 11489 49583
rect 11651 49392 11662 49950
rect 3316 49381 11662 49392
rect 3316 49366 3424 49381
rect 3162 49335 3424 49366
rect 11554 49366 11662 49381
rect 11708 49366 11816 49976
rect 11554 49335 11816 49366
rect 3162 49302 4863 49335
rect 4915 49302 4987 49335
rect 5039 49302 7277 49335
rect 7329 49302 7401 49335
rect 7453 49302 7525 49335
rect 7577 49302 7649 49335
rect 7701 49302 9939 49335
rect 9991 49302 10063 49335
rect 10115 49302 11816 49335
rect 3162 49230 11816 49302
rect 3162 49227 4863 49230
rect 4915 49227 4987 49230
rect 5039 49227 7277 49230
rect 7329 49227 7401 49230
rect 7453 49227 7525 49230
rect 7577 49227 7649 49230
rect 7701 49227 9939 49230
rect 9991 49227 10063 49230
rect 10115 49227 11816 49230
rect 3162 49181 3330 49227
rect 11648 49181 11816 49227
rect 3162 49178 4863 49181
rect 4915 49178 4987 49181
rect 5039 49178 7277 49181
rect 7329 49178 7401 49181
rect 7453 49178 7525 49181
rect 7577 49178 7649 49181
rect 7701 49178 9939 49181
rect 9991 49178 10063 49181
rect 10115 49178 11816 49181
rect 3162 49106 11816 49178
rect 3162 49073 4863 49106
rect 4915 49073 4987 49106
rect 5039 49073 7277 49106
rect 7329 49073 7401 49106
rect 7453 49073 7525 49106
rect 7577 49073 7649 49106
rect 7701 49073 9939 49106
rect 9991 49073 10063 49106
rect 10115 49073 11816 49106
rect 3162 49042 3424 49073
rect 3162 48432 3270 49042
rect 3316 49027 3424 49042
rect 11554 49042 11816 49073
rect 11554 49027 11662 49042
rect 3316 49016 11662 49027
rect 3316 48458 3327 49016
rect 3489 48825 11489 48837
rect 3489 48824 3559 48825
rect 3611 48824 3683 48825
rect 3735 48824 3807 48825
rect 3859 48824 3931 48825
rect 3983 48824 4055 48825
rect 4107 48824 4179 48825
rect 4231 48824 4303 48825
rect 4355 48824 4427 48825
rect 4479 48824 4551 48825
rect 4603 48824 4675 48825
rect 4727 48824 5180 48825
rect 5232 48824 5304 48825
rect 5356 48824 5428 48825
rect 5480 48824 5552 48825
rect 5604 48824 5676 48825
rect 5728 48824 5800 48825
rect 5852 48824 5924 48825
rect 5976 48824 6048 48825
rect 6100 48824 6172 48825
rect 6224 48824 6296 48825
rect 6348 48824 6420 48825
rect 6472 48824 6544 48825
rect 6596 48824 6668 48825
rect 6720 48824 6792 48825
rect 6844 48824 6916 48825
rect 6968 48824 7040 48825
rect 7092 48824 7886 48825
rect 7938 48824 8010 48825
rect 8062 48824 8134 48825
rect 8186 48824 8258 48825
rect 8310 48824 8382 48825
rect 8434 48824 8506 48825
rect 8558 48824 8630 48825
rect 8682 48824 8754 48825
rect 8806 48824 8878 48825
rect 8930 48824 9002 48825
rect 9054 48824 9126 48825
rect 9178 48824 9250 48825
rect 9302 48824 9374 48825
rect 9426 48824 9498 48825
rect 9550 48824 9622 48825
rect 9674 48824 9746 48825
rect 9798 48824 10251 48825
rect 10303 48824 10375 48825
rect 10427 48824 10499 48825
rect 10551 48824 10623 48825
rect 10675 48824 10747 48825
rect 10799 48824 10871 48825
rect 10923 48824 10995 48825
rect 11047 48824 11119 48825
rect 11171 48824 11243 48825
rect 11295 48824 11367 48825
rect 11419 48824 11489 48825
rect 3489 48778 3502 48824
rect 11476 48778 11489 48824
rect 3489 48773 3559 48778
rect 3611 48773 3683 48778
rect 3735 48773 3807 48778
rect 3859 48773 3931 48778
rect 3983 48773 4055 48778
rect 4107 48773 4179 48778
rect 4231 48773 4303 48778
rect 4355 48773 4427 48778
rect 4479 48773 4551 48778
rect 4603 48773 4675 48778
rect 4727 48773 5180 48778
rect 5232 48773 5304 48778
rect 5356 48773 5428 48778
rect 5480 48773 5552 48778
rect 5604 48773 5676 48778
rect 5728 48773 5800 48778
rect 5852 48773 5924 48778
rect 5976 48773 6048 48778
rect 6100 48773 6172 48778
rect 6224 48773 6296 48778
rect 6348 48773 6420 48778
rect 6472 48773 6544 48778
rect 6596 48773 6668 48778
rect 6720 48773 6792 48778
rect 6844 48773 6916 48778
rect 6968 48773 7040 48778
rect 7092 48773 7886 48778
rect 7938 48773 8010 48778
rect 8062 48773 8134 48778
rect 8186 48773 8258 48778
rect 8310 48773 8382 48778
rect 8434 48773 8506 48778
rect 8558 48773 8630 48778
rect 8682 48773 8754 48778
rect 8806 48773 8878 48778
rect 8930 48773 9002 48778
rect 9054 48773 9126 48778
rect 9178 48773 9250 48778
rect 9302 48773 9374 48778
rect 9426 48773 9498 48778
rect 9550 48773 9622 48778
rect 9674 48773 9746 48778
rect 9798 48773 10251 48778
rect 10303 48773 10375 48778
rect 10427 48773 10499 48778
rect 10551 48773 10623 48778
rect 10675 48773 10747 48778
rect 10799 48773 10871 48778
rect 10923 48773 10995 48778
rect 11047 48773 11119 48778
rect 11171 48773 11243 48778
rect 11295 48773 11367 48778
rect 11419 48773 11489 48778
rect 3489 48701 11489 48773
rect 3489 48696 3559 48701
rect 3611 48696 3683 48701
rect 3735 48696 3807 48701
rect 3859 48696 3931 48701
rect 3983 48696 4055 48701
rect 4107 48696 4179 48701
rect 4231 48696 4303 48701
rect 4355 48696 4427 48701
rect 4479 48696 4551 48701
rect 4603 48696 4675 48701
rect 4727 48696 5180 48701
rect 5232 48696 5304 48701
rect 5356 48696 5428 48701
rect 5480 48696 5552 48701
rect 5604 48696 5676 48701
rect 5728 48696 5800 48701
rect 5852 48696 5924 48701
rect 5976 48696 6048 48701
rect 6100 48696 6172 48701
rect 6224 48696 6296 48701
rect 6348 48696 6420 48701
rect 6472 48696 6544 48701
rect 6596 48696 6668 48701
rect 6720 48696 6792 48701
rect 6844 48696 6916 48701
rect 6968 48696 7040 48701
rect 7092 48696 7886 48701
rect 7938 48696 8010 48701
rect 8062 48696 8134 48701
rect 8186 48696 8258 48701
rect 8310 48696 8382 48701
rect 8434 48696 8506 48701
rect 8558 48696 8630 48701
rect 8682 48696 8754 48701
rect 8806 48696 8878 48701
rect 8930 48696 9002 48701
rect 9054 48696 9126 48701
rect 9178 48696 9250 48701
rect 9302 48696 9374 48701
rect 9426 48696 9498 48701
rect 9550 48696 9622 48701
rect 9674 48696 9746 48701
rect 9798 48696 10251 48701
rect 10303 48696 10375 48701
rect 10427 48696 10499 48701
rect 10551 48696 10623 48701
rect 10675 48696 10747 48701
rect 10799 48696 10871 48701
rect 10923 48696 10995 48701
rect 11047 48696 11119 48701
rect 11171 48696 11243 48701
rect 11295 48696 11367 48701
rect 11419 48696 11489 48701
rect 3489 48650 3502 48696
rect 11476 48650 11489 48696
rect 3489 48649 3559 48650
rect 3611 48649 3683 48650
rect 3735 48649 3807 48650
rect 3859 48649 3931 48650
rect 3983 48649 4055 48650
rect 4107 48649 4179 48650
rect 4231 48649 4303 48650
rect 4355 48649 4427 48650
rect 4479 48649 4551 48650
rect 4603 48649 4675 48650
rect 4727 48649 5180 48650
rect 5232 48649 5304 48650
rect 5356 48649 5428 48650
rect 5480 48649 5552 48650
rect 5604 48649 5676 48650
rect 5728 48649 5800 48650
rect 5852 48649 5924 48650
rect 5976 48649 6048 48650
rect 6100 48649 6172 48650
rect 6224 48649 6296 48650
rect 6348 48649 6420 48650
rect 6472 48649 6544 48650
rect 6596 48649 6668 48650
rect 6720 48649 6792 48650
rect 6844 48649 6916 48650
rect 6968 48649 7040 48650
rect 7092 48649 7886 48650
rect 7938 48649 8010 48650
rect 8062 48649 8134 48650
rect 8186 48649 8258 48650
rect 8310 48649 8382 48650
rect 8434 48649 8506 48650
rect 8558 48649 8630 48650
rect 8682 48649 8754 48650
rect 8806 48649 8878 48650
rect 8930 48649 9002 48650
rect 9054 48649 9126 48650
rect 9178 48649 9250 48650
rect 9302 48649 9374 48650
rect 9426 48649 9498 48650
rect 9550 48649 9622 48650
rect 9674 48649 9746 48650
rect 9798 48649 10251 48650
rect 10303 48649 10375 48650
rect 10427 48649 10499 48650
rect 10551 48649 10623 48650
rect 10675 48649 10747 48650
rect 10799 48649 10871 48650
rect 10923 48649 10995 48650
rect 11047 48649 11119 48650
rect 11171 48649 11243 48650
rect 11295 48649 11367 48650
rect 11419 48649 11489 48650
rect 3489 48637 11489 48649
rect 11651 48458 11662 49016
rect 3316 48447 11662 48458
rect 3316 48432 3424 48447
rect 3162 48401 3424 48432
rect 11554 48432 11662 48447
rect 11708 48432 11816 49042
rect 11554 48401 11816 48432
rect 3162 48383 4863 48401
rect 4915 48383 4987 48401
rect 5039 48383 7277 48401
rect 7329 48383 7401 48401
rect 7453 48383 7525 48401
rect 7577 48383 7649 48401
rect 7701 48383 9939 48401
rect 9991 48383 10063 48401
rect 10115 48383 11816 48401
rect 3162 48376 11816 48383
rect 11862 48376 11873 51900
rect 3105 48311 11873 48376
rect 3105 48293 4863 48311
rect 4915 48293 4987 48311
rect 5039 48293 7277 48311
rect 7329 48293 7401 48311
rect 7453 48293 7525 48311
rect 7577 48293 7649 48311
rect 7701 48293 9939 48311
rect 9991 48293 10063 48311
rect 10115 48293 11873 48311
rect 3105 48247 3142 48293
rect 11836 48247 11873 48293
rect 3105 48236 11873 48247
rect 12059 48022 12070 52254
rect 2908 48011 12070 48022
rect 2908 47988 3016 48011
rect 11962 47988 12070 48011
rect 2908 47936 2934 47988
rect 2986 47936 3016 47988
rect 11962 47936 11992 47988
rect 12044 47936 12070 47988
rect 2908 47864 3016 47936
rect 11962 47864 12070 47936
rect 2908 47812 2934 47864
rect 2986 47812 3016 47864
rect 11962 47812 11992 47864
rect 12044 47812 12070 47864
rect 2908 47740 3016 47812
rect 11962 47740 12070 47812
rect 2908 47688 2934 47740
rect 2986 47688 3016 47740
rect 11962 47688 11992 47740
rect 12044 47688 12070 47740
rect 2908 47665 3016 47688
rect 11962 47665 12070 47688
rect 12416 47665 12427 52611
rect 2551 47654 12427 47665
rect 12753 52611 14907 52622
rect 12753 47665 12764 52611
rect 14710 52586 14907 52611
rect 14710 52574 14968 52586
rect 14710 52522 14904 52574
rect 14956 52522 14968 52574
rect 14710 52466 14968 52522
rect 14710 52414 14904 52466
rect 14956 52414 14968 52466
rect 14710 52358 14968 52414
rect 14710 52306 14904 52358
rect 14956 52306 14968 52358
rect 14710 52250 14968 52306
rect 14710 52198 14904 52250
rect 14956 52198 14968 52250
rect 14710 52142 14968 52198
rect 14710 52090 14904 52142
rect 14956 52090 14968 52142
rect 14710 52034 14968 52090
rect 14710 51982 14904 52034
rect 14956 51982 14968 52034
rect 14710 51926 14968 51982
rect 14710 51874 14904 51926
rect 14956 51874 14968 51926
rect 14710 51818 14968 51874
rect 14710 51766 14904 51818
rect 14956 51766 14968 51818
rect 14710 51710 14968 51766
rect 14710 51658 14904 51710
rect 14956 51658 14968 51710
rect 14710 51622 14968 51658
rect 14710 51422 14721 51622
rect 14892 51602 14968 51622
rect 14892 51550 14904 51602
rect 14956 51550 14968 51602
rect 14892 51494 14968 51550
rect 14892 51442 14904 51494
rect 14956 51442 14968 51494
rect 14892 51422 14968 51442
rect 14710 51386 14968 51422
rect 14710 51334 14904 51386
rect 14956 51334 14968 51386
rect 14710 51278 14968 51334
rect 14710 51226 14904 51278
rect 14956 51226 14968 51278
rect 14710 51214 14968 51226
rect 14710 50422 14907 51214
rect 14710 49854 14721 50422
rect 14710 48854 14907 49854
rect 14710 48654 14721 48854
rect 14710 47665 14907 48654
rect 12753 47654 14907 47665
rect 71 42647 725 42658
rect 71 41658 268 42647
rect 257 41458 268 41658
rect 71 40458 268 41458
rect 257 40258 268 40458
rect 71 39258 268 40258
rect 257 39058 268 39258
rect 71 38186 268 39058
rect 10 38174 268 38186
rect 10 38122 22 38174
rect 74 38122 268 38174
rect 10 38066 268 38122
rect 10 38014 22 38066
rect 74 38058 268 38066
rect 74 38014 86 38058
rect 10 37958 86 38014
rect 10 37906 22 37958
rect 74 37906 86 37958
rect 10 37858 86 37906
rect 257 37858 268 38058
rect 10 37850 268 37858
rect 10 37798 22 37850
rect 74 37798 268 37850
rect 10 37742 268 37798
rect 10 37690 22 37742
rect 74 37690 268 37742
rect 10 37634 268 37690
rect 10 37582 22 37634
rect 74 37582 268 37634
rect 10 37526 268 37582
rect 10 37474 22 37526
rect 74 37474 268 37526
rect 10 37418 268 37474
rect 10 37366 22 37418
rect 74 37366 268 37418
rect 10 37310 268 37366
rect 10 37258 22 37310
rect 74 37258 268 37310
rect 10 37202 268 37258
rect 10 37150 22 37202
rect 74 37150 268 37202
rect 10 37094 268 37150
rect 10 37042 22 37094
rect 74 37042 268 37094
rect 10 36986 268 37042
rect 10 36934 22 36986
rect 74 36934 268 36986
rect 10 36878 268 36934
rect 10 36826 22 36878
rect 74 36858 268 36878
rect 74 36826 86 36858
rect 10 36814 86 36826
rect 257 36658 268 36858
rect 71 35658 268 36658
rect 257 35458 268 35658
rect 71 34458 268 35458
rect 257 34258 268 34458
rect 71 33258 268 34258
rect 257 33058 268 33258
rect 71 32058 268 33058
rect 257 31858 268 32058
rect 71 30858 268 31858
rect 257 30658 268 30858
rect 71 29658 268 30658
rect 257 29458 268 29658
rect 71 28458 268 29458
rect 257 28258 268 28458
rect 71 27258 268 28258
rect 257 27058 268 27258
rect 71 26058 268 27058
rect 257 25858 268 26058
rect 71 24858 268 25858
rect 257 24658 268 24858
rect 71 23658 268 24658
rect 257 23458 268 23658
rect 71 22458 268 23458
rect 257 21390 268 22458
rect 71 20390 268 21390
rect 257 20190 268 20390
rect 71 19190 268 20190
rect 257 18990 268 19190
rect 71 17990 268 18990
rect 257 17790 268 17990
rect 71 16790 268 17790
rect 257 16590 268 16790
rect 71 15590 268 16590
rect 257 15390 268 15590
rect 71 14390 268 15390
rect 257 14190 268 14390
rect 71 13190 268 14190
rect 257 12990 268 13190
rect 71 11990 268 12990
rect 257 11790 268 11990
rect 71 10790 268 11790
rect 257 10590 268 10790
rect 71 9590 268 10590
rect 257 9390 268 9590
rect 71 8390 268 9390
rect 257 8190 268 8390
rect 71 7190 268 8190
rect 257 6990 268 7190
rect 71 5990 268 6990
rect 257 5790 268 5990
rect 71 4790 268 5790
rect 257 4590 268 4790
rect 71 3590 268 4590
rect 257 3390 268 3590
rect 71 2390 268 3390
rect 257 2190 268 2390
rect 71 1201 268 2190
rect 714 1201 725 42647
rect 13012 42647 14907 42658
rect 13012 27201 13023 42647
rect 13969 41658 14264 42647
rect 13969 41458 13980 41658
rect 14253 41458 14264 41658
rect 13969 40458 14264 41458
rect 13969 40258 13980 40458
rect 14253 40258 14264 40458
rect 13969 39258 14264 40258
rect 13969 39058 13980 39258
rect 14253 39058 14264 39258
rect 13969 38058 14264 39058
rect 13969 37858 13980 38058
rect 14253 37858 14264 38058
rect 13969 36858 14264 37858
rect 13969 36658 13980 36858
rect 14253 36658 14264 36858
rect 13969 35658 14264 36658
rect 13969 35458 13980 35658
rect 14253 35458 14264 35658
rect 13969 34458 14264 35458
rect 13969 34258 13980 34458
rect 14253 34258 14264 34458
rect 13969 33258 14264 34258
rect 13969 33058 13980 33258
rect 14253 33058 14264 33258
rect 13969 32058 14264 33058
rect 13969 31858 13980 32058
rect 14253 31858 14264 32058
rect 13969 30858 14264 31858
rect 13969 30658 13980 30858
rect 14253 30658 14264 30858
rect 13969 29658 14264 30658
rect 13969 29458 13980 29658
rect 14253 29458 14264 29658
rect 13969 28458 14264 29458
rect 13969 28190 13980 28458
rect 14253 28190 14264 28458
rect 13969 27201 14264 28190
rect 13012 27190 14264 27201
rect 71 1190 725 1201
rect 14253 1201 14264 27190
rect 14710 41658 14907 42647
rect 14710 41458 14721 41658
rect 14710 40458 14907 41458
rect 14710 40258 14721 40458
rect 14710 39258 14907 40258
rect 14710 39058 14721 39258
rect 14710 38186 14907 39058
rect 14710 38174 14968 38186
rect 14710 38122 14904 38174
rect 14956 38122 14968 38174
rect 14710 38066 14968 38122
rect 14710 38058 14904 38066
rect 14710 37858 14721 38058
rect 14892 38014 14904 38058
rect 14956 38014 14968 38066
rect 14892 37958 14968 38014
rect 14892 37906 14904 37958
rect 14956 37906 14968 37958
rect 14892 37858 14968 37906
rect 14710 37850 14968 37858
rect 14710 37798 14904 37850
rect 14956 37798 14968 37850
rect 14710 37742 14968 37798
rect 14710 37690 14904 37742
rect 14956 37690 14968 37742
rect 14710 37634 14968 37690
rect 14710 37582 14904 37634
rect 14956 37582 14968 37634
rect 14710 37526 14968 37582
rect 14710 37474 14904 37526
rect 14956 37474 14968 37526
rect 14710 37418 14968 37474
rect 14710 37366 14904 37418
rect 14956 37366 14968 37418
rect 14710 37310 14968 37366
rect 14710 37258 14904 37310
rect 14956 37258 14968 37310
rect 14710 37202 14968 37258
rect 14710 37150 14904 37202
rect 14956 37150 14968 37202
rect 14710 37094 14968 37150
rect 14710 37042 14904 37094
rect 14956 37042 14968 37094
rect 14710 36986 14968 37042
rect 14710 36934 14904 36986
rect 14956 36934 14968 36986
rect 14710 36878 14968 36934
rect 14710 36858 14904 36878
rect 14710 36658 14721 36858
rect 14892 36826 14904 36858
rect 14956 36826 14968 36878
rect 14892 36814 14968 36826
rect 14710 35658 14907 36658
rect 14710 35458 14721 35658
rect 14710 34458 14907 35458
rect 14710 34258 14721 34458
rect 14710 33258 14907 34258
rect 14710 33058 14721 33258
rect 14710 32058 14907 33058
rect 14710 31858 14721 32058
rect 14710 30858 14907 31858
rect 14710 30658 14721 30858
rect 14710 29658 14907 30658
rect 14710 29458 14721 29658
rect 14710 28458 14907 29458
rect 14710 28258 14721 28458
rect 14710 27258 14907 28258
rect 14710 27058 14721 27258
rect 14710 26058 14907 27058
rect 14710 25858 14721 26058
rect 14710 24858 14907 25858
rect 14710 24658 14721 24858
rect 14710 23658 14907 24658
rect 14710 23458 14721 23658
rect 14710 22458 14907 23458
rect 14710 21390 14721 22458
rect 14710 20390 14907 21390
rect 14710 20190 14721 20390
rect 14710 19190 14907 20190
rect 14710 18990 14721 19190
rect 14710 17990 14907 18990
rect 14710 17790 14721 17990
rect 14710 16790 14907 17790
rect 14710 16590 14721 16790
rect 14710 15590 14907 16590
rect 14710 15390 14721 15590
rect 14710 14390 14907 15390
rect 14710 14190 14721 14390
rect 14710 13190 14907 14190
rect 14710 12990 14721 13190
rect 14710 11990 14907 12990
rect 14710 11790 14721 11990
rect 14710 10790 14907 11790
rect 14710 10590 14721 10790
rect 14710 9590 14907 10590
rect 14710 9390 14721 9590
rect 14710 8390 14907 9390
rect 14710 8190 14721 8390
rect 14710 7190 14907 8190
rect 14710 6990 14721 7190
rect 14710 5990 14907 6990
rect 14710 5790 14721 5990
rect 14710 4790 14907 5790
rect 14710 4590 14721 4790
rect 14710 3590 14907 4590
rect 14710 3390 14721 3590
rect 14710 2390 14907 3390
rect 14710 2190 14721 2390
rect 14710 1201 14907 2190
rect 14253 1190 14907 1201
<< via1 >>
rect 2501 57105 2553 57108
rect 2609 57105 2661 57108
rect 4871 57105 4923 57108
rect 4979 57105 5031 57108
rect 7247 57105 7299 57108
rect 7355 57105 7407 57108
rect 7463 57105 7515 57108
rect 7571 57105 7623 57108
rect 7679 57105 7731 57108
rect 9947 57105 9999 57108
rect 10055 57105 10107 57108
rect 12317 57105 12369 57108
rect 12425 57105 12477 57108
rect 2501 57059 2553 57105
rect 2609 57059 2661 57105
rect 4871 57059 4923 57105
rect 4979 57059 5031 57105
rect 7247 57059 7299 57105
rect 7355 57059 7407 57105
rect 7463 57059 7515 57105
rect 7571 57059 7623 57105
rect 7679 57059 7731 57105
rect 9947 57059 9999 57105
rect 10055 57059 10107 57105
rect 12317 57059 12369 57105
rect 12425 57059 12477 57105
rect 2501 57056 2553 57059
rect 2609 57056 2661 57059
rect 4871 57056 4923 57059
rect 4979 57056 5031 57059
rect 7247 57056 7299 57059
rect 7355 57056 7407 57059
rect 7463 57056 7515 57059
rect 7571 57056 7623 57059
rect 7679 57056 7731 57059
rect 9947 57056 9999 57059
rect 10055 57056 10107 57059
rect 12317 57056 12369 57059
rect 12425 57056 12477 57059
rect 917 56617 969 56669
rect 1041 56617 1093 56669
rect 1165 56617 1217 56669
rect 1289 56617 1341 56669
rect 1413 56617 1465 56669
rect 1537 56617 1589 56669
rect 1661 56617 1713 56669
rect 1785 56617 1837 56669
rect 917 56493 969 56545
rect 1041 56493 1093 56545
rect 1165 56493 1217 56545
rect 1289 56493 1341 56545
rect 1413 56493 1465 56545
rect 1537 56493 1589 56545
rect 1661 56493 1713 56545
rect 1785 56493 1837 56545
rect 917 56369 969 56421
rect 1041 56369 1093 56421
rect 1165 56369 1217 56421
rect 1289 56369 1341 56421
rect 1413 56369 1465 56421
rect 1537 56369 1589 56421
rect 1661 56369 1713 56421
rect 1785 56369 1837 56421
rect 917 56245 969 56297
rect 1041 56245 1093 56297
rect 1165 56245 1217 56297
rect 1289 56245 1341 56297
rect 1413 56245 1465 56297
rect 1537 56245 1589 56297
rect 1661 56245 1713 56297
rect 1785 56245 1837 56297
rect 917 56121 969 56173
rect 1041 56121 1093 56173
rect 1165 56121 1217 56173
rect 1289 56121 1341 56173
rect 1413 56121 1465 56173
rect 1537 56121 1589 56173
rect 1661 56121 1713 56173
rect 1785 56121 1837 56173
rect 917 55997 969 56049
rect 1041 55997 1093 56049
rect 1165 55997 1217 56049
rect 1289 55997 1341 56049
rect 1413 55997 1465 56049
rect 1537 55997 1589 56049
rect 1661 55997 1713 56049
rect 1785 55997 1837 56049
rect 917 55873 969 55925
rect 1041 55873 1093 55925
rect 1165 55873 1217 55925
rect 1289 55873 1341 55925
rect 1413 55873 1465 55925
rect 1537 55873 1589 55925
rect 1661 55873 1713 55925
rect 1785 55873 1837 55925
rect 917 55749 969 55801
rect 1041 55749 1093 55801
rect 1165 55749 1217 55801
rect 1289 55749 1341 55801
rect 1413 55749 1465 55801
rect 1537 55749 1589 55801
rect 1661 55749 1713 55801
rect 1785 55749 1837 55801
rect 917 55625 969 55677
rect 1041 55625 1093 55677
rect 1165 55625 1217 55677
rect 1289 55625 1341 55677
rect 1413 55625 1465 55677
rect 1537 55625 1589 55677
rect 1661 55625 1713 55677
rect 1785 55625 1837 55677
rect 917 55501 969 55553
rect 1041 55501 1093 55553
rect 1165 55501 1217 55553
rect 1289 55501 1341 55553
rect 1413 55501 1465 55553
rect 1537 55501 1589 55553
rect 1661 55501 1713 55553
rect 1785 55501 1837 55553
rect 917 55377 969 55429
rect 1041 55377 1093 55429
rect 1165 55377 1217 55429
rect 1289 55377 1341 55429
rect 1413 55377 1465 55429
rect 1537 55377 1589 55429
rect 1661 55377 1713 55429
rect 1785 55377 1837 55429
rect 917 55253 969 55305
rect 1041 55253 1093 55305
rect 1165 55253 1217 55305
rect 1289 55253 1341 55305
rect 1413 55253 1465 55305
rect 1537 55253 1589 55305
rect 1661 55253 1713 55305
rect 1785 55253 1837 55305
rect 917 55129 969 55181
rect 1041 55129 1093 55181
rect 1165 55129 1217 55181
rect 1289 55129 1341 55181
rect 1413 55129 1465 55181
rect 1537 55129 1589 55181
rect 1661 55129 1713 55181
rect 1785 55129 1837 55181
rect 917 55005 969 55057
rect 1041 55005 1093 55057
rect 1165 55005 1217 55057
rect 1289 55005 1341 55057
rect 1413 55005 1465 55057
rect 1537 55005 1589 55057
rect 1661 55005 1713 55057
rect 1785 55005 1837 55057
rect 917 54881 969 54933
rect 1041 54881 1093 54933
rect 1165 54881 1217 54933
rect 1289 54881 1341 54933
rect 1413 54881 1465 54933
rect 1537 54881 1589 54933
rect 1661 54881 1713 54933
rect 1785 54881 1837 54933
rect 917 54757 969 54809
rect 1041 54757 1093 54809
rect 1165 54757 1217 54809
rect 1289 54757 1341 54809
rect 1413 54757 1465 54809
rect 1537 54757 1589 54809
rect 1661 54757 1713 54809
rect 1785 54757 1837 54809
rect 917 54633 969 54685
rect 1041 54633 1093 54685
rect 1165 54633 1217 54685
rect 1289 54633 1341 54685
rect 1413 54633 1465 54685
rect 1537 54633 1589 54685
rect 1661 54633 1713 54685
rect 1785 54633 1837 54685
rect 917 54509 969 54561
rect 1041 54509 1093 54561
rect 1165 54509 1217 54561
rect 1289 54509 1341 54561
rect 1413 54509 1465 54561
rect 1537 54509 1589 54561
rect 1661 54509 1713 54561
rect 1785 54509 1837 54561
rect 917 54385 969 54437
rect 1041 54385 1093 54437
rect 1165 54385 1217 54437
rect 1289 54385 1341 54437
rect 1413 54385 1465 54437
rect 1537 54385 1589 54437
rect 1661 54385 1713 54437
rect 1785 54385 1837 54437
rect 917 54261 969 54313
rect 1041 54261 1093 54313
rect 1165 54261 1217 54313
rect 1289 54261 1341 54313
rect 1413 54261 1465 54313
rect 1537 54261 1589 54313
rect 1661 54261 1713 54313
rect 1785 54261 1837 54313
rect 917 54137 969 54189
rect 1041 54137 1093 54189
rect 1165 54137 1217 54189
rect 1289 54137 1341 54189
rect 1413 54137 1465 54189
rect 1537 54137 1589 54189
rect 1661 54137 1713 54189
rect 1785 54137 1837 54189
rect 917 54013 969 54065
rect 1041 54013 1093 54065
rect 1165 54013 1217 54065
rect 1289 54013 1341 54065
rect 1413 54013 1465 54065
rect 1537 54013 1589 54065
rect 1661 54013 1713 54065
rect 1785 54013 1837 54065
rect 917 53889 969 53941
rect 1041 53889 1093 53941
rect 1165 53889 1217 53941
rect 1289 53889 1341 53941
rect 1413 53889 1465 53941
rect 1537 53889 1589 53941
rect 1661 53889 1713 53941
rect 1785 53889 1837 53941
rect 917 53765 969 53817
rect 1041 53765 1093 53817
rect 1165 53765 1217 53817
rect 1289 53765 1341 53817
rect 1413 53765 1465 53817
rect 1537 53765 1589 53817
rect 1661 53765 1713 53817
rect 1785 53765 1837 53817
rect 917 53641 969 53693
rect 1041 53641 1093 53693
rect 1165 53641 1217 53693
rect 1289 53641 1341 53693
rect 1413 53641 1465 53693
rect 1537 53641 1589 53693
rect 1661 53641 1713 53693
rect 1785 53641 1837 53693
rect 2833 56617 2885 56669
rect 2957 56617 3009 56669
rect 3081 56617 3133 56669
rect 3205 56617 3257 56669
rect 3329 56617 3381 56669
rect 3453 56617 3505 56669
rect 3577 56617 3629 56669
rect 3701 56617 3753 56669
rect 2833 56493 2885 56545
rect 2957 56493 3009 56545
rect 3081 56493 3133 56545
rect 3205 56493 3257 56545
rect 3329 56493 3381 56545
rect 3453 56493 3505 56545
rect 3577 56493 3629 56545
rect 3701 56493 3753 56545
rect 2833 56369 2885 56421
rect 2957 56369 3009 56421
rect 3081 56369 3133 56421
rect 3205 56369 3257 56421
rect 3329 56369 3381 56421
rect 3453 56369 3505 56421
rect 3577 56369 3629 56421
rect 3701 56369 3753 56421
rect 2833 56245 2885 56297
rect 2957 56245 3009 56297
rect 3081 56245 3133 56297
rect 3205 56245 3257 56297
rect 3329 56245 3381 56297
rect 3453 56245 3505 56297
rect 3577 56245 3629 56297
rect 3701 56245 3753 56297
rect 2833 56121 2885 56173
rect 2957 56121 3009 56173
rect 3081 56121 3133 56173
rect 3205 56121 3257 56173
rect 3329 56121 3381 56173
rect 3453 56121 3505 56173
rect 3577 56121 3629 56173
rect 3701 56121 3753 56173
rect 2833 55997 2885 56049
rect 2957 55997 3009 56049
rect 3081 55997 3133 56049
rect 3205 55997 3257 56049
rect 3329 55997 3381 56049
rect 3453 55997 3505 56049
rect 3577 55997 3629 56049
rect 3701 55997 3753 56049
rect 2833 55873 2885 55925
rect 2957 55873 3009 55925
rect 3081 55873 3133 55925
rect 3205 55873 3257 55925
rect 3329 55873 3381 55925
rect 3453 55873 3505 55925
rect 3577 55873 3629 55925
rect 3701 55873 3753 55925
rect 2833 55749 2885 55801
rect 2957 55749 3009 55801
rect 3081 55749 3133 55801
rect 3205 55749 3257 55801
rect 3329 55749 3381 55801
rect 3453 55749 3505 55801
rect 3577 55749 3629 55801
rect 3701 55749 3753 55801
rect 2833 55625 2885 55677
rect 2957 55625 3009 55677
rect 3081 55625 3133 55677
rect 3205 55625 3257 55677
rect 3329 55625 3381 55677
rect 3453 55625 3505 55677
rect 3577 55625 3629 55677
rect 3701 55625 3753 55677
rect 2833 55501 2885 55553
rect 2957 55501 3009 55553
rect 3081 55501 3133 55553
rect 3205 55501 3257 55553
rect 3329 55501 3381 55553
rect 3453 55501 3505 55553
rect 3577 55501 3629 55553
rect 3701 55501 3753 55553
rect 2833 55377 2885 55429
rect 2957 55377 3009 55429
rect 3081 55377 3133 55429
rect 3205 55377 3257 55429
rect 3329 55377 3381 55429
rect 3453 55377 3505 55429
rect 3577 55377 3629 55429
rect 3701 55377 3753 55429
rect 2833 55253 2885 55305
rect 2957 55253 3009 55305
rect 3081 55253 3133 55305
rect 3205 55253 3257 55305
rect 3329 55253 3381 55305
rect 3453 55253 3505 55305
rect 3577 55253 3629 55305
rect 3701 55253 3753 55305
rect 2833 55129 2885 55181
rect 2957 55129 3009 55181
rect 3081 55129 3133 55181
rect 3205 55129 3257 55181
rect 3329 55129 3381 55181
rect 3453 55129 3505 55181
rect 3577 55129 3629 55181
rect 3701 55129 3753 55181
rect 2833 55005 2885 55057
rect 2957 55005 3009 55057
rect 3081 55005 3133 55057
rect 3205 55005 3257 55057
rect 3329 55005 3381 55057
rect 3453 55005 3505 55057
rect 3577 55005 3629 55057
rect 3701 55005 3753 55057
rect 2833 54881 2885 54933
rect 2957 54881 3009 54933
rect 3081 54881 3133 54933
rect 3205 54881 3257 54933
rect 3329 54881 3381 54933
rect 3453 54881 3505 54933
rect 3577 54881 3629 54933
rect 3701 54881 3753 54933
rect 2833 54757 2885 54809
rect 2957 54757 3009 54809
rect 3081 54757 3133 54809
rect 3205 54757 3257 54809
rect 3329 54757 3381 54809
rect 3453 54757 3505 54809
rect 3577 54757 3629 54809
rect 3701 54757 3753 54809
rect 2833 54633 2885 54685
rect 2957 54633 3009 54685
rect 3081 54633 3133 54685
rect 3205 54633 3257 54685
rect 3329 54633 3381 54685
rect 3453 54633 3505 54685
rect 3577 54633 3629 54685
rect 3701 54633 3753 54685
rect 2833 54509 2885 54561
rect 2957 54509 3009 54561
rect 3081 54509 3133 54561
rect 3205 54509 3257 54561
rect 3329 54509 3381 54561
rect 3453 54509 3505 54561
rect 3577 54509 3629 54561
rect 3701 54509 3753 54561
rect 2833 54385 2885 54437
rect 2957 54385 3009 54437
rect 3081 54385 3133 54437
rect 3205 54385 3257 54437
rect 3329 54385 3381 54437
rect 3453 54385 3505 54437
rect 3577 54385 3629 54437
rect 3701 54385 3753 54437
rect 2833 54261 2885 54313
rect 2957 54261 3009 54313
rect 3081 54261 3133 54313
rect 3205 54261 3257 54313
rect 3329 54261 3381 54313
rect 3453 54261 3505 54313
rect 3577 54261 3629 54313
rect 3701 54261 3753 54313
rect 2833 54137 2885 54189
rect 2957 54137 3009 54189
rect 3081 54137 3133 54189
rect 3205 54137 3257 54189
rect 3329 54137 3381 54189
rect 3453 54137 3505 54189
rect 3577 54137 3629 54189
rect 3701 54137 3753 54189
rect 2833 54013 2885 54065
rect 2957 54013 3009 54065
rect 3081 54013 3133 54065
rect 3205 54013 3257 54065
rect 3329 54013 3381 54065
rect 3453 54013 3505 54065
rect 3577 54013 3629 54065
rect 3701 54013 3753 54065
rect 2833 53889 2885 53941
rect 2957 53889 3009 53941
rect 3081 53889 3133 53941
rect 3205 53889 3257 53941
rect 3329 53889 3381 53941
rect 3453 53889 3505 53941
rect 3577 53889 3629 53941
rect 3701 53889 3753 53941
rect 2833 53765 2885 53817
rect 2957 53765 3009 53817
rect 3081 53765 3133 53817
rect 3205 53765 3257 53817
rect 3329 53765 3381 53817
rect 3453 53765 3505 53817
rect 3577 53765 3629 53817
rect 3701 53765 3753 53817
rect 2833 53641 2885 53693
rect 2957 53641 3009 53693
rect 3081 53641 3133 53693
rect 3205 53641 3257 53693
rect 3329 53641 3381 53693
rect 3453 53641 3505 53693
rect 3577 53641 3629 53693
rect 3701 53641 3753 53693
rect 4340 56617 4392 56669
rect 4464 56617 4516 56669
rect 4588 56617 4640 56669
rect 4712 56617 4764 56669
rect 4340 56493 4392 56545
rect 4464 56493 4516 56545
rect 4588 56493 4640 56545
rect 4712 56493 4764 56545
rect 4340 56369 4392 56421
rect 4464 56369 4516 56421
rect 4588 56369 4640 56421
rect 4712 56369 4764 56421
rect 4340 56245 4392 56297
rect 4464 56245 4516 56297
rect 4588 56245 4640 56297
rect 4712 56245 4764 56297
rect 4340 56121 4392 56173
rect 4464 56121 4516 56173
rect 4588 56121 4640 56173
rect 4712 56121 4764 56173
rect 4340 55997 4392 56049
rect 4464 55997 4516 56049
rect 4588 55997 4640 56049
rect 4712 55997 4764 56049
rect 4340 55873 4392 55925
rect 4464 55873 4516 55925
rect 4588 55873 4640 55925
rect 4712 55873 4764 55925
rect 4340 55749 4392 55801
rect 4464 55749 4516 55801
rect 4588 55749 4640 55801
rect 4712 55749 4764 55801
rect 4340 55625 4392 55677
rect 4464 55625 4516 55677
rect 4588 55625 4640 55677
rect 4712 55625 4764 55677
rect 4340 55501 4392 55553
rect 4464 55501 4516 55553
rect 4588 55501 4640 55553
rect 4712 55501 4764 55553
rect 4340 55377 4392 55429
rect 4464 55377 4516 55429
rect 4588 55377 4640 55429
rect 4712 55377 4764 55429
rect 4340 55253 4392 55305
rect 4464 55253 4516 55305
rect 4588 55253 4640 55305
rect 4712 55253 4764 55305
rect 4340 55129 4392 55181
rect 4464 55129 4516 55181
rect 4588 55129 4640 55181
rect 4712 55129 4764 55181
rect 4340 55005 4392 55057
rect 4464 55005 4516 55057
rect 4588 55005 4640 55057
rect 4712 55005 4764 55057
rect 4340 54881 4392 54933
rect 4464 54881 4516 54933
rect 4588 54881 4640 54933
rect 4712 54881 4764 54933
rect 4340 54757 4392 54809
rect 4464 54757 4516 54809
rect 4588 54757 4640 54809
rect 4712 54757 4764 54809
rect 4340 54633 4392 54685
rect 4464 54633 4516 54685
rect 4588 54633 4640 54685
rect 4712 54633 4764 54685
rect 4340 54509 4392 54561
rect 4464 54509 4516 54561
rect 4588 54509 4640 54561
rect 4712 54509 4764 54561
rect 4340 54385 4392 54437
rect 4464 54385 4516 54437
rect 4588 54385 4640 54437
rect 4712 54385 4764 54437
rect 4340 54261 4392 54313
rect 4464 54261 4516 54313
rect 4588 54261 4640 54313
rect 4712 54261 4764 54313
rect 4340 54137 4392 54189
rect 4464 54137 4516 54189
rect 4588 54137 4640 54189
rect 4712 54137 4764 54189
rect 4340 54013 4392 54065
rect 4464 54013 4516 54065
rect 4588 54013 4640 54065
rect 4712 54013 4764 54065
rect 4340 53889 4392 53941
rect 4464 53889 4516 53941
rect 4588 53889 4640 53941
rect 4712 53889 4764 53941
rect 4340 53765 4392 53817
rect 4464 53765 4516 53817
rect 4588 53765 4640 53817
rect 4712 53765 4764 53817
rect 4340 53641 4392 53693
rect 4464 53641 4516 53693
rect 4588 53641 4640 53693
rect 4712 53641 4764 53693
rect 6297 56617 6349 56669
rect 6421 56617 6473 56669
rect 6545 56617 6597 56669
rect 6669 56617 6721 56669
rect 6793 56617 6845 56669
rect 6917 56617 6969 56669
rect 7041 56617 7093 56669
rect 6297 56493 6349 56545
rect 6421 56493 6473 56545
rect 6545 56493 6597 56545
rect 6669 56493 6721 56545
rect 6793 56493 6845 56545
rect 6917 56493 6969 56545
rect 7041 56493 7093 56545
rect 6297 56369 6349 56421
rect 6421 56369 6473 56421
rect 6545 56369 6597 56421
rect 6669 56369 6721 56421
rect 6793 56369 6845 56421
rect 6917 56369 6969 56421
rect 7041 56369 7093 56421
rect 6297 56245 6349 56297
rect 6421 56245 6473 56297
rect 6545 56245 6597 56297
rect 6669 56245 6721 56297
rect 6793 56245 6845 56297
rect 6917 56245 6969 56297
rect 7041 56245 7093 56297
rect 6297 56121 6349 56173
rect 6421 56121 6473 56173
rect 6545 56121 6597 56173
rect 6669 56121 6721 56173
rect 6793 56121 6845 56173
rect 6917 56121 6969 56173
rect 7041 56121 7093 56173
rect 6297 55997 6349 56049
rect 6421 55997 6473 56049
rect 6545 55997 6597 56049
rect 6669 55997 6721 56049
rect 6793 55997 6845 56049
rect 6917 55997 6969 56049
rect 7041 55997 7093 56049
rect 6297 55873 6349 55925
rect 6421 55873 6473 55925
rect 6545 55873 6597 55925
rect 6669 55873 6721 55925
rect 6793 55873 6845 55925
rect 6917 55873 6969 55925
rect 7041 55873 7093 55925
rect 6297 55749 6349 55801
rect 6421 55749 6473 55801
rect 6545 55749 6597 55801
rect 6669 55749 6721 55801
rect 6793 55749 6845 55801
rect 6917 55749 6969 55801
rect 7041 55749 7093 55801
rect 6297 55625 6349 55677
rect 6421 55625 6473 55677
rect 6545 55625 6597 55677
rect 6669 55625 6721 55677
rect 6793 55625 6845 55677
rect 6917 55625 6969 55677
rect 7041 55625 7093 55677
rect 6297 55501 6349 55553
rect 6421 55501 6473 55553
rect 6545 55501 6597 55553
rect 6669 55501 6721 55553
rect 6793 55501 6845 55553
rect 6917 55501 6969 55553
rect 7041 55501 7093 55553
rect 6297 55377 6349 55429
rect 6421 55377 6473 55429
rect 6545 55377 6597 55429
rect 6669 55377 6721 55429
rect 6793 55377 6845 55429
rect 6917 55377 6969 55429
rect 7041 55377 7093 55429
rect 6297 55253 6349 55305
rect 6421 55253 6473 55305
rect 6545 55253 6597 55305
rect 6669 55253 6721 55305
rect 6793 55253 6845 55305
rect 6917 55253 6969 55305
rect 7041 55253 7093 55305
rect 6297 55129 6349 55181
rect 6421 55129 6473 55181
rect 6545 55129 6597 55181
rect 6669 55129 6721 55181
rect 6793 55129 6845 55181
rect 6917 55129 6969 55181
rect 7041 55129 7093 55181
rect 6297 55005 6349 55057
rect 6421 55005 6473 55057
rect 6545 55005 6597 55057
rect 6669 55005 6721 55057
rect 6793 55005 6845 55057
rect 6917 55005 6969 55057
rect 7041 55005 7093 55057
rect 6297 54881 6349 54933
rect 6421 54881 6473 54933
rect 6545 54881 6597 54933
rect 6669 54881 6721 54933
rect 6793 54881 6845 54933
rect 6917 54881 6969 54933
rect 7041 54881 7093 54933
rect 6297 54757 6349 54809
rect 6421 54757 6473 54809
rect 6545 54757 6597 54809
rect 6669 54757 6721 54809
rect 6793 54757 6845 54809
rect 6917 54757 6969 54809
rect 7041 54757 7093 54809
rect 6297 54633 6349 54685
rect 6421 54633 6473 54685
rect 6545 54633 6597 54685
rect 6669 54633 6721 54685
rect 6793 54633 6845 54685
rect 6917 54633 6969 54685
rect 7041 54633 7093 54685
rect 6297 54509 6349 54561
rect 6421 54509 6473 54561
rect 6545 54509 6597 54561
rect 6669 54509 6721 54561
rect 6793 54509 6845 54561
rect 6917 54509 6969 54561
rect 7041 54509 7093 54561
rect 6297 54385 6349 54437
rect 6421 54385 6473 54437
rect 6545 54385 6597 54437
rect 6669 54385 6721 54437
rect 6793 54385 6845 54437
rect 6917 54385 6969 54437
rect 7041 54385 7093 54437
rect 6297 54261 6349 54313
rect 6421 54261 6473 54313
rect 6545 54261 6597 54313
rect 6669 54261 6721 54313
rect 6793 54261 6845 54313
rect 6917 54261 6969 54313
rect 7041 54261 7093 54313
rect 6297 54137 6349 54189
rect 6421 54137 6473 54189
rect 6545 54137 6597 54189
rect 6669 54137 6721 54189
rect 6793 54137 6845 54189
rect 6917 54137 6969 54189
rect 7041 54137 7093 54189
rect 6297 54013 6349 54065
rect 6421 54013 6473 54065
rect 6545 54013 6597 54065
rect 6669 54013 6721 54065
rect 6793 54013 6845 54065
rect 6917 54013 6969 54065
rect 7041 54013 7093 54065
rect 6297 53889 6349 53941
rect 6421 53889 6473 53941
rect 6545 53889 6597 53941
rect 6669 53889 6721 53941
rect 6793 53889 6845 53941
rect 6917 53889 6969 53941
rect 7041 53889 7093 53941
rect 6297 53765 6349 53817
rect 6421 53765 6473 53817
rect 6545 53765 6597 53817
rect 6669 53765 6721 53817
rect 6793 53765 6845 53817
rect 6917 53765 6969 53817
rect 7041 53765 7093 53817
rect 6297 53641 6349 53693
rect 6421 53641 6473 53693
rect 6545 53641 6597 53693
rect 6669 53641 6721 53693
rect 6793 53641 6845 53693
rect 6917 53641 6969 53693
rect 7041 53641 7093 53693
rect 7885 56617 7937 56669
rect 8009 56617 8061 56669
rect 8133 56617 8185 56669
rect 8257 56617 8309 56669
rect 8381 56617 8433 56669
rect 8505 56617 8557 56669
rect 8629 56617 8681 56669
rect 7885 56493 7937 56545
rect 8009 56493 8061 56545
rect 8133 56493 8185 56545
rect 8257 56493 8309 56545
rect 8381 56493 8433 56545
rect 8505 56493 8557 56545
rect 8629 56493 8681 56545
rect 7885 56369 7937 56421
rect 8009 56369 8061 56421
rect 8133 56369 8185 56421
rect 8257 56369 8309 56421
rect 8381 56369 8433 56421
rect 8505 56369 8557 56421
rect 8629 56369 8681 56421
rect 7885 56245 7937 56297
rect 8009 56245 8061 56297
rect 8133 56245 8185 56297
rect 8257 56245 8309 56297
rect 8381 56245 8433 56297
rect 8505 56245 8557 56297
rect 8629 56245 8681 56297
rect 7885 56121 7937 56173
rect 8009 56121 8061 56173
rect 8133 56121 8185 56173
rect 8257 56121 8309 56173
rect 8381 56121 8433 56173
rect 8505 56121 8557 56173
rect 8629 56121 8681 56173
rect 7885 55997 7937 56049
rect 8009 55997 8061 56049
rect 8133 55997 8185 56049
rect 8257 55997 8309 56049
rect 8381 55997 8433 56049
rect 8505 55997 8557 56049
rect 8629 55997 8681 56049
rect 7885 55873 7937 55925
rect 8009 55873 8061 55925
rect 8133 55873 8185 55925
rect 8257 55873 8309 55925
rect 8381 55873 8433 55925
rect 8505 55873 8557 55925
rect 8629 55873 8681 55925
rect 7885 55749 7937 55801
rect 8009 55749 8061 55801
rect 8133 55749 8185 55801
rect 8257 55749 8309 55801
rect 8381 55749 8433 55801
rect 8505 55749 8557 55801
rect 8629 55749 8681 55801
rect 7885 55625 7937 55677
rect 8009 55625 8061 55677
rect 8133 55625 8185 55677
rect 8257 55625 8309 55677
rect 8381 55625 8433 55677
rect 8505 55625 8557 55677
rect 8629 55625 8681 55677
rect 7885 55501 7937 55553
rect 8009 55501 8061 55553
rect 8133 55501 8185 55553
rect 8257 55501 8309 55553
rect 8381 55501 8433 55553
rect 8505 55501 8557 55553
rect 8629 55501 8681 55553
rect 7885 55377 7937 55429
rect 8009 55377 8061 55429
rect 8133 55377 8185 55429
rect 8257 55377 8309 55429
rect 8381 55377 8433 55429
rect 8505 55377 8557 55429
rect 8629 55377 8681 55429
rect 7885 55253 7937 55305
rect 8009 55253 8061 55305
rect 8133 55253 8185 55305
rect 8257 55253 8309 55305
rect 8381 55253 8433 55305
rect 8505 55253 8557 55305
rect 8629 55253 8681 55305
rect 7885 55129 7937 55181
rect 8009 55129 8061 55181
rect 8133 55129 8185 55181
rect 8257 55129 8309 55181
rect 8381 55129 8433 55181
rect 8505 55129 8557 55181
rect 8629 55129 8681 55181
rect 7885 55005 7937 55057
rect 8009 55005 8061 55057
rect 8133 55005 8185 55057
rect 8257 55005 8309 55057
rect 8381 55005 8433 55057
rect 8505 55005 8557 55057
rect 8629 55005 8681 55057
rect 7885 54881 7937 54933
rect 8009 54881 8061 54933
rect 8133 54881 8185 54933
rect 8257 54881 8309 54933
rect 8381 54881 8433 54933
rect 8505 54881 8557 54933
rect 8629 54881 8681 54933
rect 7885 54757 7937 54809
rect 8009 54757 8061 54809
rect 8133 54757 8185 54809
rect 8257 54757 8309 54809
rect 8381 54757 8433 54809
rect 8505 54757 8557 54809
rect 8629 54757 8681 54809
rect 7885 54633 7937 54685
rect 8009 54633 8061 54685
rect 8133 54633 8185 54685
rect 8257 54633 8309 54685
rect 8381 54633 8433 54685
rect 8505 54633 8557 54685
rect 8629 54633 8681 54685
rect 7885 54509 7937 54561
rect 8009 54509 8061 54561
rect 8133 54509 8185 54561
rect 8257 54509 8309 54561
rect 8381 54509 8433 54561
rect 8505 54509 8557 54561
rect 8629 54509 8681 54561
rect 7885 54385 7937 54437
rect 8009 54385 8061 54437
rect 8133 54385 8185 54437
rect 8257 54385 8309 54437
rect 8381 54385 8433 54437
rect 8505 54385 8557 54437
rect 8629 54385 8681 54437
rect 7885 54261 7937 54313
rect 8009 54261 8061 54313
rect 8133 54261 8185 54313
rect 8257 54261 8309 54313
rect 8381 54261 8433 54313
rect 8505 54261 8557 54313
rect 8629 54261 8681 54313
rect 7885 54137 7937 54189
rect 8009 54137 8061 54189
rect 8133 54137 8185 54189
rect 8257 54137 8309 54189
rect 8381 54137 8433 54189
rect 8505 54137 8557 54189
rect 8629 54137 8681 54189
rect 7885 54013 7937 54065
rect 8009 54013 8061 54065
rect 8133 54013 8185 54065
rect 8257 54013 8309 54065
rect 8381 54013 8433 54065
rect 8505 54013 8557 54065
rect 8629 54013 8681 54065
rect 7885 53889 7937 53941
rect 8009 53889 8061 53941
rect 8133 53889 8185 53941
rect 8257 53889 8309 53941
rect 8381 53889 8433 53941
rect 8505 53889 8557 53941
rect 8629 53889 8681 53941
rect 7885 53765 7937 53817
rect 8009 53765 8061 53817
rect 8133 53765 8185 53817
rect 8257 53765 8309 53817
rect 8381 53765 8433 53817
rect 8505 53765 8557 53817
rect 8629 53765 8681 53817
rect 7885 53641 7937 53693
rect 8009 53641 8061 53693
rect 8133 53641 8185 53693
rect 8257 53641 8309 53693
rect 8381 53641 8433 53693
rect 8505 53641 8557 53693
rect 8629 53641 8681 53693
rect 10214 56617 10266 56669
rect 10338 56617 10390 56669
rect 10462 56617 10514 56669
rect 10586 56617 10638 56669
rect 10214 56493 10266 56545
rect 10338 56493 10390 56545
rect 10462 56493 10514 56545
rect 10586 56493 10638 56545
rect 10214 56369 10266 56421
rect 10338 56369 10390 56421
rect 10462 56369 10514 56421
rect 10586 56369 10638 56421
rect 10214 56245 10266 56297
rect 10338 56245 10390 56297
rect 10462 56245 10514 56297
rect 10586 56245 10638 56297
rect 10214 56121 10266 56173
rect 10338 56121 10390 56173
rect 10462 56121 10514 56173
rect 10586 56121 10638 56173
rect 10214 55997 10266 56049
rect 10338 55997 10390 56049
rect 10462 55997 10514 56049
rect 10586 55997 10638 56049
rect 10214 55873 10266 55925
rect 10338 55873 10390 55925
rect 10462 55873 10514 55925
rect 10586 55873 10638 55925
rect 10214 55749 10266 55801
rect 10338 55749 10390 55801
rect 10462 55749 10514 55801
rect 10586 55749 10638 55801
rect 10214 55625 10266 55677
rect 10338 55625 10390 55677
rect 10462 55625 10514 55677
rect 10586 55625 10638 55677
rect 10214 55501 10266 55553
rect 10338 55501 10390 55553
rect 10462 55501 10514 55553
rect 10586 55501 10638 55553
rect 10214 55377 10266 55429
rect 10338 55377 10390 55429
rect 10462 55377 10514 55429
rect 10586 55377 10638 55429
rect 10214 55253 10266 55305
rect 10338 55253 10390 55305
rect 10462 55253 10514 55305
rect 10586 55253 10638 55305
rect 10214 55129 10266 55181
rect 10338 55129 10390 55181
rect 10462 55129 10514 55181
rect 10586 55129 10638 55181
rect 10214 55005 10266 55057
rect 10338 55005 10390 55057
rect 10462 55005 10514 55057
rect 10586 55005 10638 55057
rect 10214 54881 10266 54933
rect 10338 54881 10390 54933
rect 10462 54881 10514 54933
rect 10586 54881 10638 54933
rect 10214 54757 10266 54809
rect 10338 54757 10390 54809
rect 10462 54757 10514 54809
rect 10586 54757 10638 54809
rect 10214 54633 10266 54685
rect 10338 54633 10390 54685
rect 10462 54633 10514 54685
rect 10586 54633 10638 54685
rect 10214 54509 10266 54561
rect 10338 54509 10390 54561
rect 10462 54509 10514 54561
rect 10586 54509 10638 54561
rect 10214 54385 10266 54437
rect 10338 54385 10390 54437
rect 10462 54385 10514 54437
rect 10586 54385 10638 54437
rect 10214 54261 10266 54313
rect 10338 54261 10390 54313
rect 10462 54261 10514 54313
rect 10586 54261 10638 54313
rect 10214 54137 10266 54189
rect 10338 54137 10390 54189
rect 10462 54137 10514 54189
rect 10586 54137 10638 54189
rect 10214 54013 10266 54065
rect 10338 54013 10390 54065
rect 10462 54013 10514 54065
rect 10586 54013 10638 54065
rect 10214 53889 10266 53941
rect 10338 53889 10390 53941
rect 10462 53889 10514 53941
rect 10586 53889 10638 53941
rect 10214 53765 10266 53817
rect 10338 53765 10390 53817
rect 10462 53765 10514 53817
rect 10586 53765 10638 53817
rect 10214 53641 10266 53693
rect 10338 53641 10390 53693
rect 10462 53641 10514 53693
rect 10586 53641 10638 53693
rect 11225 56617 11277 56669
rect 11349 56617 11401 56669
rect 11473 56617 11525 56669
rect 11597 56617 11649 56669
rect 11721 56617 11773 56669
rect 11845 56617 11897 56669
rect 11969 56617 12021 56669
rect 12093 56617 12145 56669
rect 11225 56493 11277 56545
rect 11349 56493 11401 56545
rect 11473 56493 11525 56545
rect 11597 56493 11649 56545
rect 11721 56493 11773 56545
rect 11845 56493 11897 56545
rect 11969 56493 12021 56545
rect 12093 56493 12145 56545
rect 11225 56369 11277 56421
rect 11349 56369 11401 56421
rect 11473 56369 11525 56421
rect 11597 56369 11649 56421
rect 11721 56369 11773 56421
rect 11845 56369 11897 56421
rect 11969 56369 12021 56421
rect 12093 56369 12145 56421
rect 11225 56245 11277 56297
rect 11349 56245 11401 56297
rect 11473 56245 11525 56297
rect 11597 56245 11649 56297
rect 11721 56245 11773 56297
rect 11845 56245 11897 56297
rect 11969 56245 12021 56297
rect 12093 56245 12145 56297
rect 11225 56121 11277 56173
rect 11349 56121 11401 56173
rect 11473 56121 11525 56173
rect 11597 56121 11649 56173
rect 11721 56121 11773 56173
rect 11845 56121 11897 56173
rect 11969 56121 12021 56173
rect 12093 56121 12145 56173
rect 11225 55997 11277 56049
rect 11349 55997 11401 56049
rect 11473 55997 11525 56049
rect 11597 55997 11649 56049
rect 11721 55997 11773 56049
rect 11845 55997 11897 56049
rect 11969 55997 12021 56049
rect 12093 55997 12145 56049
rect 11225 55873 11277 55925
rect 11349 55873 11401 55925
rect 11473 55873 11525 55925
rect 11597 55873 11649 55925
rect 11721 55873 11773 55925
rect 11845 55873 11897 55925
rect 11969 55873 12021 55925
rect 12093 55873 12145 55925
rect 11225 55749 11277 55801
rect 11349 55749 11401 55801
rect 11473 55749 11525 55801
rect 11597 55749 11649 55801
rect 11721 55749 11773 55801
rect 11845 55749 11897 55801
rect 11969 55749 12021 55801
rect 12093 55749 12145 55801
rect 11225 55625 11277 55677
rect 11349 55625 11401 55677
rect 11473 55625 11525 55677
rect 11597 55625 11649 55677
rect 11721 55625 11773 55677
rect 11845 55625 11897 55677
rect 11969 55625 12021 55677
rect 12093 55625 12145 55677
rect 11225 55501 11277 55553
rect 11349 55501 11401 55553
rect 11473 55501 11525 55553
rect 11597 55501 11649 55553
rect 11721 55501 11773 55553
rect 11845 55501 11897 55553
rect 11969 55501 12021 55553
rect 12093 55501 12145 55553
rect 11225 55377 11277 55429
rect 11349 55377 11401 55429
rect 11473 55377 11525 55429
rect 11597 55377 11649 55429
rect 11721 55377 11773 55429
rect 11845 55377 11897 55429
rect 11969 55377 12021 55429
rect 12093 55377 12145 55429
rect 11225 55253 11277 55305
rect 11349 55253 11401 55305
rect 11473 55253 11525 55305
rect 11597 55253 11649 55305
rect 11721 55253 11773 55305
rect 11845 55253 11897 55305
rect 11969 55253 12021 55305
rect 12093 55253 12145 55305
rect 11225 55129 11277 55181
rect 11349 55129 11401 55181
rect 11473 55129 11525 55181
rect 11597 55129 11649 55181
rect 11721 55129 11773 55181
rect 11845 55129 11897 55181
rect 11969 55129 12021 55181
rect 12093 55129 12145 55181
rect 11225 55005 11277 55057
rect 11349 55005 11401 55057
rect 11473 55005 11525 55057
rect 11597 55005 11649 55057
rect 11721 55005 11773 55057
rect 11845 55005 11897 55057
rect 11969 55005 12021 55057
rect 12093 55005 12145 55057
rect 11225 54881 11277 54933
rect 11349 54881 11401 54933
rect 11473 54881 11525 54933
rect 11597 54881 11649 54933
rect 11721 54881 11773 54933
rect 11845 54881 11897 54933
rect 11969 54881 12021 54933
rect 12093 54881 12145 54933
rect 11225 54757 11277 54809
rect 11349 54757 11401 54809
rect 11473 54757 11525 54809
rect 11597 54757 11649 54809
rect 11721 54757 11773 54809
rect 11845 54757 11897 54809
rect 11969 54757 12021 54809
rect 12093 54757 12145 54809
rect 11225 54633 11277 54685
rect 11349 54633 11401 54685
rect 11473 54633 11525 54685
rect 11597 54633 11649 54685
rect 11721 54633 11773 54685
rect 11845 54633 11897 54685
rect 11969 54633 12021 54685
rect 12093 54633 12145 54685
rect 11225 54509 11277 54561
rect 11349 54509 11401 54561
rect 11473 54509 11525 54561
rect 11597 54509 11649 54561
rect 11721 54509 11773 54561
rect 11845 54509 11897 54561
rect 11969 54509 12021 54561
rect 12093 54509 12145 54561
rect 11225 54385 11277 54437
rect 11349 54385 11401 54437
rect 11473 54385 11525 54437
rect 11597 54385 11649 54437
rect 11721 54385 11773 54437
rect 11845 54385 11897 54437
rect 11969 54385 12021 54437
rect 12093 54385 12145 54437
rect 11225 54261 11277 54313
rect 11349 54261 11401 54313
rect 11473 54261 11525 54313
rect 11597 54261 11649 54313
rect 11721 54261 11773 54313
rect 11845 54261 11897 54313
rect 11969 54261 12021 54313
rect 12093 54261 12145 54313
rect 11225 54137 11277 54189
rect 11349 54137 11401 54189
rect 11473 54137 11525 54189
rect 11597 54137 11649 54189
rect 11721 54137 11773 54189
rect 11845 54137 11897 54189
rect 11969 54137 12021 54189
rect 12093 54137 12145 54189
rect 11225 54013 11277 54065
rect 11349 54013 11401 54065
rect 11473 54013 11525 54065
rect 11597 54013 11649 54065
rect 11721 54013 11773 54065
rect 11845 54013 11897 54065
rect 11969 54013 12021 54065
rect 12093 54013 12145 54065
rect 11225 53889 11277 53941
rect 11349 53889 11401 53941
rect 11473 53889 11525 53941
rect 11597 53889 11649 53941
rect 11721 53889 11773 53941
rect 11845 53889 11897 53941
rect 11969 53889 12021 53941
rect 12093 53889 12145 53941
rect 11225 53765 11277 53817
rect 11349 53765 11401 53817
rect 11473 53765 11525 53817
rect 11597 53765 11649 53817
rect 11721 53765 11773 53817
rect 11845 53765 11897 53817
rect 11969 53765 12021 53817
rect 12093 53765 12145 53817
rect 11225 53641 11277 53693
rect 11349 53641 11401 53693
rect 11473 53641 11525 53693
rect 11597 53641 11649 53693
rect 11721 53641 11773 53693
rect 11845 53641 11897 53693
rect 11969 53641 12021 53693
rect 12093 53641 12145 53693
rect 13141 56617 13193 56669
rect 13265 56617 13317 56669
rect 13389 56617 13441 56669
rect 13513 56617 13565 56669
rect 13637 56617 13689 56669
rect 13761 56617 13813 56669
rect 13885 56617 13937 56669
rect 14009 56617 14061 56669
rect 13141 56493 13193 56545
rect 13265 56493 13317 56545
rect 13389 56493 13441 56545
rect 13513 56493 13565 56545
rect 13637 56493 13689 56545
rect 13761 56493 13813 56545
rect 13885 56493 13937 56545
rect 14009 56493 14061 56545
rect 13141 56369 13193 56421
rect 13265 56369 13317 56421
rect 13389 56369 13441 56421
rect 13513 56369 13565 56421
rect 13637 56369 13689 56421
rect 13761 56369 13813 56421
rect 13885 56369 13937 56421
rect 14009 56369 14061 56421
rect 13141 56245 13193 56297
rect 13265 56245 13317 56297
rect 13389 56245 13441 56297
rect 13513 56245 13565 56297
rect 13637 56245 13689 56297
rect 13761 56245 13813 56297
rect 13885 56245 13937 56297
rect 14009 56245 14061 56297
rect 13141 56121 13193 56173
rect 13265 56121 13317 56173
rect 13389 56121 13441 56173
rect 13513 56121 13565 56173
rect 13637 56121 13689 56173
rect 13761 56121 13813 56173
rect 13885 56121 13937 56173
rect 14009 56121 14061 56173
rect 13141 55997 13193 56049
rect 13265 55997 13317 56049
rect 13389 55997 13441 56049
rect 13513 55997 13565 56049
rect 13637 55997 13689 56049
rect 13761 55997 13813 56049
rect 13885 55997 13937 56049
rect 14009 55997 14061 56049
rect 13141 55873 13193 55925
rect 13265 55873 13317 55925
rect 13389 55873 13441 55925
rect 13513 55873 13565 55925
rect 13637 55873 13689 55925
rect 13761 55873 13813 55925
rect 13885 55873 13937 55925
rect 14009 55873 14061 55925
rect 13141 55749 13193 55801
rect 13265 55749 13317 55801
rect 13389 55749 13441 55801
rect 13513 55749 13565 55801
rect 13637 55749 13689 55801
rect 13761 55749 13813 55801
rect 13885 55749 13937 55801
rect 14009 55749 14061 55801
rect 13141 55625 13193 55677
rect 13265 55625 13317 55677
rect 13389 55625 13441 55677
rect 13513 55625 13565 55677
rect 13637 55625 13689 55677
rect 13761 55625 13813 55677
rect 13885 55625 13937 55677
rect 14009 55625 14061 55677
rect 13141 55501 13193 55553
rect 13265 55501 13317 55553
rect 13389 55501 13441 55553
rect 13513 55501 13565 55553
rect 13637 55501 13689 55553
rect 13761 55501 13813 55553
rect 13885 55501 13937 55553
rect 14009 55501 14061 55553
rect 13141 55377 13193 55429
rect 13265 55377 13317 55429
rect 13389 55377 13441 55429
rect 13513 55377 13565 55429
rect 13637 55377 13689 55429
rect 13761 55377 13813 55429
rect 13885 55377 13937 55429
rect 14009 55377 14061 55429
rect 13141 55253 13193 55305
rect 13265 55253 13317 55305
rect 13389 55253 13441 55305
rect 13513 55253 13565 55305
rect 13637 55253 13689 55305
rect 13761 55253 13813 55305
rect 13885 55253 13937 55305
rect 14009 55253 14061 55305
rect 13141 55129 13193 55181
rect 13265 55129 13317 55181
rect 13389 55129 13441 55181
rect 13513 55129 13565 55181
rect 13637 55129 13689 55181
rect 13761 55129 13813 55181
rect 13885 55129 13937 55181
rect 14009 55129 14061 55181
rect 13141 55005 13193 55057
rect 13265 55005 13317 55057
rect 13389 55005 13441 55057
rect 13513 55005 13565 55057
rect 13637 55005 13689 55057
rect 13761 55005 13813 55057
rect 13885 55005 13937 55057
rect 14009 55005 14061 55057
rect 13141 54881 13193 54933
rect 13265 54881 13317 54933
rect 13389 54881 13441 54933
rect 13513 54881 13565 54933
rect 13637 54881 13689 54933
rect 13761 54881 13813 54933
rect 13885 54881 13937 54933
rect 14009 54881 14061 54933
rect 13141 54757 13193 54809
rect 13265 54757 13317 54809
rect 13389 54757 13441 54809
rect 13513 54757 13565 54809
rect 13637 54757 13689 54809
rect 13761 54757 13813 54809
rect 13885 54757 13937 54809
rect 14009 54757 14061 54809
rect 13141 54633 13193 54685
rect 13265 54633 13317 54685
rect 13389 54633 13441 54685
rect 13513 54633 13565 54685
rect 13637 54633 13689 54685
rect 13761 54633 13813 54685
rect 13885 54633 13937 54685
rect 14009 54633 14061 54685
rect 13141 54509 13193 54561
rect 13265 54509 13317 54561
rect 13389 54509 13441 54561
rect 13513 54509 13565 54561
rect 13637 54509 13689 54561
rect 13761 54509 13813 54561
rect 13885 54509 13937 54561
rect 14009 54509 14061 54561
rect 13141 54385 13193 54437
rect 13265 54385 13317 54437
rect 13389 54385 13441 54437
rect 13513 54385 13565 54437
rect 13637 54385 13689 54437
rect 13761 54385 13813 54437
rect 13885 54385 13937 54437
rect 14009 54385 14061 54437
rect 13141 54261 13193 54313
rect 13265 54261 13317 54313
rect 13389 54261 13441 54313
rect 13513 54261 13565 54313
rect 13637 54261 13689 54313
rect 13761 54261 13813 54313
rect 13885 54261 13937 54313
rect 14009 54261 14061 54313
rect 13141 54137 13193 54189
rect 13265 54137 13317 54189
rect 13389 54137 13441 54189
rect 13513 54137 13565 54189
rect 13637 54137 13689 54189
rect 13761 54137 13813 54189
rect 13885 54137 13937 54189
rect 14009 54137 14061 54189
rect 13141 54013 13193 54065
rect 13265 54013 13317 54065
rect 13389 54013 13441 54065
rect 13513 54013 13565 54065
rect 13637 54013 13689 54065
rect 13761 54013 13813 54065
rect 13885 54013 13937 54065
rect 14009 54013 14061 54065
rect 13141 53889 13193 53941
rect 13265 53889 13317 53941
rect 13389 53889 13441 53941
rect 13513 53889 13565 53941
rect 13637 53889 13689 53941
rect 13761 53889 13813 53941
rect 13885 53889 13937 53941
rect 14009 53889 14061 53941
rect 13141 53765 13193 53817
rect 13265 53765 13317 53817
rect 13389 53765 13441 53817
rect 13513 53765 13565 53817
rect 13637 53765 13689 53817
rect 13761 53765 13813 53817
rect 13885 53765 13937 53817
rect 14009 53765 14061 53817
rect 13141 53641 13193 53693
rect 13265 53641 13317 53693
rect 13389 53641 13441 53693
rect 13513 53641 13565 53693
rect 13637 53641 13689 53693
rect 13761 53641 13813 53693
rect 13885 53641 13937 53693
rect 14009 53641 14061 53693
rect 2501 53432 2553 53484
rect 2609 53432 2661 53484
rect 4871 53432 4923 53484
rect 4979 53432 5031 53484
rect 7247 53432 7299 53484
rect 7355 53432 7407 53484
rect 7463 53432 7515 53484
rect 7571 53432 7623 53484
rect 7679 53432 7731 53484
rect 9947 53432 9999 53484
rect 10055 53432 10107 53484
rect 12317 53432 12369 53484
rect 12425 53432 12477 53484
rect 2501 53324 2553 53376
rect 2609 53324 2661 53376
rect 4871 53324 4923 53376
rect 4979 53324 5031 53376
rect 7247 53324 7299 53376
rect 7355 53324 7407 53376
rect 7463 53324 7515 53376
rect 7571 53324 7623 53376
rect 7679 53324 7731 53376
rect 9947 53324 9999 53376
rect 10055 53324 10107 53376
rect 12317 53324 12369 53376
rect 12425 53324 12477 53376
rect 2501 53251 2553 53268
rect 2609 53251 2661 53268
rect 4871 53251 4923 53268
rect 4979 53251 5031 53268
rect 7247 53251 7299 53268
rect 7355 53251 7407 53268
rect 7463 53251 7515 53268
rect 7571 53251 7623 53268
rect 7679 53251 7731 53268
rect 9947 53251 9999 53268
rect 10055 53251 10107 53268
rect 12317 53251 12369 53268
rect 12425 53251 12477 53268
rect 2501 53216 2553 53251
rect 2609 53216 2661 53251
rect 4871 53216 4923 53251
rect 4979 53216 5031 53251
rect 7247 53216 7299 53251
rect 7355 53216 7407 53251
rect 7463 53216 7515 53251
rect 7571 53216 7623 53251
rect 7679 53216 7731 53251
rect 9947 53216 9999 53251
rect 10055 53216 10107 53251
rect 12317 53216 12369 53251
rect 12425 53216 12477 53251
rect 22 52522 74 52574
rect 22 52414 74 52466
rect 22 52306 74 52358
rect 22 52198 74 52250
rect 22 52090 74 52142
rect 22 51982 74 52034
rect 22 51874 74 51926
rect 22 51766 74 51818
rect 22 51658 74 51710
rect 22 51550 74 51602
rect 22 51442 74 51494
rect 22 51334 74 51386
rect 22 51226 74 51278
rect 2810 52536 2862 52588
rect 2934 52536 2986 52588
rect 3058 52536 3110 52588
rect 3182 52536 3234 52588
rect 3306 52536 3358 52588
rect 3430 52536 3482 52588
rect 3554 52536 3606 52588
rect 3678 52536 3730 52588
rect 3802 52536 3854 52588
rect 3926 52536 3978 52588
rect 4050 52536 4102 52588
rect 4174 52536 4226 52588
rect 4298 52536 4350 52588
rect 4422 52536 4474 52588
rect 4546 52536 4598 52588
rect 4670 52536 4722 52588
rect 5180 52536 5232 52588
rect 5304 52536 5356 52588
rect 5428 52536 5480 52588
rect 5552 52536 5604 52588
rect 5676 52536 5728 52588
rect 5800 52536 5852 52588
rect 5924 52536 5976 52588
rect 6048 52536 6100 52588
rect 6172 52536 6224 52588
rect 6296 52536 6348 52588
rect 6420 52536 6472 52588
rect 6544 52536 6596 52588
rect 6668 52536 6720 52588
rect 6792 52536 6844 52588
rect 6916 52536 6968 52588
rect 7040 52536 7092 52588
rect 7886 52536 7938 52588
rect 8010 52536 8062 52588
rect 8134 52536 8186 52588
rect 8258 52536 8310 52588
rect 8382 52536 8434 52588
rect 8506 52536 8558 52588
rect 8630 52536 8682 52588
rect 8754 52536 8806 52588
rect 8878 52536 8930 52588
rect 9002 52536 9054 52588
rect 9126 52536 9178 52588
rect 9250 52536 9302 52588
rect 9374 52536 9426 52588
rect 9498 52536 9550 52588
rect 9622 52536 9674 52588
rect 9746 52536 9798 52588
rect 10256 52536 10308 52588
rect 10380 52536 10432 52588
rect 10504 52536 10556 52588
rect 10628 52536 10680 52588
rect 10752 52536 10804 52588
rect 10876 52536 10928 52588
rect 11000 52536 11052 52588
rect 11124 52536 11176 52588
rect 11248 52536 11300 52588
rect 11372 52536 11424 52588
rect 11496 52536 11548 52588
rect 11620 52536 11672 52588
rect 11744 52536 11796 52588
rect 11868 52536 11920 52588
rect 11992 52536 12044 52588
rect 12116 52536 12168 52588
rect 2810 52412 2862 52464
rect 2934 52412 2986 52464
rect 3058 52412 3110 52464
rect 3182 52412 3234 52464
rect 3306 52412 3358 52464
rect 3430 52412 3482 52464
rect 3554 52412 3606 52464
rect 3678 52412 3730 52464
rect 3802 52412 3854 52464
rect 3926 52412 3978 52464
rect 4050 52412 4102 52464
rect 4174 52412 4226 52464
rect 4298 52412 4350 52464
rect 4422 52412 4474 52464
rect 4546 52412 4598 52464
rect 4670 52412 4722 52464
rect 5180 52412 5232 52464
rect 5304 52412 5356 52464
rect 5428 52412 5480 52464
rect 5552 52412 5604 52464
rect 5676 52412 5728 52464
rect 5800 52412 5852 52464
rect 5924 52412 5976 52464
rect 6048 52412 6100 52464
rect 6172 52412 6224 52464
rect 6296 52412 6348 52464
rect 6420 52412 6472 52464
rect 6544 52412 6596 52464
rect 6668 52412 6720 52464
rect 6792 52412 6844 52464
rect 6916 52412 6968 52464
rect 7040 52412 7092 52464
rect 7886 52412 7938 52464
rect 8010 52412 8062 52464
rect 8134 52412 8186 52464
rect 8258 52412 8310 52464
rect 8382 52412 8434 52464
rect 8506 52412 8558 52464
rect 8630 52412 8682 52464
rect 8754 52412 8806 52464
rect 8878 52412 8930 52464
rect 9002 52412 9054 52464
rect 9126 52412 9178 52464
rect 9250 52412 9302 52464
rect 9374 52412 9426 52464
rect 9498 52412 9550 52464
rect 9622 52412 9674 52464
rect 9746 52412 9798 52464
rect 10256 52412 10308 52464
rect 10380 52412 10432 52464
rect 10504 52412 10556 52464
rect 10628 52412 10680 52464
rect 10752 52412 10804 52464
rect 10876 52412 10928 52464
rect 11000 52412 11052 52464
rect 11124 52412 11176 52464
rect 11248 52412 11300 52464
rect 11372 52412 11424 52464
rect 11496 52412 11548 52464
rect 11620 52412 11672 52464
rect 11744 52412 11796 52464
rect 11868 52412 11920 52464
rect 11992 52412 12044 52464
rect 12116 52412 12168 52464
rect 2810 52288 2862 52340
rect 2934 52288 2986 52340
rect 3058 52288 3110 52340
rect 3182 52288 3234 52340
rect 3306 52288 3358 52340
rect 3430 52288 3482 52340
rect 3554 52288 3606 52340
rect 3678 52288 3730 52340
rect 3802 52288 3854 52340
rect 3926 52288 3978 52340
rect 4050 52288 4102 52340
rect 4174 52288 4226 52340
rect 4298 52288 4350 52340
rect 4422 52288 4474 52340
rect 4546 52288 4598 52340
rect 4670 52288 4722 52340
rect 5180 52288 5232 52340
rect 5304 52288 5356 52340
rect 5428 52288 5480 52340
rect 5552 52288 5604 52340
rect 5676 52288 5728 52340
rect 5800 52288 5852 52340
rect 5924 52288 5976 52340
rect 6048 52288 6100 52340
rect 6172 52288 6224 52340
rect 6296 52288 6348 52340
rect 6420 52288 6472 52340
rect 6544 52288 6596 52340
rect 6668 52288 6720 52340
rect 6792 52288 6844 52340
rect 6916 52288 6968 52340
rect 7040 52288 7092 52340
rect 7886 52288 7938 52340
rect 8010 52288 8062 52340
rect 8134 52288 8186 52340
rect 8258 52288 8310 52340
rect 8382 52288 8434 52340
rect 8506 52288 8558 52340
rect 8630 52288 8682 52340
rect 8754 52288 8806 52340
rect 8878 52288 8930 52340
rect 9002 52288 9054 52340
rect 9126 52288 9178 52340
rect 9250 52288 9302 52340
rect 9374 52288 9426 52340
rect 9498 52288 9550 52340
rect 9622 52288 9674 52340
rect 9746 52288 9798 52340
rect 10256 52288 10308 52340
rect 10380 52288 10432 52340
rect 10504 52288 10556 52340
rect 10628 52288 10680 52340
rect 10752 52288 10804 52340
rect 10876 52288 10928 52340
rect 11000 52288 11052 52340
rect 11124 52288 11176 52340
rect 11248 52288 11300 52340
rect 11372 52288 11424 52340
rect 11496 52288 11548 52340
rect 11620 52288 11672 52340
rect 11744 52288 11796 52340
rect 11868 52288 11920 52340
rect 11992 52288 12044 52340
rect 12116 52288 12168 52340
rect 4863 51983 4915 52017
rect 4987 51983 5039 52017
rect 7277 51983 7329 52017
rect 7401 51983 7453 52017
rect 7525 51983 7577 52017
rect 7649 51983 7701 52017
rect 9939 51983 9991 52017
rect 10063 51983 10115 52017
rect 4863 51965 4915 51983
rect 4987 51965 5039 51983
rect 7277 51965 7329 51983
rect 7401 51965 7453 51983
rect 7525 51965 7577 51983
rect 7649 51965 7701 51983
rect 9939 51965 9991 51983
rect 10063 51965 10115 51983
rect 4863 51875 4915 51893
rect 4987 51875 5039 51893
rect 7277 51875 7329 51893
rect 7401 51875 7453 51893
rect 7525 51875 7577 51893
rect 7649 51875 7701 51893
rect 9939 51875 9991 51893
rect 10063 51875 10115 51893
rect 4863 51841 4915 51875
rect 4987 51841 5039 51875
rect 7277 51841 7329 51875
rect 7401 51841 7453 51875
rect 7525 51841 7577 51875
rect 7649 51841 7701 51875
rect 9939 51841 9991 51875
rect 10063 51841 10115 51875
rect 3559 51626 3611 51627
rect 3683 51626 3735 51627
rect 3807 51626 3859 51627
rect 3931 51626 3983 51627
rect 4055 51626 4107 51627
rect 4179 51626 4231 51627
rect 4303 51626 4355 51627
rect 4427 51626 4479 51627
rect 4551 51626 4603 51627
rect 4675 51626 4727 51627
rect 5180 51626 5232 51627
rect 5304 51626 5356 51627
rect 5428 51626 5480 51627
rect 5552 51626 5604 51627
rect 5676 51626 5728 51627
rect 5800 51626 5852 51627
rect 5924 51626 5976 51627
rect 6048 51626 6100 51627
rect 6172 51626 6224 51627
rect 6296 51626 6348 51627
rect 6420 51626 6472 51627
rect 6544 51626 6596 51627
rect 6668 51626 6720 51627
rect 6792 51626 6844 51627
rect 6916 51626 6968 51627
rect 7040 51626 7092 51627
rect 7886 51626 7938 51627
rect 8010 51626 8062 51627
rect 8134 51626 8186 51627
rect 8258 51626 8310 51627
rect 8382 51626 8434 51627
rect 8506 51626 8558 51627
rect 8630 51626 8682 51627
rect 8754 51626 8806 51627
rect 8878 51626 8930 51627
rect 9002 51626 9054 51627
rect 9126 51626 9178 51627
rect 9250 51626 9302 51627
rect 9374 51626 9426 51627
rect 9498 51626 9550 51627
rect 9622 51626 9674 51627
rect 9746 51626 9798 51627
rect 10251 51626 10303 51627
rect 10375 51626 10427 51627
rect 10499 51626 10551 51627
rect 10623 51626 10675 51627
rect 10747 51626 10799 51627
rect 10871 51626 10923 51627
rect 10995 51626 11047 51627
rect 11119 51626 11171 51627
rect 11243 51626 11295 51627
rect 11367 51626 11419 51627
rect 3559 51580 3611 51626
rect 3683 51580 3735 51626
rect 3807 51580 3859 51626
rect 3931 51580 3983 51626
rect 4055 51580 4107 51626
rect 4179 51580 4231 51626
rect 4303 51580 4355 51626
rect 4427 51580 4479 51626
rect 4551 51580 4603 51626
rect 4675 51580 4727 51626
rect 5180 51580 5232 51626
rect 5304 51580 5356 51626
rect 5428 51580 5480 51626
rect 5552 51580 5604 51626
rect 5676 51580 5728 51626
rect 5800 51580 5852 51626
rect 5924 51580 5976 51626
rect 6048 51580 6100 51626
rect 6172 51580 6224 51626
rect 6296 51580 6348 51626
rect 6420 51580 6472 51626
rect 6544 51580 6596 51626
rect 6668 51580 6720 51626
rect 6792 51580 6844 51626
rect 6916 51580 6968 51626
rect 7040 51580 7092 51626
rect 7886 51580 7938 51626
rect 8010 51580 8062 51626
rect 8134 51580 8186 51626
rect 8258 51580 8310 51626
rect 8382 51580 8434 51626
rect 8506 51580 8558 51626
rect 8630 51580 8682 51626
rect 8754 51580 8806 51626
rect 8878 51580 8930 51626
rect 9002 51580 9054 51626
rect 9126 51580 9178 51626
rect 9250 51580 9302 51626
rect 9374 51580 9426 51626
rect 9498 51580 9550 51626
rect 9622 51580 9674 51626
rect 9746 51580 9798 51626
rect 10251 51580 10303 51626
rect 10375 51580 10427 51626
rect 10499 51580 10551 51626
rect 10623 51580 10675 51626
rect 10747 51580 10799 51626
rect 10871 51580 10923 51626
rect 10995 51580 11047 51626
rect 11119 51580 11171 51626
rect 11243 51580 11295 51626
rect 11367 51580 11419 51626
rect 3559 51575 3611 51580
rect 3683 51575 3735 51580
rect 3807 51575 3859 51580
rect 3931 51575 3983 51580
rect 4055 51575 4107 51580
rect 4179 51575 4231 51580
rect 4303 51575 4355 51580
rect 4427 51575 4479 51580
rect 4551 51575 4603 51580
rect 4675 51575 4727 51580
rect 5180 51575 5232 51580
rect 5304 51575 5356 51580
rect 5428 51575 5480 51580
rect 5552 51575 5604 51580
rect 5676 51575 5728 51580
rect 5800 51575 5852 51580
rect 5924 51575 5976 51580
rect 6048 51575 6100 51580
rect 6172 51575 6224 51580
rect 6296 51575 6348 51580
rect 6420 51575 6472 51580
rect 6544 51575 6596 51580
rect 6668 51575 6720 51580
rect 6792 51575 6844 51580
rect 6916 51575 6968 51580
rect 7040 51575 7092 51580
rect 7886 51575 7938 51580
rect 8010 51575 8062 51580
rect 8134 51575 8186 51580
rect 8258 51575 8310 51580
rect 8382 51575 8434 51580
rect 8506 51575 8558 51580
rect 8630 51575 8682 51580
rect 8754 51575 8806 51580
rect 8878 51575 8930 51580
rect 9002 51575 9054 51580
rect 9126 51575 9178 51580
rect 9250 51575 9302 51580
rect 9374 51575 9426 51580
rect 9498 51575 9550 51580
rect 9622 51575 9674 51580
rect 9746 51575 9798 51580
rect 10251 51575 10303 51580
rect 10375 51575 10427 51580
rect 10499 51575 10551 51580
rect 10623 51575 10675 51580
rect 10747 51575 10799 51580
rect 10871 51575 10923 51580
rect 10995 51575 11047 51580
rect 11119 51575 11171 51580
rect 11243 51575 11295 51580
rect 11367 51575 11419 51580
rect 3559 51498 3611 51503
rect 3683 51498 3735 51503
rect 3807 51498 3859 51503
rect 3931 51498 3983 51503
rect 4055 51498 4107 51503
rect 4179 51498 4231 51503
rect 4303 51498 4355 51503
rect 4427 51498 4479 51503
rect 4551 51498 4603 51503
rect 4675 51498 4727 51503
rect 5180 51498 5232 51503
rect 5304 51498 5356 51503
rect 5428 51498 5480 51503
rect 5552 51498 5604 51503
rect 5676 51498 5728 51503
rect 5800 51498 5852 51503
rect 5924 51498 5976 51503
rect 6048 51498 6100 51503
rect 6172 51498 6224 51503
rect 6296 51498 6348 51503
rect 6420 51498 6472 51503
rect 6544 51498 6596 51503
rect 6668 51498 6720 51503
rect 6792 51498 6844 51503
rect 6916 51498 6968 51503
rect 7040 51498 7092 51503
rect 7886 51498 7938 51503
rect 8010 51498 8062 51503
rect 8134 51498 8186 51503
rect 8258 51498 8310 51503
rect 8382 51498 8434 51503
rect 8506 51498 8558 51503
rect 8630 51498 8682 51503
rect 8754 51498 8806 51503
rect 8878 51498 8930 51503
rect 9002 51498 9054 51503
rect 9126 51498 9178 51503
rect 9250 51498 9302 51503
rect 9374 51498 9426 51503
rect 9498 51498 9550 51503
rect 9622 51498 9674 51503
rect 9746 51498 9798 51503
rect 10251 51498 10303 51503
rect 10375 51498 10427 51503
rect 10499 51498 10551 51503
rect 10623 51498 10675 51503
rect 10747 51498 10799 51503
rect 10871 51498 10923 51503
rect 10995 51498 11047 51503
rect 11119 51498 11171 51503
rect 11243 51498 11295 51503
rect 11367 51498 11419 51503
rect 3559 51452 3611 51498
rect 3683 51452 3735 51498
rect 3807 51452 3859 51498
rect 3931 51452 3983 51498
rect 4055 51452 4107 51498
rect 4179 51452 4231 51498
rect 4303 51452 4355 51498
rect 4427 51452 4479 51498
rect 4551 51452 4603 51498
rect 4675 51452 4727 51498
rect 5180 51452 5232 51498
rect 5304 51452 5356 51498
rect 5428 51452 5480 51498
rect 5552 51452 5604 51498
rect 5676 51452 5728 51498
rect 5800 51452 5852 51498
rect 5924 51452 5976 51498
rect 6048 51452 6100 51498
rect 6172 51452 6224 51498
rect 6296 51452 6348 51498
rect 6420 51452 6472 51498
rect 6544 51452 6596 51498
rect 6668 51452 6720 51498
rect 6792 51452 6844 51498
rect 6916 51452 6968 51498
rect 7040 51452 7092 51498
rect 7886 51452 7938 51498
rect 8010 51452 8062 51498
rect 8134 51452 8186 51498
rect 8258 51452 8310 51498
rect 8382 51452 8434 51498
rect 8506 51452 8558 51498
rect 8630 51452 8682 51498
rect 8754 51452 8806 51498
rect 8878 51452 8930 51498
rect 9002 51452 9054 51498
rect 9126 51452 9178 51498
rect 9250 51452 9302 51498
rect 9374 51452 9426 51498
rect 9498 51452 9550 51498
rect 9622 51452 9674 51498
rect 9746 51452 9798 51498
rect 10251 51452 10303 51498
rect 10375 51452 10427 51498
rect 10499 51452 10551 51498
rect 10623 51452 10675 51498
rect 10747 51452 10799 51498
rect 10871 51452 10923 51498
rect 10995 51452 11047 51498
rect 11119 51452 11171 51498
rect 11243 51452 11295 51498
rect 11367 51452 11419 51498
rect 3559 51451 3611 51452
rect 3683 51451 3735 51452
rect 3807 51451 3859 51452
rect 3931 51451 3983 51452
rect 4055 51451 4107 51452
rect 4179 51451 4231 51452
rect 4303 51451 4355 51452
rect 4427 51451 4479 51452
rect 4551 51451 4603 51452
rect 4675 51451 4727 51452
rect 5180 51451 5232 51452
rect 5304 51451 5356 51452
rect 5428 51451 5480 51452
rect 5552 51451 5604 51452
rect 5676 51451 5728 51452
rect 5800 51451 5852 51452
rect 5924 51451 5976 51452
rect 6048 51451 6100 51452
rect 6172 51451 6224 51452
rect 6296 51451 6348 51452
rect 6420 51451 6472 51452
rect 6544 51451 6596 51452
rect 6668 51451 6720 51452
rect 6792 51451 6844 51452
rect 6916 51451 6968 51452
rect 7040 51451 7092 51452
rect 7886 51451 7938 51452
rect 8010 51451 8062 51452
rect 8134 51451 8186 51452
rect 8258 51451 8310 51452
rect 8382 51451 8434 51452
rect 8506 51451 8558 51452
rect 8630 51451 8682 51452
rect 8754 51451 8806 51452
rect 8878 51451 8930 51452
rect 9002 51451 9054 51452
rect 9126 51451 9178 51452
rect 9250 51451 9302 51452
rect 9374 51451 9426 51452
rect 9498 51451 9550 51452
rect 9622 51451 9674 51452
rect 9746 51451 9798 51452
rect 10251 51451 10303 51452
rect 10375 51451 10427 51452
rect 10499 51451 10551 51452
rect 10623 51451 10675 51452
rect 10747 51451 10799 51452
rect 10871 51451 10923 51452
rect 10995 51451 11047 51452
rect 11119 51451 11171 51452
rect 11243 51451 11295 51452
rect 11367 51451 11419 51452
rect 4863 51203 4915 51222
rect 4987 51203 5039 51222
rect 7277 51203 7329 51222
rect 7401 51203 7453 51222
rect 7525 51203 7577 51222
rect 7649 51203 7701 51222
rect 9939 51203 9991 51222
rect 10063 51203 10115 51222
rect 4863 51170 4915 51203
rect 4987 51170 5039 51203
rect 7277 51170 7329 51203
rect 7401 51170 7453 51203
rect 7525 51170 7577 51203
rect 7649 51170 7701 51203
rect 9939 51170 9991 51203
rect 10063 51170 10115 51203
rect 4863 51095 4915 51098
rect 4987 51095 5039 51098
rect 7277 51095 7329 51098
rect 7401 51095 7453 51098
rect 7525 51095 7577 51098
rect 7649 51095 7701 51098
rect 9939 51095 9991 51098
rect 10063 51095 10115 51098
rect 4863 51049 4915 51095
rect 4987 51049 5039 51095
rect 7277 51049 7329 51095
rect 7401 51049 7453 51095
rect 7525 51049 7577 51095
rect 7649 51049 7701 51095
rect 9939 51049 9991 51095
rect 10063 51049 10115 51095
rect 4863 51046 4915 51049
rect 4987 51046 5039 51049
rect 7277 51046 7329 51049
rect 7401 51046 7453 51049
rect 7525 51046 7577 51049
rect 7649 51046 7701 51049
rect 9939 51046 9991 51049
rect 10063 51046 10115 51049
rect 4863 50941 4915 50974
rect 4987 50941 5039 50974
rect 7277 50941 7329 50974
rect 7401 50941 7453 50974
rect 7525 50941 7577 50974
rect 7649 50941 7701 50974
rect 9939 50941 9991 50974
rect 10063 50941 10115 50974
rect 4863 50922 4915 50941
rect 4987 50922 5039 50941
rect 7277 50922 7329 50941
rect 7401 50922 7453 50941
rect 7525 50922 7577 50941
rect 7649 50922 7701 50941
rect 9939 50922 9991 50941
rect 10063 50922 10115 50941
rect 3559 50692 3611 50693
rect 3683 50692 3735 50693
rect 3807 50692 3859 50693
rect 3931 50692 3983 50693
rect 4055 50692 4107 50693
rect 4179 50692 4231 50693
rect 4303 50692 4355 50693
rect 4427 50692 4479 50693
rect 4551 50692 4603 50693
rect 4675 50692 4727 50693
rect 5180 50692 5232 50693
rect 5304 50692 5356 50693
rect 5428 50692 5480 50693
rect 5552 50692 5604 50693
rect 5676 50692 5728 50693
rect 5800 50692 5852 50693
rect 5924 50692 5976 50693
rect 6048 50692 6100 50693
rect 6172 50692 6224 50693
rect 6296 50692 6348 50693
rect 6420 50692 6472 50693
rect 6544 50692 6596 50693
rect 6668 50692 6720 50693
rect 6792 50692 6844 50693
rect 6916 50692 6968 50693
rect 7040 50692 7092 50693
rect 7886 50692 7938 50693
rect 8010 50692 8062 50693
rect 8134 50692 8186 50693
rect 8258 50692 8310 50693
rect 8382 50692 8434 50693
rect 8506 50692 8558 50693
rect 8630 50692 8682 50693
rect 8754 50692 8806 50693
rect 8878 50692 8930 50693
rect 9002 50692 9054 50693
rect 9126 50692 9178 50693
rect 9250 50692 9302 50693
rect 9374 50692 9426 50693
rect 9498 50692 9550 50693
rect 9622 50692 9674 50693
rect 9746 50692 9798 50693
rect 10251 50692 10303 50693
rect 10375 50692 10427 50693
rect 10499 50692 10551 50693
rect 10623 50692 10675 50693
rect 10747 50692 10799 50693
rect 10871 50692 10923 50693
rect 10995 50692 11047 50693
rect 11119 50692 11171 50693
rect 11243 50692 11295 50693
rect 11367 50692 11419 50693
rect 3559 50646 3611 50692
rect 3683 50646 3735 50692
rect 3807 50646 3859 50692
rect 3931 50646 3983 50692
rect 4055 50646 4107 50692
rect 4179 50646 4231 50692
rect 4303 50646 4355 50692
rect 4427 50646 4479 50692
rect 4551 50646 4603 50692
rect 4675 50646 4727 50692
rect 5180 50646 5232 50692
rect 5304 50646 5356 50692
rect 5428 50646 5480 50692
rect 5552 50646 5604 50692
rect 5676 50646 5728 50692
rect 5800 50646 5852 50692
rect 5924 50646 5976 50692
rect 6048 50646 6100 50692
rect 6172 50646 6224 50692
rect 6296 50646 6348 50692
rect 6420 50646 6472 50692
rect 6544 50646 6596 50692
rect 6668 50646 6720 50692
rect 6792 50646 6844 50692
rect 6916 50646 6968 50692
rect 7040 50646 7092 50692
rect 7886 50646 7938 50692
rect 8010 50646 8062 50692
rect 8134 50646 8186 50692
rect 8258 50646 8310 50692
rect 8382 50646 8434 50692
rect 8506 50646 8558 50692
rect 8630 50646 8682 50692
rect 8754 50646 8806 50692
rect 8878 50646 8930 50692
rect 9002 50646 9054 50692
rect 9126 50646 9178 50692
rect 9250 50646 9302 50692
rect 9374 50646 9426 50692
rect 9498 50646 9550 50692
rect 9622 50646 9674 50692
rect 9746 50646 9798 50692
rect 10251 50646 10303 50692
rect 10375 50646 10427 50692
rect 10499 50646 10551 50692
rect 10623 50646 10675 50692
rect 10747 50646 10799 50692
rect 10871 50646 10923 50692
rect 10995 50646 11047 50692
rect 11119 50646 11171 50692
rect 11243 50646 11295 50692
rect 11367 50646 11419 50692
rect 3559 50641 3611 50646
rect 3683 50641 3735 50646
rect 3807 50641 3859 50646
rect 3931 50641 3983 50646
rect 4055 50641 4107 50646
rect 4179 50641 4231 50646
rect 4303 50641 4355 50646
rect 4427 50641 4479 50646
rect 4551 50641 4603 50646
rect 4675 50641 4727 50646
rect 5180 50641 5232 50646
rect 5304 50641 5356 50646
rect 5428 50641 5480 50646
rect 5552 50641 5604 50646
rect 5676 50641 5728 50646
rect 5800 50641 5852 50646
rect 5924 50641 5976 50646
rect 6048 50641 6100 50646
rect 6172 50641 6224 50646
rect 6296 50641 6348 50646
rect 6420 50641 6472 50646
rect 6544 50641 6596 50646
rect 6668 50641 6720 50646
rect 6792 50641 6844 50646
rect 6916 50641 6968 50646
rect 7040 50641 7092 50646
rect 7886 50641 7938 50646
rect 8010 50641 8062 50646
rect 8134 50641 8186 50646
rect 8258 50641 8310 50646
rect 8382 50641 8434 50646
rect 8506 50641 8558 50646
rect 8630 50641 8682 50646
rect 8754 50641 8806 50646
rect 8878 50641 8930 50646
rect 9002 50641 9054 50646
rect 9126 50641 9178 50646
rect 9250 50641 9302 50646
rect 9374 50641 9426 50646
rect 9498 50641 9550 50646
rect 9622 50641 9674 50646
rect 9746 50641 9798 50646
rect 10251 50641 10303 50646
rect 10375 50641 10427 50646
rect 10499 50641 10551 50646
rect 10623 50641 10675 50646
rect 10747 50641 10799 50646
rect 10871 50641 10923 50646
rect 10995 50641 11047 50646
rect 11119 50641 11171 50646
rect 11243 50641 11295 50646
rect 11367 50641 11419 50646
rect 3559 50564 3611 50569
rect 3683 50564 3735 50569
rect 3807 50564 3859 50569
rect 3931 50564 3983 50569
rect 4055 50564 4107 50569
rect 4179 50564 4231 50569
rect 4303 50564 4355 50569
rect 4427 50564 4479 50569
rect 4551 50564 4603 50569
rect 4675 50564 4727 50569
rect 5180 50564 5232 50569
rect 5304 50564 5356 50569
rect 5428 50564 5480 50569
rect 5552 50564 5604 50569
rect 5676 50564 5728 50569
rect 5800 50564 5852 50569
rect 5924 50564 5976 50569
rect 6048 50564 6100 50569
rect 6172 50564 6224 50569
rect 6296 50564 6348 50569
rect 6420 50564 6472 50569
rect 6544 50564 6596 50569
rect 6668 50564 6720 50569
rect 6792 50564 6844 50569
rect 6916 50564 6968 50569
rect 7040 50564 7092 50569
rect 7886 50564 7938 50569
rect 8010 50564 8062 50569
rect 8134 50564 8186 50569
rect 8258 50564 8310 50569
rect 8382 50564 8434 50569
rect 8506 50564 8558 50569
rect 8630 50564 8682 50569
rect 8754 50564 8806 50569
rect 8878 50564 8930 50569
rect 9002 50564 9054 50569
rect 9126 50564 9178 50569
rect 9250 50564 9302 50569
rect 9374 50564 9426 50569
rect 9498 50564 9550 50569
rect 9622 50564 9674 50569
rect 9746 50564 9798 50569
rect 10251 50564 10303 50569
rect 10375 50564 10427 50569
rect 10499 50564 10551 50569
rect 10623 50564 10675 50569
rect 10747 50564 10799 50569
rect 10871 50564 10923 50569
rect 10995 50564 11047 50569
rect 11119 50564 11171 50569
rect 11243 50564 11295 50569
rect 11367 50564 11419 50569
rect 3559 50518 3611 50564
rect 3683 50518 3735 50564
rect 3807 50518 3859 50564
rect 3931 50518 3983 50564
rect 4055 50518 4107 50564
rect 4179 50518 4231 50564
rect 4303 50518 4355 50564
rect 4427 50518 4479 50564
rect 4551 50518 4603 50564
rect 4675 50518 4727 50564
rect 5180 50518 5232 50564
rect 5304 50518 5356 50564
rect 5428 50518 5480 50564
rect 5552 50518 5604 50564
rect 5676 50518 5728 50564
rect 5800 50518 5852 50564
rect 5924 50518 5976 50564
rect 6048 50518 6100 50564
rect 6172 50518 6224 50564
rect 6296 50518 6348 50564
rect 6420 50518 6472 50564
rect 6544 50518 6596 50564
rect 6668 50518 6720 50564
rect 6792 50518 6844 50564
rect 6916 50518 6968 50564
rect 7040 50518 7092 50564
rect 7886 50518 7938 50564
rect 8010 50518 8062 50564
rect 8134 50518 8186 50564
rect 8258 50518 8310 50564
rect 8382 50518 8434 50564
rect 8506 50518 8558 50564
rect 8630 50518 8682 50564
rect 8754 50518 8806 50564
rect 8878 50518 8930 50564
rect 9002 50518 9054 50564
rect 9126 50518 9178 50564
rect 9250 50518 9302 50564
rect 9374 50518 9426 50564
rect 9498 50518 9550 50564
rect 9622 50518 9674 50564
rect 9746 50518 9798 50564
rect 10251 50518 10303 50564
rect 10375 50518 10427 50564
rect 10499 50518 10551 50564
rect 10623 50518 10675 50564
rect 10747 50518 10799 50564
rect 10871 50518 10923 50564
rect 10995 50518 11047 50564
rect 11119 50518 11171 50564
rect 11243 50518 11295 50564
rect 11367 50518 11419 50564
rect 3559 50517 3611 50518
rect 3683 50517 3735 50518
rect 3807 50517 3859 50518
rect 3931 50517 3983 50518
rect 4055 50517 4107 50518
rect 4179 50517 4231 50518
rect 4303 50517 4355 50518
rect 4427 50517 4479 50518
rect 4551 50517 4603 50518
rect 4675 50517 4727 50518
rect 5180 50517 5232 50518
rect 5304 50517 5356 50518
rect 5428 50517 5480 50518
rect 5552 50517 5604 50518
rect 5676 50517 5728 50518
rect 5800 50517 5852 50518
rect 5924 50517 5976 50518
rect 6048 50517 6100 50518
rect 6172 50517 6224 50518
rect 6296 50517 6348 50518
rect 6420 50517 6472 50518
rect 6544 50517 6596 50518
rect 6668 50517 6720 50518
rect 6792 50517 6844 50518
rect 6916 50517 6968 50518
rect 7040 50517 7092 50518
rect 7886 50517 7938 50518
rect 8010 50517 8062 50518
rect 8134 50517 8186 50518
rect 8258 50517 8310 50518
rect 8382 50517 8434 50518
rect 8506 50517 8558 50518
rect 8630 50517 8682 50518
rect 8754 50517 8806 50518
rect 8878 50517 8930 50518
rect 9002 50517 9054 50518
rect 9126 50517 9178 50518
rect 9250 50517 9302 50518
rect 9374 50517 9426 50518
rect 9498 50517 9550 50518
rect 9622 50517 9674 50518
rect 9746 50517 9798 50518
rect 10251 50517 10303 50518
rect 10375 50517 10427 50518
rect 10499 50517 10551 50518
rect 10623 50517 10675 50518
rect 10747 50517 10799 50518
rect 10871 50517 10923 50518
rect 10995 50517 11047 50518
rect 11119 50517 11171 50518
rect 11243 50517 11295 50518
rect 11367 50517 11419 50518
rect 4863 50269 4915 50288
rect 4987 50269 5039 50288
rect 7277 50269 7329 50288
rect 7401 50269 7453 50288
rect 7525 50269 7577 50288
rect 7649 50269 7701 50288
rect 9939 50269 9991 50288
rect 10063 50269 10115 50288
rect 4863 50236 4915 50269
rect 4987 50236 5039 50269
rect 7277 50236 7329 50269
rect 7401 50236 7453 50269
rect 7525 50236 7577 50269
rect 7649 50236 7701 50269
rect 9939 50236 9991 50269
rect 10063 50236 10115 50269
rect 4863 50161 4915 50164
rect 4987 50161 5039 50164
rect 7277 50161 7329 50164
rect 7401 50161 7453 50164
rect 7525 50161 7577 50164
rect 7649 50161 7701 50164
rect 9939 50161 9991 50164
rect 10063 50161 10115 50164
rect 4863 50115 4915 50161
rect 4987 50115 5039 50161
rect 7277 50115 7329 50161
rect 7401 50115 7453 50161
rect 7525 50115 7577 50161
rect 7649 50115 7701 50161
rect 9939 50115 9991 50161
rect 10063 50115 10115 50161
rect 4863 50112 4915 50115
rect 4987 50112 5039 50115
rect 7277 50112 7329 50115
rect 7401 50112 7453 50115
rect 7525 50112 7577 50115
rect 7649 50112 7701 50115
rect 9939 50112 9991 50115
rect 10063 50112 10115 50115
rect 4863 50007 4915 50040
rect 4987 50007 5039 50040
rect 7277 50007 7329 50040
rect 7401 50007 7453 50040
rect 7525 50007 7577 50040
rect 7649 50007 7701 50040
rect 9939 50007 9991 50040
rect 10063 50007 10115 50040
rect 4863 49988 4915 50007
rect 4987 49988 5039 50007
rect 7277 49988 7329 50007
rect 7401 49988 7453 50007
rect 7525 49988 7577 50007
rect 7649 49988 7701 50007
rect 9939 49988 9991 50007
rect 10063 49988 10115 50007
rect 3559 49758 3611 49759
rect 3683 49758 3735 49759
rect 3807 49758 3859 49759
rect 3931 49758 3983 49759
rect 4055 49758 4107 49759
rect 4179 49758 4231 49759
rect 4303 49758 4355 49759
rect 4427 49758 4479 49759
rect 4551 49758 4603 49759
rect 4675 49758 4727 49759
rect 5180 49758 5232 49759
rect 5304 49758 5356 49759
rect 5428 49758 5480 49759
rect 5552 49758 5604 49759
rect 5676 49758 5728 49759
rect 5800 49758 5852 49759
rect 5924 49758 5976 49759
rect 6048 49758 6100 49759
rect 6172 49758 6224 49759
rect 6296 49758 6348 49759
rect 6420 49758 6472 49759
rect 6544 49758 6596 49759
rect 6668 49758 6720 49759
rect 6792 49758 6844 49759
rect 6916 49758 6968 49759
rect 7040 49758 7092 49759
rect 7886 49758 7938 49759
rect 8010 49758 8062 49759
rect 8134 49758 8186 49759
rect 8258 49758 8310 49759
rect 8382 49758 8434 49759
rect 8506 49758 8558 49759
rect 8630 49758 8682 49759
rect 8754 49758 8806 49759
rect 8878 49758 8930 49759
rect 9002 49758 9054 49759
rect 9126 49758 9178 49759
rect 9250 49758 9302 49759
rect 9374 49758 9426 49759
rect 9498 49758 9550 49759
rect 9622 49758 9674 49759
rect 9746 49758 9798 49759
rect 10251 49758 10303 49759
rect 10375 49758 10427 49759
rect 10499 49758 10551 49759
rect 10623 49758 10675 49759
rect 10747 49758 10799 49759
rect 10871 49758 10923 49759
rect 10995 49758 11047 49759
rect 11119 49758 11171 49759
rect 11243 49758 11295 49759
rect 11367 49758 11419 49759
rect 3559 49712 3611 49758
rect 3683 49712 3735 49758
rect 3807 49712 3859 49758
rect 3931 49712 3983 49758
rect 4055 49712 4107 49758
rect 4179 49712 4231 49758
rect 4303 49712 4355 49758
rect 4427 49712 4479 49758
rect 4551 49712 4603 49758
rect 4675 49712 4727 49758
rect 5180 49712 5232 49758
rect 5304 49712 5356 49758
rect 5428 49712 5480 49758
rect 5552 49712 5604 49758
rect 5676 49712 5728 49758
rect 5800 49712 5852 49758
rect 5924 49712 5976 49758
rect 6048 49712 6100 49758
rect 6172 49712 6224 49758
rect 6296 49712 6348 49758
rect 6420 49712 6472 49758
rect 6544 49712 6596 49758
rect 6668 49712 6720 49758
rect 6792 49712 6844 49758
rect 6916 49712 6968 49758
rect 7040 49712 7092 49758
rect 7886 49712 7938 49758
rect 8010 49712 8062 49758
rect 8134 49712 8186 49758
rect 8258 49712 8310 49758
rect 8382 49712 8434 49758
rect 8506 49712 8558 49758
rect 8630 49712 8682 49758
rect 8754 49712 8806 49758
rect 8878 49712 8930 49758
rect 9002 49712 9054 49758
rect 9126 49712 9178 49758
rect 9250 49712 9302 49758
rect 9374 49712 9426 49758
rect 9498 49712 9550 49758
rect 9622 49712 9674 49758
rect 9746 49712 9798 49758
rect 10251 49712 10303 49758
rect 10375 49712 10427 49758
rect 10499 49712 10551 49758
rect 10623 49712 10675 49758
rect 10747 49712 10799 49758
rect 10871 49712 10923 49758
rect 10995 49712 11047 49758
rect 11119 49712 11171 49758
rect 11243 49712 11295 49758
rect 11367 49712 11419 49758
rect 3559 49707 3611 49712
rect 3683 49707 3735 49712
rect 3807 49707 3859 49712
rect 3931 49707 3983 49712
rect 4055 49707 4107 49712
rect 4179 49707 4231 49712
rect 4303 49707 4355 49712
rect 4427 49707 4479 49712
rect 4551 49707 4603 49712
rect 4675 49707 4727 49712
rect 5180 49707 5232 49712
rect 5304 49707 5356 49712
rect 5428 49707 5480 49712
rect 5552 49707 5604 49712
rect 5676 49707 5728 49712
rect 5800 49707 5852 49712
rect 5924 49707 5976 49712
rect 6048 49707 6100 49712
rect 6172 49707 6224 49712
rect 6296 49707 6348 49712
rect 6420 49707 6472 49712
rect 6544 49707 6596 49712
rect 6668 49707 6720 49712
rect 6792 49707 6844 49712
rect 6916 49707 6968 49712
rect 7040 49707 7092 49712
rect 7886 49707 7938 49712
rect 8010 49707 8062 49712
rect 8134 49707 8186 49712
rect 8258 49707 8310 49712
rect 8382 49707 8434 49712
rect 8506 49707 8558 49712
rect 8630 49707 8682 49712
rect 8754 49707 8806 49712
rect 8878 49707 8930 49712
rect 9002 49707 9054 49712
rect 9126 49707 9178 49712
rect 9250 49707 9302 49712
rect 9374 49707 9426 49712
rect 9498 49707 9550 49712
rect 9622 49707 9674 49712
rect 9746 49707 9798 49712
rect 10251 49707 10303 49712
rect 10375 49707 10427 49712
rect 10499 49707 10551 49712
rect 10623 49707 10675 49712
rect 10747 49707 10799 49712
rect 10871 49707 10923 49712
rect 10995 49707 11047 49712
rect 11119 49707 11171 49712
rect 11243 49707 11295 49712
rect 11367 49707 11419 49712
rect 3559 49630 3611 49635
rect 3683 49630 3735 49635
rect 3807 49630 3859 49635
rect 3931 49630 3983 49635
rect 4055 49630 4107 49635
rect 4179 49630 4231 49635
rect 4303 49630 4355 49635
rect 4427 49630 4479 49635
rect 4551 49630 4603 49635
rect 4675 49630 4727 49635
rect 5180 49630 5232 49635
rect 5304 49630 5356 49635
rect 5428 49630 5480 49635
rect 5552 49630 5604 49635
rect 5676 49630 5728 49635
rect 5800 49630 5852 49635
rect 5924 49630 5976 49635
rect 6048 49630 6100 49635
rect 6172 49630 6224 49635
rect 6296 49630 6348 49635
rect 6420 49630 6472 49635
rect 6544 49630 6596 49635
rect 6668 49630 6720 49635
rect 6792 49630 6844 49635
rect 6916 49630 6968 49635
rect 7040 49630 7092 49635
rect 7886 49630 7938 49635
rect 8010 49630 8062 49635
rect 8134 49630 8186 49635
rect 8258 49630 8310 49635
rect 8382 49630 8434 49635
rect 8506 49630 8558 49635
rect 8630 49630 8682 49635
rect 8754 49630 8806 49635
rect 8878 49630 8930 49635
rect 9002 49630 9054 49635
rect 9126 49630 9178 49635
rect 9250 49630 9302 49635
rect 9374 49630 9426 49635
rect 9498 49630 9550 49635
rect 9622 49630 9674 49635
rect 9746 49630 9798 49635
rect 10251 49630 10303 49635
rect 10375 49630 10427 49635
rect 10499 49630 10551 49635
rect 10623 49630 10675 49635
rect 10747 49630 10799 49635
rect 10871 49630 10923 49635
rect 10995 49630 11047 49635
rect 11119 49630 11171 49635
rect 11243 49630 11295 49635
rect 11367 49630 11419 49635
rect 3559 49584 3611 49630
rect 3683 49584 3735 49630
rect 3807 49584 3859 49630
rect 3931 49584 3983 49630
rect 4055 49584 4107 49630
rect 4179 49584 4231 49630
rect 4303 49584 4355 49630
rect 4427 49584 4479 49630
rect 4551 49584 4603 49630
rect 4675 49584 4727 49630
rect 5180 49584 5232 49630
rect 5304 49584 5356 49630
rect 5428 49584 5480 49630
rect 5552 49584 5604 49630
rect 5676 49584 5728 49630
rect 5800 49584 5852 49630
rect 5924 49584 5976 49630
rect 6048 49584 6100 49630
rect 6172 49584 6224 49630
rect 6296 49584 6348 49630
rect 6420 49584 6472 49630
rect 6544 49584 6596 49630
rect 6668 49584 6720 49630
rect 6792 49584 6844 49630
rect 6916 49584 6968 49630
rect 7040 49584 7092 49630
rect 7886 49584 7938 49630
rect 8010 49584 8062 49630
rect 8134 49584 8186 49630
rect 8258 49584 8310 49630
rect 8382 49584 8434 49630
rect 8506 49584 8558 49630
rect 8630 49584 8682 49630
rect 8754 49584 8806 49630
rect 8878 49584 8930 49630
rect 9002 49584 9054 49630
rect 9126 49584 9178 49630
rect 9250 49584 9302 49630
rect 9374 49584 9426 49630
rect 9498 49584 9550 49630
rect 9622 49584 9674 49630
rect 9746 49584 9798 49630
rect 10251 49584 10303 49630
rect 10375 49584 10427 49630
rect 10499 49584 10551 49630
rect 10623 49584 10675 49630
rect 10747 49584 10799 49630
rect 10871 49584 10923 49630
rect 10995 49584 11047 49630
rect 11119 49584 11171 49630
rect 11243 49584 11295 49630
rect 11367 49584 11419 49630
rect 3559 49583 3611 49584
rect 3683 49583 3735 49584
rect 3807 49583 3859 49584
rect 3931 49583 3983 49584
rect 4055 49583 4107 49584
rect 4179 49583 4231 49584
rect 4303 49583 4355 49584
rect 4427 49583 4479 49584
rect 4551 49583 4603 49584
rect 4675 49583 4727 49584
rect 5180 49583 5232 49584
rect 5304 49583 5356 49584
rect 5428 49583 5480 49584
rect 5552 49583 5604 49584
rect 5676 49583 5728 49584
rect 5800 49583 5852 49584
rect 5924 49583 5976 49584
rect 6048 49583 6100 49584
rect 6172 49583 6224 49584
rect 6296 49583 6348 49584
rect 6420 49583 6472 49584
rect 6544 49583 6596 49584
rect 6668 49583 6720 49584
rect 6792 49583 6844 49584
rect 6916 49583 6968 49584
rect 7040 49583 7092 49584
rect 7886 49583 7938 49584
rect 8010 49583 8062 49584
rect 8134 49583 8186 49584
rect 8258 49583 8310 49584
rect 8382 49583 8434 49584
rect 8506 49583 8558 49584
rect 8630 49583 8682 49584
rect 8754 49583 8806 49584
rect 8878 49583 8930 49584
rect 9002 49583 9054 49584
rect 9126 49583 9178 49584
rect 9250 49583 9302 49584
rect 9374 49583 9426 49584
rect 9498 49583 9550 49584
rect 9622 49583 9674 49584
rect 9746 49583 9798 49584
rect 10251 49583 10303 49584
rect 10375 49583 10427 49584
rect 10499 49583 10551 49584
rect 10623 49583 10675 49584
rect 10747 49583 10799 49584
rect 10871 49583 10923 49584
rect 10995 49583 11047 49584
rect 11119 49583 11171 49584
rect 11243 49583 11295 49584
rect 11367 49583 11419 49584
rect 4863 49335 4915 49354
rect 4987 49335 5039 49354
rect 7277 49335 7329 49354
rect 7401 49335 7453 49354
rect 7525 49335 7577 49354
rect 7649 49335 7701 49354
rect 9939 49335 9991 49354
rect 10063 49335 10115 49354
rect 4863 49302 4915 49335
rect 4987 49302 5039 49335
rect 7277 49302 7329 49335
rect 7401 49302 7453 49335
rect 7525 49302 7577 49335
rect 7649 49302 7701 49335
rect 9939 49302 9991 49335
rect 10063 49302 10115 49335
rect 4863 49227 4915 49230
rect 4987 49227 5039 49230
rect 7277 49227 7329 49230
rect 7401 49227 7453 49230
rect 7525 49227 7577 49230
rect 7649 49227 7701 49230
rect 9939 49227 9991 49230
rect 10063 49227 10115 49230
rect 4863 49181 4915 49227
rect 4987 49181 5039 49227
rect 7277 49181 7329 49227
rect 7401 49181 7453 49227
rect 7525 49181 7577 49227
rect 7649 49181 7701 49227
rect 9939 49181 9991 49227
rect 10063 49181 10115 49227
rect 4863 49178 4915 49181
rect 4987 49178 5039 49181
rect 7277 49178 7329 49181
rect 7401 49178 7453 49181
rect 7525 49178 7577 49181
rect 7649 49178 7701 49181
rect 9939 49178 9991 49181
rect 10063 49178 10115 49181
rect 4863 49073 4915 49106
rect 4987 49073 5039 49106
rect 7277 49073 7329 49106
rect 7401 49073 7453 49106
rect 7525 49073 7577 49106
rect 7649 49073 7701 49106
rect 9939 49073 9991 49106
rect 10063 49073 10115 49106
rect 4863 49054 4915 49073
rect 4987 49054 5039 49073
rect 7277 49054 7329 49073
rect 7401 49054 7453 49073
rect 7525 49054 7577 49073
rect 7649 49054 7701 49073
rect 9939 49054 9991 49073
rect 10063 49054 10115 49073
rect 3559 48824 3611 48825
rect 3683 48824 3735 48825
rect 3807 48824 3859 48825
rect 3931 48824 3983 48825
rect 4055 48824 4107 48825
rect 4179 48824 4231 48825
rect 4303 48824 4355 48825
rect 4427 48824 4479 48825
rect 4551 48824 4603 48825
rect 4675 48824 4727 48825
rect 5180 48824 5232 48825
rect 5304 48824 5356 48825
rect 5428 48824 5480 48825
rect 5552 48824 5604 48825
rect 5676 48824 5728 48825
rect 5800 48824 5852 48825
rect 5924 48824 5976 48825
rect 6048 48824 6100 48825
rect 6172 48824 6224 48825
rect 6296 48824 6348 48825
rect 6420 48824 6472 48825
rect 6544 48824 6596 48825
rect 6668 48824 6720 48825
rect 6792 48824 6844 48825
rect 6916 48824 6968 48825
rect 7040 48824 7092 48825
rect 7886 48824 7938 48825
rect 8010 48824 8062 48825
rect 8134 48824 8186 48825
rect 8258 48824 8310 48825
rect 8382 48824 8434 48825
rect 8506 48824 8558 48825
rect 8630 48824 8682 48825
rect 8754 48824 8806 48825
rect 8878 48824 8930 48825
rect 9002 48824 9054 48825
rect 9126 48824 9178 48825
rect 9250 48824 9302 48825
rect 9374 48824 9426 48825
rect 9498 48824 9550 48825
rect 9622 48824 9674 48825
rect 9746 48824 9798 48825
rect 10251 48824 10303 48825
rect 10375 48824 10427 48825
rect 10499 48824 10551 48825
rect 10623 48824 10675 48825
rect 10747 48824 10799 48825
rect 10871 48824 10923 48825
rect 10995 48824 11047 48825
rect 11119 48824 11171 48825
rect 11243 48824 11295 48825
rect 11367 48824 11419 48825
rect 3559 48778 3611 48824
rect 3683 48778 3735 48824
rect 3807 48778 3859 48824
rect 3931 48778 3983 48824
rect 4055 48778 4107 48824
rect 4179 48778 4231 48824
rect 4303 48778 4355 48824
rect 4427 48778 4479 48824
rect 4551 48778 4603 48824
rect 4675 48778 4727 48824
rect 5180 48778 5232 48824
rect 5304 48778 5356 48824
rect 5428 48778 5480 48824
rect 5552 48778 5604 48824
rect 5676 48778 5728 48824
rect 5800 48778 5852 48824
rect 5924 48778 5976 48824
rect 6048 48778 6100 48824
rect 6172 48778 6224 48824
rect 6296 48778 6348 48824
rect 6420 48778 6472 48824
rect 6544 48778 6596 48824
rect 6668 48778 6720 48824
rect 6792 48778 6844 48824
rect 6916 48778 6968 48824
rect 7040 48778 7092 48824
rect 7886 48778 7938 48824
rect 8010 48778 8062 48824
rect 8134 48778 8186 48824
rect 8258 48778 8310 48824
rect 8382 48778 8434 48824
rect 8506 48778 8558 48824
rect 8630 48778 8682 48824
rect 8754 48778 8806 48824
rect 8878 48778 8930 48824
rect 9002 48778 9054 48824
rect 9126 48778 9178 48824
rect 9250 48778 9302 48824
rect 9374 48778 9426 48824
rect 9498 48778 9550 48824
rect 9622 48778 9674 48824
rect 9746 48778 9798 48824
rect 10251 48778 10303 48824
rect 10375 48778 10427 48824
rect 10499 48778 10551 48824
rect 10623 48778 10675 48824
rect 10747 48778 10799 48824
rect 10871 48778 10923 48824
rect 10995 48778 11047 48824
rect 11119 48778 11171 48824
rect 11243 48778 11295 48824
rect 11367 48778 11419 48824
rect 3559 48773 3611 48778
rect 3683 48773 3735 48778
rect 3807 48773 3859 48778
rect 3931 48773 3983 48778
rect 4055 48773 4107 48778
rect 4179 48773 4231 48778
rect 4303 48773 4355 48778
rect 4427 48773 4479 48778
rect 4551 48773 4603 48778
rect 4675 48773 4727 48778
rect 5180 48773 5232 48778
rect 5304 48773 5356 48778
rect 5428 48773 5480 48778
rect 5552 48773 5604 48778
rect 5676 48773 5728 48778
rect 5800 48773 5852 48778
rect 5924 48773 5976 48778
rect 6048 48773 6100 48778
rect 6172 48773 6224 48778
rect 6296 48773 6348 48778
rect 6420 48773 6472 48778
rect 6544 48773 6596 48778
rect 6668 48773 6720 48778
rect 6792 48773 6844 48778
rect 6916 48773 6968 48778
rect 7040 48773 7092 48778
rect 7886 48773 7938 48778
rect 8010 48773 8062 48778
rect 8134 48773 8186 48778
rect 8258 48773 8310 48778
rect 8382 48773 8434 48778
rect 8506 48773 8558 48778
rect 8630 48773 8682 48778
rect 8754 48773 8806 48778
rect 8878 48773 8930 48778
rect 9002 48773 9054 48778
rect 9126 48773 9178 48778
rect 9250 48773 9302 48778
rect 9374 48773 9426 48778
rect 9498 48773 9550 48778
rect 9622 48773 9674 48778
rect 9746 48773 9798 48778
rect 10251 48773 10303 48778
rect 10375 48773 10427 48778
rect 10499 48773 10551 48778
rect 10623 48773 10675 48778
rect 10747 48773 10799 48778
rect 10871 48773 10923 48778
rect 10995 48773 11047 48778
rect 11119 48773 11171 48778
rect 11243 48773 11295 48778
rect 11367 48773 11419 48778
rect 3559 48696 3611 48701
rect 3683 48696 3735 48701
rect 3807 48696 3859 48701
rect 3931 48696 3983 48701
rect 4055 48696 4107 48701
rect 4179 48696 4231 48701
rect 4303 48696 4355 48701
rect 4427 48696 4479 48701
rect 4551 48696 4603 48701
rect 4675 48696 4727 48701
rect 5180 48696 5232 48701
rect 5304 48696 5356 48701
rect 5428 48696 5480 48701
rect 5552 48696 5604 48701
rect 5676 48696 5728 48701
rect 5800 48696 5852 48701
rect 5924 48696 5976 48701
rect 6048 48696 6100 48701
rect 6172 48696 6224 48701
rect 6296 48696 6348 48701
rect 6420 48696 6472 48701
rect 6544 48696 6596 48701
rect 6668 48696 6720 48701
rect 6792 48696 6844 48701
rect 6916 48696 6968 48701
rect 7040 48696 7092 48701
rect 7886 48696 7938 48701
rect 8010 48696 8062 48701
rect 8134 48696 8186 48701
rect 8258 48696 8310 48701
rect 8382 48696 8434 48701
rect 8506 48696 8558 48701
rect 8630 48696 8682 48701
rect 8754 48696 8806 48701
rect 8878 48696 8930 48701
rect 9002 48696 9054 48701
rect 9126 48696 9178 48701
rect 9250 48696 9302 48701
rect 9374 48696 9426 48701
rect 9498 48696 9550 48701
rect 9622 48696 9674 48701
rect 9746 48696 9798 48701
rect 10251 48696 10303 48701
rect 10375 48696 10427 48701
rect 10499 48696 10551 48701
rect 10623 48696 10675 48701
rect 10747 48696 10799 48701
rect 10871 48696 10923 48701
rect 10995 48696 11047 48701
rect 11119 48696 11171 48701
rect 11243 48696 11295 48701
rect 11367 48696 11419 48701
rect 3559 48650 3611 48696
rect 3683 48650 3735 48696
rect 3807 48650 3859 48696
rect 3931 48650 3983 48696
rect 4055 48650 4107 48696
rect 4179 48650 4231 48696
rect 4303 48650 4355 48696
rect 4427 48650 4479 48696
rect 4551 48650 4603 48696
rect 4675 48650 4727 48696
rect 5180 48650 5232 48696
rect 5304 48650 5356 48696
rect 5428 48650 5480 48696
rect 5552 48650 5604 48696
rect 5676 48650 5728 48696
rect 5800 48650 5852 48696
rect 5924 48650 5976 48696
rect 6048 48650 6100 48696
rect 6172 48650 6224 48696
rect 6296 48650 6348 48696
rect 6420 48650 6472 48696
rect 6544 48650 6596 48696
rect 6668 48650 6720 48696
rect 6792 48650 6844 48696
rect 6916 48650 6968 48696
rect 7040 48650 7092 48696
rect 7886 48650 7938 48696
rect 8010 48650 8062 48696
rect 8134 48650 8186 48696
rect 8258 48650 8310 48696
rect 8382 48650 8434 48696
rect 8506 48650 8558 48696
rect 8630 48650 8682 48696
rect 8754 48650 8806 48696
rect 8878 48650 8930 48696
rect 9002 48650 9054 48696
rect 9126 48650 9178 48696
rect 9250 48650 9302 48696
rect 9374 48650 9426 48696
rect 9498 48650 9550 48696
rect 9622 48650 9674 48696
rect 9746 48650 9798 48696
rect 10251 48650 10303 48696
rect 10375 48650 10427 48696
rect 10499 48650 10551 48696
rect 10623 48650 10675 48696
rect 10747 48650 10799 48696
rect 10871 48650 10923 48696
rect 10995 48650 11047 48696
rect 11119 48650 11171 48696
rect 11243 48650 11295 48696
rect 11367 48650 11419 48696
rect 3559 48649 3611 48650
rect 3683 48649 3735 48650
rect 3807 48649 3859 48650
rect 3931 48649 3983 48650
rect 4055 48649 4107 48650
rect 4179 48649 4231 48650
rect 4303 48649 4355 48650
rect 4427 48649 4479 48650
rect 4551 48649 4603 48650
rect 4675 48649 4727 48650
rect 5180 48649 5232 48650
rect 5304 48649 5356 48650
rect 5428 48649 5480 48650
rect 5552 48649 5604 48650
rect 5676 48649 5728 48650
rect 5800 48649 5852 48650
rect 5924 48649 5976 48650
rect 6048 48649 6100 48650
rect 6172 48649 6224 48650
rect 6296 48649 6348 48650
rect 6420 48649 6472 48650
rect 6544 48649 6596 48650
rect 6668 48649 6720 48650
rect 6792 48649 6844 48650
rect 6916 48649 6968 48650
rect 7040 48649 7092 48650
rect 7886 48649 7938 48650
rect 8010 48649 8062 48650
rect 8134 48649 8186 48650
rect 8258 48649 8310 48650
rect 8382 48649 8434 48650
rect 8506 48649 8558 48650
rect 8630 48649 8682 48650
rect 8754 48649 8806 48650
rect 8878 48649 8930 48650
rect 9002 48649 9054 48650
rect 9126 48649 9178 48650
rect 9250 48649 9302 48650
rect 9374 48649 9426 48650
rect 9498 48649 9550 48650
rect 9622 48649 9674 48650
rect 9746 48649 9798 48650
rect 10251 48649 10303 48650
rect 10375 48649 10427 48650
rect 10499 48649 10551 48650
rect 10623 48649 10675 48650
rect 10747 48649 10799 48650
rect 10871 48649 10923 48650
rect 10995 48649 11047 48650
rect 11119 48649 11171 48650
rect 11243 48649 11295 48650
rect 11367 48649 11419 48650
rect 4863 48401 4915 48435
rect 4987 48401 5039 48435
rect 7277 48401 7329 48435
rect 7401 48401 7453 48435
rect 7525 48401 7577 48435
rect 7649 48401 7701 48435
rect 9939 48401 9991 48435
rect 10063 48401 10115 48435
rect 4863 48383 4915 48401
rect 4987 48383 5039 48401
rect 7277 48383 7329 48401
rect 7401 48383 7453 48401
rect 7525 48383 7577 48401
rect 7649 48383 7701 48401
rect 9939 48383 9991 48401
rect 10063 48383 10115 48401
rect 4863 48293 4915 48311
rect 4987 48293 5039 48311
rect 7277 48293 7329 48311
rect 7401 48293 7453 48311
rect 7525 48293 7577 48311
rect 7649 48293 7701 48311
rect 9939 48293 9991 48311
rect 10063 48293 10115 48311
rect 4863 48259 4915 48293
rect 4987 48259 5039 48293
rect 7277 48259 7329 48293
rect 7401 48259 7453 48293
rect 7525 48259 7577 48293
rect 7649 48259 7701 48293
rect 9939 48259 9991 48293
rect 10063 48259 10115 48293
rect 2810 47936 2862 47988
rect 2934 47936 2986 47988
rect 3058 47936 3110 47988
rect 3182 47936 3234 47988
rect 3306 47936 3358 47988
rect 3430 47936 3482 47988
rect 3554 47936 3606 47988
rect 3678 47936 3730 47988
rect 3802 47936 3854 47988
rect 3926 47936 3978 47988
rect 4050 47936 4102 47988
rect 4174 47936 4226 47988
rect 4298 47936 4350 47988
rect 4422 47936 4474 47988
rect 4546 47936 4598 47988
rect 4670 47936 4722 47988
rect 5180 47936 5232 47988
rect 5304 47936 5356 47988
rect 5428 47936 5480 47988
rect 5552 47936 5604 47988
rect 5676 47936 5728 47988
rect 5800 47936 5852 47988
rect 5924 47936 5976 47988
rect 6048 47936 6100 47988
rect 6172 47936 6224 47988
rect 6296 47936 6348 47988
rect 6420 47936 6472 47988
rect 6544 47936 6596 47988
rect 6668 47936 6720 47988
rect 6792 47936 6844 47988
rect 6916 47936 6968 47988
rect 7040 47936 7092 47988
rect 7886 47936 7938 47988
rect 8010 47936 8062 47988
rect 8134 47936 8186 47988
rect 8258 47936 8310 47988
rect 8382 47936 8434 47988
rect 8506 47936 8558 47988
rect 8630 47936 8682 47988
rect 8754 47936 8806 47988
rect 8878 47936 8930 47988
rect 9002 47936 9054 47988
rect 9126 47936 9178 47988
rect 9250 47936 9302 47988
rect 9374 47936 9426 47988
rect 9498 47936 9550 47988
rect 9622 47936 9674 47988
rect 9746 47936 9798 47988
rect 10256 47936 10308 47988
rect 10380 47936 10432 47988
rect 10504 47936 10556 47988
rect 10628 47936 10680 47988
rect 10752 47936 10804 47988
rect 10876 47936 10928 47988
rect 11000 47936 11052 47988
rect 11124 47936 11176 47988
rect 11248 47936 11300 47988
rect 11372 47936 11424 47988
rect 11496 47936 11548 47988
rect 11620 47936 11672 47988
rect 11744 47936 11796 47988
rect 11868 47936 11920 47988
rect 11992 47936 12044 47988
rect 12116 47936 12168 47988
rect 2810 47812 2862 47864
rect 2934 47812 2986 47864
rect 3058 47812 3110 47864
rect 3182 47812 3234 47864
rect 3306 47812 3358 47864
rect 3430 47812 3482 47864
rect 3554 47812 3606 47864
rect 3678 47812 3730 47864
rect 3802 47812 3854 47864
rect 3926 47812 3978 47864
rect 4050 47812 4102 47864
rect 4174 47812 4226 47864
rect 4298 47812 4350 47864
rect 4422 47812 4474 47864
rect 4546 47812 4598 47864
rect 4670 47812 4722 47864
rect 5180 47812 5232 47864
rect 5304 47812 5356 47864
rect 5428 47812 5480 47864
rect 5552 47812 5604 47864
rect 5676 47812 5728 47864
rect 5800 47812 5852 47864
rect 5924 47812 5976 47864
rect 6048 47812 6100 47864
rect 6172 47812 6224 47864
rect 6296 47812 6348 47864
rect 6420 47812 6472 47864
rect 6544 47812 6596 47864
rect 6668 47812 6720 47864
rect 6792 47812 6844 47864
rect 6916 47812 6968 47864
rect 7040 47812 7092 47864
rect 7886 47812 7938 47864
rect 8010 47812 8062 47864
rect 8134 47812 8186 47864
rect 8258 47812 8310 47864
rect 8382 47812 8434 47864
rect 8506 47812 8558 47864
rect 8630 47812 8682 47864
rect 8754 47812 8806 47864
rect 8878 47812 8930 47864
rect 9002 47812 9054 47864
rect 9126 47812 9178 47864
rect 9250 47812 9302 47864
rect 9374 47812 9426 47864
rect 9498 47812 9550 47864
rect 9622 47812 9674 47864
rect 9746 47812 9798 47864
rect 10256 47812 10308 47864
rect 10380 47812 10432 47864
rect 10504 47812 10556 47864
rect 10628 47812 10680 47864
rect 10752 47812 10804 47864
rect 10876 47812 10928 47864
rect 11000 47812 11052 47864
rect 11124 47812 11176 47864
rect 11248 47812 11300 47864
rect 11372 47812 11424 47864
rect 11496 47812 11548 47864
rect 11620 47812 11672 47864
rect 11744 47812 11796 47864
rect 11868 47812 11920 47864
rect 11992 47812 12044 47864
rect 12116 47812 12168 47864
rect 2810 47688 2862 47740
rect 2934 47688 2986 47740
rect 3058 47688 3110 47740
rect 3182 47688 3234 47740
rect 3306 47688 3358 47740
rect 3430 47688 3482 47740
rect 3554 47688 3606 47740
rect 3678 47688 3730 47740
rect 3802 47688 3854 47740
rect 3926 47688 3978 47740
rect 4050 47688 4102 47740
rect 4174 47688 4226 47740
rect 4298 47688 4350 47740
rect 4422 47688 4474 47740
rect 4546 47688 4598 47740
rect 4670 47688 4722 47740
rect 5180 47688 5232 47740
rect 5304 47688 5356 47740
rect 5428 47688 5480 47740
rect 5552 47688 5604 47740
rect 5676 47688 5728 47740
rect 5800 47688 5852 47740
rect 5924 47688 5976 47740
rect 6048 47688 6100 47740
rect 6172 47688 6224 47740
rect 6296 47688 6348 47740
rect 6420 47688 6472 47740
rect 6544 47688 6596 47740
rect 6668 47688 6720 47740
rect 6792 47688 6844 47740
rect 6916 47688 6968 47740
rect 7040 47688 7092 47740
rect 7886 47688 7938 47740
rect 8010 47688 8062 47740
rect 8134 47688 8186 47740
rect 8258 47688 8310 47740
rect 8382 47688 8434 47740
rect 8506 47688 8558 47740
rect 8630 47688 8682 47740
rect 8754 47688 8806 47740
rect 8878 47688 8930 47740
rect 9002 47688 9054 47740
rect 9126 47688 9178 47740
rect 9250 47688 9302 47740
rect 9374 47688 9426 47740
rect 9498 47688 9550 47740
rect 9622 47688 9674 47740
rect 9746 47688 9798 47740
rect 10256 47688 10308 47740
rect 10380 47688 10432 47740
rect 10504 47688 10556 47740
rect 10628 47688 10680 47740
rect 10752 47688 10804 47740
rect 10876 47688 10928 47740
rect 11000 47688 11052 47740
rect 11124 47688 11176 47740
rect 11248 47688 11300 47740
rect 11372 47688 11424 47740
rect 11496 47688 11548 47740
rect 11620 47688 11672 47740
rect 11744 47688 11796 47740
rect 11868 47688 11920 47740
rect 11992 47688 12044 47740
rect 12116 47688 12168 47740
rect 14904 52522 14956 52574
rect 14904 52414 14956 52466
rect 14904 52306 14956 52358
rect 14904 52198 14956 52250
rect 14904 52090 14956 52142
rect 14904 51982 14956 52034
rect 14904 51874 14956 51926
rect 14904 51766 14956 51818
rect 14904 51658 14956 51710
rect 14904 51550 14956 51602
rect 14904 51442 14956 51494
rect 14904 51334 14956 51386
rect 14904 51226 14956 51278
rect 22 38122 74 38174
rect 22 38014 74 38066
rect 22 37906 74 37958
rect 22 37798 74 37850
rect 22 37690 74 37742
rect 22 37582 74 37634
rect 22 37474 74 37526
rect 22 37366 74 37418
rect 22 37258 74 37310
rect 22 37150 74 37202
rect 22 37042 74 37094
rect 22 36934 74 36986
rect 22 36826 74 36878
rect 14904 38122 14956 38174
rect 14904 38014 14956 38066
rect 14904 37906 14956 37958
rect 14904 37798 14956 37850
rect 14904 37690 14956 37742
rect 14904 37582 14956 37634
rect 14904 37474 14956 37526
rect 14904 37366 14956 37418
rect 14904 37258 14956 37310
rect 14904 37150 14956 37202
rect 14904 37042 14956 37094
rect 14904 36934 14956 36986
rect 14904 36826 14956 36878
<< metal2 >>
rect 261 56669 2161 57600
rect 261 56617 917 56669
rect 969 56617 1041 56669
rect 1093 56617 1165 56669
rect 1217 56617 1289 56669
rect 1341 56617 1413 56669
rect 1465 56617 1537 56669
rect 1589 56617 1661 56669
rect 1713 56617 1785 56669
rect 1837 56617 2161 56669
rect 261 56545 2161 56617
rect 261 56493 917 56545
rect 969 56493 1041 56545
rect 1093 56493 1165 56545
rect 1217 56493 1289 56545
rect 1341 56493 1413 56545
rect 1465 56493 1537 56545
rect 1589 56493 1661 56545
rect 1713 56493 1785 56545
rect 1837 56493 2161 56545
rect 261 56421 2161 56493
rect 261 56369 917 56421
rect 969 56369 1041 56421
rect 1093 56369 1165 56421
rect 1217 56369 1289 56421
rect 1341 56369 1413 56421
rect 1465 56369 1537 56421
rect 1589 56369 1661 56421
rect 1713 56369 1785 56421
rect 1837 56369 2161 56421
rect 261 56297 2161 56369
rect 261 56245 917 56297
rect 969 56245 1041 56297
rect 1093 56245 1165 56297
rect 1217 56245 1289 56297
rect 1341 56245 1413 56297
rect 1465 56245 1537 56297
rect 1589 56245 1661 56297
rect 1713 56245 1785 56297
rect 1837 56245 2161 56297
rect 261 56173 2161 56245
rect 261 56121 917 56173
rect 969 56121 1041 56173
rect 1093 56121 1165 56173
rect 1217 56121 1289 56173
rect 1341 56121 1413 56173
rect 1465 56121 1537 56173
rect 1589 56121 1661 56173
rect 1713 56121 1785 56173
rect 1837 56121 2161 56173
rect 261 56049 2161 56121
rect 261 55997 917 56049
rect 969 55997 1041 56049
rect 1093 55997 1165 56049
rect 1217 55997 1289 56049
rect 1341 55997 1413 56049
rect 1465 55997 1537 56049
rect 1589 55997 1661 56049
rect 1713 55997 1785 56049
rect 1837 55997 2161 56049
rect 261 55925 2161 55997
rect 261 55873 917 55925
rect 969 55873 1041 55925
rect 1093 55873 1165 55925
rect 1217 55873 1289 55925
rect 1341 55873 1413 55925
rect 1465 55873 1537 55925
rect 1589 55873 1661 55925
rect 1713 55873 1785 55925
rect 1837 55873 2161 55925
rect 261 55801 2161 55873
rect 261 55749 917 55801
rect 969 55749 1041 55801
rect 1093 55749 1165 55801
rect 1217 55749 1289 55801
rect 1341 55749 1413 55801
rect 1465 55749 1537 55801
rect 1589 55749 1661 55801
rect 1713 55749 1785 55801
rect 1837 55749 2161 55801
rect 261 55677 2161 55749
rect 261 55625 917 55677
rect 969 55625 1041 55677
rect 1093 55625 1165 55677
rect 1217 55625 1289 55677
rect 1341 55625 1413 55677
rect 1465 55625 1537 55677
rect 1589 55625 1661 55677
rect 1713 55625 1785 55677
rect 1837 55625 2161 55677
rect 261 55553 2161 55625
rect 261 55501 917 55553
rect 969 55501 1041 55553
rect 1093 55501 1165 55553
rect 1217 55501 1289 55553
rect 1341 55501 1413 55553
rect 1465 55501 1537 55553
rect 1589 55501 1661 55553
rect 1713 55501 1785 55553
rect 1837 55501 2161 55553
rect 261 55429 2161 55501
rect 261 55377 917 55429
rect 969 55377 1041 55429
rect 1093 55377 1165 55429
rect 1217 55377 1289 55429
rect 1341 55377 1413 55429
rect 1465 55377 1537 55429
rect 1589 55377 1661 55429
rect 1713 55377 1785 55429
rect 1837 55377 2161 55429
rect 261 55305 2161 55377
rect 261 55253 917 55305
rect 969 55253 1041 55305
rect 1093 55253 1165 55305
rect 1217 55253 1289 55305
rect 1341 55253 1413 55305
rect 1465 55253 1537 55305
rect 1589 55253 1661 55305
rect 1713 55253 1785 55305
rect 1837 55253 2161 55305
rect 261 55181 2161 55253
rect 261 55129 917 55181
rect 969 55129 1041 55181
rect 1093 55129 1165 55181
rect 1217 55129 1289 55181
rect 1341 55129 1413 55181
rect 1465 55129 1537 55181
rect 1589 55129 1661 55181
rect 1713 55129 1785 55181
rect 1837 55129 2161 55181
rect 261 55057 2161 55129
rect 261 55005 917 55057
rect 969 55005 1041 55057
rect 1093 55005 1165 55057
rect 1217 55005 1289 55057
rect 1341 55005 1413 55057
rect 1465 55005 1537 55057
rect 1589 55005 1661 55057
rect 1713 55005 1785 55057
rect 1837 55005 2161 55057
rect 261 54933 2161 55005
rect 261 54881 917 54933
rect 969 54881 1041 54933
rect 1093 54881 1165 54933
rect 1217 54881 1289 54933
rect 1341 54881 1413 54933
rect 1465 54881 1537 54933
rect 1589 54881 1661 54933
rect 1713 54881 1785 54933
rect 1837 54881 2161 54933
rect 261 54809 2161 54881
rect 261 54757 917 54809
rect 969 54757 1041 54809
rect 1093 54757 1165 54809
rect 1217 54757 1289 54809
rect 1341 54757 1413 54809
rect 1465 54757 1537 54809
rect 1589 54757 1661 54809
rect 1713 54757 1785 54809
rect 1837 54757 2161 54809
rect 261 54685 2161 54757
rect 261 54633 917 54685
rect 969 54633 1041 54685
rect 1093 54633 1165 54685
rect 1217 54633 1289 54685
rect 1341 54633 1413 54685
rect 1465 54633 1537 54685
rect 1589 54633 1661 54685
rect 1713 54633 1785 54685
rect 1837 54633 2161 54685
rect 261 54561 2161 54633
rect 261 54509 917 54561
rect 969 54509 1041 54561
rect 1093 54509 1165 54561
rect 1217 54509 1289 54561
rect 1341 54509 1413 54561
rect 1465 54509 1537 54561
rect 1589 54509 1661 54561
rect 1713 54509 1785 54561
rect 1837 54509 2161 54561
rect 261 54437 2161 54509
rect 261 54385 917 54437
rect 969 54385 1041 54437
rect 1093 54385 1165 54437
rect 1217 54385 1289 54437
rect 1341 54385 1413 54437
rect 1465 54385 1537 54437
rect 1589 54385 1661 54437
rect 1713 54385 1785 54437
rect 1837 54385 2161 54437
rect 261 54313 2161 54385
rect 261 54261 917 54313
rect 969 54261 1041 54313
rect 1093 54261 1165 54313
rect 1217 54261 1289 54313
rect 1341 54261 1413 54313
rect 1465 54261 1537 54313
rect 1589 54261 1661 54313
rect 1713 54261 1785 54313
rect 1837 54261 2161 54313
rect 261 54189 2161 54261
rect 261 54137 917 54189
rect 969 54137 1041 54189
rect 1093 54137 1165 54189
rect 1217 54137 1289 54189
rect 1341 54137 1413 54189
rect 1465 54137 1537 54189
rect 1589 54137 1661 54189
rect 1713 54137 1785 54189
rect 1837 54137 2161 54189
rect 261 54065 2161 54137
rect 261 54013 917 54065
rect 969 54013 1041 54065
rect 1093 54013 1165 54065
rect 1217 54013 1289 54065
rect 1341 54013 1413 54065
rect 1465 54013 1537 54065
rect 1589 54013 1661 54065
rect 1713 54013 1785 54065
rect 1837 54013 2161 54065
rect 261 53941 2161 54013
rect 261 53889 917 53941
rect 969 53889 1041 53941
rect 1093 53889 1165 53941
rect 1217 53889 1289 53941
rect 1341 53889 1413 53941
rect 1465 53889 1537 53941
rect 1589 53889 1661 53941
rect 1713 53889 1785 53941
rect 1837 53889 2161 53941
rect 261 53817 2161 53889
rect 261 53765 917 53817
rect 969 53765 1041 53817
rect 1093 53765 1165 53817
rect 1217 53765 1289 53817
rect 1341 53765 1413 53817
rect 1465 53765 1537 53817
rect 1589 53765 1661 53817
rect 1713 53765 1785 53817
rect 1837 53765 2161 53817
rect 261 53693 2161 53765
rect 261 53641 917 53693
rect 969 53641 1041 53693
rect 1093 53641 1165 53693
rect 1217 53641 1289 53693
rect 1341 53641 1413 53693
rect 1465 53641 1537 53693
rect 1589 53641 1661 53693
rect 1713 53641 1785 53693
rect 1837 53641 2161 53693
rect -11 52576 86 52600
rect -11 51224 20 52576
rect 76 51224 86 52576
rect -11 51200 86 51224
rect 261 50948 2161 53641
rect 2481 57108 2681 57278
rect 2481 57056 2501 57108
rect 2553 57056 2609 57108
rect 2661 57056 2681 57108
rect 2481 53484 2681 57056
rect 2481 53432 2501 53484
rect 2553 53432 2609 53484
rect 2661 53432 2681 53484
rect 2481 53376 2681 53432
rect 2481 53324 2501 53376
rect 2553 53324 2609 53376
rect 2661 53324 2681 53376
rect 2481 53268 2681 53324
rect 2481 53216 2501 53268
rect 2553 53216 2609 53268
rect 2661 53216 2681 53268
rect 261 50892 315 50948
rect 371 50892 439 50948
rect 495 50892 563 50948
rect 619 50892 687 50948
rect 743 50892 811 50948
rect 867 50892 935 50948
rect 991 50892 1059 50948
rect 1115 50892 1183 50948
rect 1239 50892 1307 50948
rect 1363 50892 1431 50948
rect 1487 50892 1555 50948
rect 1611 50892 1679 50948
rect 1735 50892 1803 50948
rect 1859 50892 1927 50948
rect 1983 50892 2051 50948
rect 2107 50892 2161 50948
rect 261 50824 2161 50892
rect 261 50768 315 50824
rect 371 50768 439 50824
rect 495 50768 563 50824
rect 619 50768 687 50824
rect 743 50768 811 50824
rect 867 50768 935 50824
rect 991 50768 1059 50824
rect 1115 50768 1183 50824
rect 1239 50768 1307 50824
rect 1363 50768 1431 50824
rect 1487 50768 1555 50824
rect 1611 50768 1679 50824
rect 1735 50768 1803 50824
rect 1859 50768 1927 50824
rect 1983 50768 2051 50824
rect 2107 50768 2161 50824
rect 261 50700 2161 50768
rect 261 50644 315 50700
rect 371 50644 439 50700
rect 495 50644 563 50700
rect 619 50644 687 50700
rect 743 50644 811 50700
rect 867 50644 935 50700
rect 991 50644 1059 50700
rect 1115 50644 1183 50700
rect 1239 50644 1307 50700
rect 1363 50644 1431 50700
rect 1487 50644 1555 50700
rect 1611 50644 1679 50700
rect 1735 50644 1803 50700
rect 1859 50644 1927 50700
rect 1983 50644 2051 50700
rect 2107 50644 2161 50700
rect 261 50576 2161 50644
rect 261 50520 315 50576
rect 371 50520 439 50576
rect 495 50520 563 50576
rect 619 50520 687 50576
rect 743 50520 811 50576
rect 867 50520 935 50576
rect 991 50520 1059 50576
rect 1115 50520 1183 50576
rect 1239 50520 1307 50576
rect 1363 50520 1431 50576
rect 1487 50520 1555 50576
rect 1611 50520 1679 50576
rect 1735 50520 1803 50576
rect 1859 50520 1927 50576
rect 1983 50520 2051 50576
rect 2107 50520 2161 50576
rect 261 50452 2161 50520
rect 261 50396 315 50452
rect 371 50396 439 50452
rect 495 50396 563 50452
rect 619 50396 687 50452
rect 743 50396 811 50452
rect 867 50396 935 50452
rect 991 50396 1059 50452
rect 1115 50396 1183 50452
rect 1239 50396 1307 50452
rect 1363 50396 1431 50452
rect 1487 50396 1555 50452
rect 1611 50396 1679 50452
rect 1735 50396 1803 50452
rect 1859 50396 1927 50452
rect 1983 50396 2051 50452
rect 2107 50396 2161 50452
rect 261 50328 2161 50396
rect 261 50272 315 50328
rect 371 50272 439 50328
rect 495 50272 563 50328
rect 619 50272 687 50328
rect 743 50272 811 50328
rect 867 50272 935 50328
rect 991 50272 1059 50328
rect 1115 50272 1183 50328
rect 1239 50272 1307 50328
rect 1363 50272 1431 50328
rect 1487 50272 1555 50328
rect 1611 50272 1679 50328
rect 1735 50272 1803 50328
rect 1859 50272 1927 50328
rect 1983 50272 2051 50328
rect 2107 50272 2161 50328
rect 261 50204 2161 50272
rect 261 50148 315 50204
rect 371 50148 439 50204
rect 495 50148 563 50204
rect 619 50148 687 50204
rect 743 50148 811 50204
rect 867 50148 935 50204
rect 991 50148 1059 50204
rect 1115 50148 1183 50204
rect 1239 50148 1307 50204
rect 1363 50148 1431 50204
rect 1487 50148 1555 50204
rect 1611 50148 1679 50204
rect 1735 50148 1803 50204
rect 1859 50148 1927 50204
rect 1983 50148 2051 50204
rect 2107 50148 2161 50204
rect 261 50080 2161 50148
rect 261 50024 315 50080
rect 371 50024 439 50080
rect 495 50024 563 50080
rect 619 50024 687 50080
rect 743 50024 811 50080
rect 867 50024 935 50080
rect 991 50024 1059 50080
rect 1115 50024 1183 50080
rect 1239 50024 1307 50080
rect 1363 50024 1431 50080
rect 1487 50024 1555 50080
rect 1611 50024 1679 50080
rect 1735 50024 1803 50080
rect 1859 50024 1927 50080
rect 1983 50024 2051 50080
rect 2107 50024 2161 50080
rect 261 49956 2161 50024
rect 261 49900 315 49956
rect 371 49900 439 49956
rect 495 49900 563 49956
rect 619 49900 687 49956
rect 743 49900 811 49956
rect 867 49900 935 49956
rect 991 49900 1059 49956
rect 1115 49900 1183 49956
rect 1239 49900 1307 49956
rect 1363 49900 1431 49956
rect 1487 49900 1555 49956
rect 1611 49900 1679 49956
rect 1735 49900 1803 49956
rect 1859 49900 1927 49956
rect 1983 49900 2051 49956
rect 2107 49900 2161 49956
rect 261 49832 2161 49900
rect 261 49776 315 49832
rect 371 49776 439 49832
rect 495 49776 563 49832
rect 619 49776 687 49832
rect 743 49776 811 49832
rect 867 49776 935 49832
rect 991 49776 1059 49832
rect 1115 49776 1183 49832
rect 1239 49776 1307 49832
rect 1363 49776 1431 49832
rect 1487 49776 1555 49832
rect 1611 49776 1679 49832
rect 1735 49776 1803 49832
rect 1859 49776 1927 49832
rect 1983 49776 2051 49832
rect 2107 49776 2161 49832
rect 261 49708 2161 49776
rect 261 49652 315 49708
rect 371 49652 439 49708
rect 495 49652 563 49708
rect 619 49652 687 49708
rect 743 49652 811 49708
rect 867 49652 935 49708
rect 991 49652 1059 49708
rect 1115 49652 1183 49708
rect 1239 49652 1307 49708
rect 1363 49652 1431 49708
rect 1487 49652 1555 49708
rect 1611 49652 1679 49708
rect 1735 49652 1803 49708
rect 1859 49652 1927 49708
rect 1983 49652 2051 49708
rect 2107 49652 2161 49708
rect 261 46430 2161 49652
rect 2279 52521 2355 52600
rect 2279 52465 2289 52521
rect 2345 52465 2355 52521
rect 2279 52389 2355 52465
rect 2279 52333 2289 52389
rect 2345 52333 2355 52389
rect 2279 52257 2355 52333
rect 2279 52201 2289 52257
rect 2345 52201 2355 52257
rect 2279 52125 2355 52201
rect 2279 52069 2289 52125
rect 2345 52069 2355 52125
rect 2279 51993 2355 52069
rect 2279 51937 2289 51993
rect 2345 51937 2355 51993
rect 2279 51861 2355 51937
rect 2279 51805 2289 51861
rect 2345 51805 2355 51861
rect 2279 51729 2355 51805
rect 2279 51673 2289 51729
rect 2345 51673 2355 51729
rect 2279 51597 2355 51673
rect 2279 51541 2289 51597
rect 2345 51541 2355 51597
rect 2279 51465 2355 51541
rect 2279 51409 2289 51465
rect 2345 51409 2355 51465
rect 2279 51333 2355 51409
rect 2279 51277 2289 51333
rect 2345 51277 2355 51333
rect 305 43242 2117 44558
rect 305 41642 2117 42958
rect 309 41358 2161 41360
rect 305 40050 2161 41358
rect 305 40042 2117 40050
rect 305 39748 2117 39758
rect 305 39692 315 39748
rect 371 39692 439 39748
rect 495 39692 563 39748
rect 619 39692 687 39748
rect 743 39692 811 39748
rect 867 39692 935 39748
rect 991 39692 1059 39748
rect 1115 39692 1183 39748
rect 1239 39692 1307 39748
rect 1363 39692 1431 39748
rect 1487 39692 1555 39748
rect 1611 39692 1679 39748
rect 1735 39692 1803 39748
rect 1859 39692 1927 39748
rect 1983 39692 2051 39748
rect 2107 39692 2117 39748
rect 305 39624 2117 39692
rect 305 39568 315 39624
rect 371 39568 439 39624
rect 495 39568 563 39624
rect 619 39568 687 39624
rect 743 39568 811 39624
rect 867 39568 935 39624
rect 991 39568 1059 39624
rect 1115 39568 1183 39624
rect 1239 39568 1307 39624
rect 1363 39568 1431 39624
rect 1487 39568 1555 39624
rect 1611 39568 1679 39624
rect 1735 39568 1803 39624
rect 1859 39568 1927 39624
rect 1983 39568 2051 39624
rect 2107 39568 2117 39624
rect 305 39500 2117 39568
rect 305 39444 315 39500
rect 371 39444 439 39500
rect 495 39444 563 39500
rect 619 39444 687 39500
rect 743 39444 811 39500
rect 867 39444 935 39500
rect 991 39444 1059 39500
rect 1115 39444 1183 39500
rect 1239 39444 1307 39500
rect 1363 39444 1431 39500
rect 1487 39444 1555 39500
rect 1611 39444 1679 39500
rect 1735 39444 1803 39500
rect 1859 39444 1927 39500
rect 1983 39444 2051 39500
rect 2107 39444 2117 39500
rect 305 39376 2117 39444
rect 305 39320 315 39376
rect 371 39320 439 39376
rect 495 39320 563 39376
rect 619 39320 687 39376
rect 743 39320 811 39376
rect 867 39320 935 39376
rect 991 39320 1059 39376
rect 1115 39320 1183 39376
rect 1239 39320 1307 39376
rect 1363 39320 1431 39376
rect 1487 39320 1555 39376
rect 1611 39320 1679 39376
rect 1735 39320 1803 39376
rect 1859 39320 1927 39376
rect 1983 39320 2051 39376
rect 2107 39320 2117 39376
rect 305 39252 2117 39320
rect 305 39196 315 39252
rect 371 39196 439 39252
rect 495 39196 563 39252
rect 619 39196 687 39252
rect 743 39196 811 39252
rect 867 39196 935 39252
rect 991 39196 1059 39252
rect 1115 39196 1183 39252
rect 1239 39196 1307 39252
rect 1363 39196 1431 39252
rect 1487 39196 1555 39252
rect 1611 39196 1679 39252
rect 1735 39196 1803 39252
rect 1859 39196 1927 39252
rect 1983 39196 2051 39252
rect 2107 39196 2117 39252
rect 305 39128 2117 39196
rect 305 39072 315 39128
rect 371 39072 439 39128
rect 495 39072 563 39128
rect 619 39072 687 39128
rect 743 39072 811 39128
rect 867 39072 935 39128
rect 991 39072 1059 39128
rect 1115 39072 1183 39128
rect 1239 39072 1307 39128
rect 1363 39072 1431 39128
rect 1487 39072 1555 39128
rect 1611 39072 1679 39128
rect 1735 39072 1803 39128
rect 1859 39072 1927 39128
rect 1983 39072 2051 39128
rect 2107 39072 2117 39128
rect 305 39004 2117 39072
rect 305 38948 315 39004
rect 371 38948 439 39004
rect 495 38948 563 39004
rect 619 38948 687 39004
rect 743 38948 811 39004
rect 867 38948 935 39004
rect 991 38948 1059 39004
rect 1115 38948 1183 39004
rect 1239 38948 1307 39004
rect 1363 38948 1431 39004
rect 1487 38948 1555 39004
rect 1611 38948 1679 39004
rect 1735 38948 1803 39004
rect 1859 38948 1927 39004
rect 1983 38948 2051 39004
rect 2107 38948 2117 39004
rect 305 38880 2117 38948
rect 305 38824 315 38880
rect 371 38824 439 38880
rect 495 38824 563 38880
rect 619 38824 687 38880
rect 743 38824 811 38880
rect 867 38824 935 38880
rect 991 38824 1059 38880
rect 1115 38824 1183 38880
rect 1239 38824 1307 38880
rect 1363 38824 1431 38880
rect 1487 38824 1555 38880
rect 1611 38824 1679 38880
rect 1735 38824 1803 38880
rect 1859 38824 1927 38880
rect 1983 38824 2051 38880
rect 2107 38824 2117 38880
rect 305 38756 2117 38824
rect 305 38700 315 38756
rect 371 38700 439 38756
rect 495 38700 563 38756
rect 619 38700 687 38756
rect 743 38700 811 38756
rect 867 38700 935 38756
rect 991 38700 1059 38756
rect 1115 38700 1183 38756
rect 1239 38700 1307 38756
rect 1363 38700 1431 38756
rect 1487 38700 1555 38756
rect 1611 38700 1679 38756
rect 1735 38700 1803 38756
rect 1859 38700 1927 38756
rect 1983 38700 2051 38756
rect 2107 38700 2117 38756
rect 305 38632 2117 38700
rect 305 38576 315 38632
rect 371 38576 439 38632
rect 495 38576 563 38632
rect 619 38576 687 38632
rect 743 38576 811 38632
rect 867 38576 935 38632
rect 991 38576 1059 38632
rect 1115 38576 1183 38632
rect 1239 38576 1307 38632
rect 1363 38576 1431 38632
rect 1487 38576 1555 38632
rect 1611 38576 1679 38632
rect 1735 38576 1803 38632
rect 1859 38576 1927 38632
rect 1983 38576 2051 38632
rect 2107 38576 2117 38632
rect 305 38508 2117 38576
rect 305 38452 315 38508
rect 371 38452 439 38508
rect 495 38452 563 38508
rect 619 38452 687 38508
rect 743 38452 811 38508
rect 867 38452 935 38508
rect 991 38452 1059 38508
rect 1115 38452 1183 38508
rect 1239 38452 1307 38508
rect 1363 38452 1431 38508
rect 1487 38452 1555 38508
rect 1611 38452 1679 38508
rect 1735 38452 1803 38508
rect 1859 38452 1927 38508
rect 1983 38452 2051 38508
rect 2107 38452 2117 38508
rect 305 38442 2117 38452
rect -11 38176 86 38200
rect -11 36824 20 38176
rect 76 36824 86 38176
rect -11 36800 86 36824
rect 2279 38135 2355 51277
rect 2481 52548 2681 53216
rect 2481 52492 2491 52548
rect 2547 52492 2615 52548
rect 2671 52492 2681 52548
rect 2481 52424 2681 52492
rect 2481 52368 2491 52424
rect 2547 52368 2615 52424
rect 2671 52368 2681 52424
rect 2481 52300 2681 52368
rect 2481 52244 2491 52300
rect 2547 52244 2615 52300
rect 2671 52244 2681 52300
rect 2481 52176 2681 52244
rect 2481 52120 2491 52176
rect 2547 52120 2615 52176
rect 2671 52120 2681 52176
rect 2481 52052 2681 52120
rect 2481 51996 2491 52052
rect 2547 51996 2615 52052
rect 2671 51996 2681 52052
rect 2481 51928 2681 51996
rect 2481 51872 2491 51928
rect 2547 51872 2615 51928
rect 2671 51872 2681 51928
rect 2481 51804 2681 51872
rect 2481 51748 2491 51804
rect 2547 51748 2615 51804
rect 2671 51748 2681 51804
rect 2481 51680 2681 51748
rect 2481 51624 2491 51680
rect 2547 51624 2615 51680
rect 2671 51624 2681 51680
rect 2481 51556 2681 51624
rect 2481 51500 2491 51556
rect 2547 51500 2615 51556
rect 2671 51500 2681 51556
rect 2481 51432 2681 51500
rect 2481 51376 2491 51432
rect 2547 51376 2615 51432
rect 2671 51376 2681 51432
rect 2481 51308 2681 51376
rect 2481 51252 2491 51308
rect 2547 51252 2615 51308
rect 2671 51252 2681 51308
rect 2481 46430 2681 51252
rect 2741 56669 4791 57600
rect 2741 56617 2833 56669
rect 2885 56617 2957 56669
rect 3009 56617 3081 56669
rect 3133 56617 3205 56669
rect 3257 56617 3329 56669
rect 3381 56617 3453 56669
rect 3505 56617 3577 56669
rect 3629 56617 3701 56669
rect 3753 56617 4340 56669
rect 4392 56617 4464 56669
rect 4516 56617 4588 56669
rect 4640 56617 4712 56669
rect 4764 56617 4791 56669
rect 2741 56545 4791 56617
rect 2741 56493 2833 56545
rect 2885 56493 2957 56545
rect 3009 56493 3081 56545
rect 3133 56493 3205 56545
rect 3257 56493 3329 56545
rect 3381 56493 3453 56545
rect 3505 56493 3577 56545
rect 3629 56493 3701 56545
rect 3753 56493 4340 56545
rect 4392 56493 4464 56545
rect 4516 56493 4588 56545
rect 4640 56493 4712 56545
rect 4764 56493 4791 56545
rect 2741 56421 4791 56493
rect 2741 56369 2833 56421
rect 2885 56369 2957 56421
rect 3009 56369 3081 56421
rect 3133 56369 3205 56421
rect 3257 56369 3329 56421
rect 3381 56369 3453 56421
rect 3505 56369 3577 56421
rect 3629 56369 3701 56421
rect 3753 56369 4340 56421
rect 4392 56369 4464 56421
rect 4516 56369 4588 56421
rect 4640 56369 4712 56421
rect 4764 56369 4791 56421
rect 2741 56297 4791 56369
rect 2741 56245 2833 56297
rect 2885 56245 2957 56297
rect 3009 56245 3081 56297
rect 3133 56245 3205 56297
rect 3257 56245 3329 56297
rect 3381 56245 3453 56297
rect 3505 56245 3577 56297
rect 3629 56245 3701 56297
rect 3753 56245 4340 56297
rect 4392 56245 4464 56297
rect 4516 56245 4588 56297
rect 4640 56245 4712 56297
rect 4764 56245 4791 56297
rect 2741 56173 4791 56245
rect 2741 56121 2833 56173
rect 2885 56121 2957 56173
rect 3009 56121 3081 56173
rect 3133 56121 3205 56173
rect 3257 56121 3329 56173
rect 3381 56121 3453 56173
rect 3505 56121 3577 56173
rect 3629 56121 3701 56173
rect 3753 56121 4340 56173
rect 4392 56121 4464 56173
rect 4516 56121 4588 56173
rect 4640 56121 4712 56173
rect 4764 56121 4791 56173
rect 2741 56049 4791 56121
rect 2741 55997 2833 56049
rect 2885 55997 2957 56049
rect 3009 55997 3081 56049
rect 3133 55997 3205 56049
rect 3257 55997 3329 56049
rect 3381 55997 3453 56049
rect 3505 55997 3577 56049
rect 3629 55997 3701 56049
rect 3753 55997 4340 56049
rect 4392 55997 4464 56049
rect 4516 55997 4588 56049
rect 4640 55997 4712 56049
rect 4764 55997 4791 56049
rect 2741 55925 4791 55997
rect 2741 55873 2833 55925
rect 2885 55873 2957 55925
rect 3009 55873 3081 55925
rect 3133 55873 3205 55925
rect 3257 55873 3329 55925
rect 3381 55873 3453 55925
rect 3505 55873 3577 55925
rect 3629 55873 3701 55925
rect 3753 55873 4340 55925
rect 4392 55873 4464 55925
rect 4516 55873 4588 55925
rect 4640 55873 4712 55925
rect 4764 55873 4791 55925
rect 2741 55801 4791 55873
rect 2741 55749 2833 55801
rect 2885 55749 2957 55801
rect 3009 55749 3081 55801
rect 3133 55749 3205 55801
rect 3257 55749 3329 55801
rect 3381 55749 3453 55801
rect 3505 55749 3577 55801
rect 3629 55749 3701 55801
rect 3753 55749 4340 55801
rect 4392 55749 4464 55801
rect 4516 55749 4588 55801
rect 4640 55749 4712 55801
rect 4764 55749 4791 55801
rect 2741 55677 4791 55749
rect 2741 55625 2833 55677
rect 2885 55625 2957 55677
rect 3009 55625 3081 55677
rect 3133 55625 3205 55677
rect 3257 55625 3329 55677
rect 3381 55625 3453 55677
rect 3505 55625 3577 55677
rect 3629 55625 3701 55677
rect 3753 55625 4340 55677
rect 4392 55625 4464 55677
rect 4516 55625 4588 55677
rect 4640 55625 4712 55677
rect 4764 55625 4791 55677
rect 2741 55553 4791 55625
rect 2741 55501 2833 55553
rect 2885 55501 2957 55553
rect 3009 55501 3081 55553
rect 3133 55501 3205 55553
rect 3257 55501 3329 55553
rect 3381 55501 3453 55553
rect 3505 55501 3577 55553
rect 3629 55501 3701 55553
rect 3753 55501 4340 55553
rect 4392 55501 4464 55553
rect 4516 55501 4588 55553
rect 4640 55501 4712 55553
rect 4764 55501 4791 55553
rect 2741 55429 4791 55501
rect 2741 55377 2833 55429
rect 2885 55377 2957 55429
rect 3009 55377 3081 55429
rect 3133 55377 3205 55429
rect 3257 55377 3329 55429
rect 3381 55377 3453 55429
rect 3505 55377 3577 55429
rect 3629 55377 3701 55429
rect 3753 55377 4340 55429
rect 4392 55377 4464 55429
rect 4516 55377 4588 55429
rect 4640 55377 4712 55429
rect 4764 55377 4791 55429
rect 2741 55305 4791 55377
rect 2741 55253 2833 55305
rect 2885 55253 2957 55305
rect 3009 55253 3081 55305
rect 3133 55253 3205 55305
rect 3257 55253 3329 55305
rect 3381 55253 3453 55305
rect 3505 55253 3577 55305
rect 3629 55253 3701 55305
rect 3753 55253 4340 55305
rect 4392 55253 4464 55305
rect 4516 55253 4588 55305
rect 4640 55253 4712 55305
rect 4764 55253 4791 55305
rect 2741 55181 4791 55253
rect 2741 55129 2833 55181
rect 2885 55129 2957 55181
rect 3009 55129 3081 55181
rect 3133 55129 3205 55181
rect 3257 55129 3329 55181
rect 3381 55129 3453 55181
rect 3505 55129 3577 55181
rect 3629 55129 3701 55181
rect 3753 55129 4340 55181
rect 4392 55129 4464 55181
rect 4516 55129 4588 55181
rect 4640 55129 4712 55181
rect 4764 55129 4791 55181
rect 2741 55057 4791 55129
rect 2741 55005 2833 55057
rect 2885 55005 2957 55057
rect 3009 55005 3081 55057
rect 3133 55005 3205 55057
rect 3257 55005 3329 55057
rect 3381 55005 3453 55057
rect 3505 55005 3577 55057
rect 3629 55005 3701 55057
rect 3753 55005 4340 55057
rect 4392 55005 4464 55057
rect 4516 55005 4588 55057
rect 4640 55005 4712 55057
rect 4764 55005 4791 55057
rect 2741 54933 4791 55005
rect 2741 54881 2833 54933
rect 2885 54881 2957 54933
rect 3009 54881 3081 54933
rect 3133 54881 3205 54933
rect 3257 54881 3329 54933
rect 3381 54881 3453 54933
rect 3505 54881 3577 54933
rect 3629 54881 3701 54933
rect 3753 54881 4340 54933
rect 4392 54881 4464 54933
rect 4516 54881 4588 54933
rect 4640 54881 4712 54933
rect 4764 54881 4791 54933
rect 2741 54809 4791 54881
rect 2741 54757 2833 54809
rect 2885 54757 2957 54809
rect 3009 54757 3081 54809
rect 3133 54757 3205 54809
rect 3257 54757 3329 54809
rect 3381 54757 3453 54809
rect 3505 54757 3577 54809
rect 3629 54757 3701 54809
rect 3753 54757 4340 54809
rect 4392 54757 4464 54809
rect 4516 54757 4588 54809
rect 4640 54757 4712 54809
rect 4764 54757 4791 54809
rect 2741 54685 4791 54757
rect 2741 54633 2833 54685
rect 2885 54633 2957 54685
rect 3009 54633 3081 54685
rect 3133 54633 3205 54685
rect 3257 54633 3329 54685
rect 3381 54633 3453 54685
rect 3505 54633 3577 54685
rect 3629 54633 3701 54685
rect 3753 54633 4340 54685
rect 4392 54633 4464 54685
rect 4516 54633 4588 54685
rect 4640 54633 4712 54685
rect 4764 54633 4791 54685
rect 2741 54561 4791 54633
rect 2741 54509 2833 54561
rect 2885 54509 2957 54561
rect 3009 54509 3081 54561
rect 3133 54509 3205 54561
rect 3257 54509 3329 54561
rect 3381 54509 3453 54561
rect 3505 54509 3577 54561
rect 3629 54509 3701 54561
rect 3753 54509 4340 54561
rect 4392 54509 4464 54561
rect 4516 54509 4588 54561
rect 4640 54509 4712 54561
rect 4764 54509 4791 54561
rect 2741 54437 4791 54509
rect 2741 54385 2833 54437
rect 2885 54385 2957 54437
rect 3009 54385 3081 54437
rect 3133 54385 3205 54437
rect 3257 54385 3329 54437
rect 3381 54385 3453 54437
rect 3505 54385 3577 54437
rect 3629 54385 3701 54437
rect 3753 54385 4340 54437
rect 4392 54385 4464 54437
rect 4516 54385 4588 54437
rect 4640 54385 4712 54437
rect 4764 54385 4791 54437
rect 2741 54313 4791 54385
rect 2741 54261 2833 54313
rect 2885 54261 2957 54313
rect 3009 54261 3081 54313
rect 3133 54261 3205 54313
rect 3257 54261 3329 54313
rect 3381 54261 3453 54313
rect 3505 54261 3577 54313
rect 3629 54261 3701 54313
rect 3753 54261 4340 54313
rect 4392 54261 4464 54313
rect 4516 54261 4588 54313
rect 4640 54261 4712 54313
rect 4764 54261 4791 54313
rect 2741 54189 4791 54261
rect 2741 54137 2833 54189
rect 2885 54137 2957 54189
rect 3009 54137 3081 54189
rect 3133 54137 3205 54189
rect 3257 54137 3329 54189
rect 3381 54137 3453 54189
rect 3505 54137 3577 54189
rect 3629 54137 3701 54189
rect 3753 54137 4340 54189
rect 4392 54137 4464 54189
rect 4516 54137 4588 54189
rect 4640 54137 4712 54189
rect 4764 54137 4791 54189
rect 2741 54065 4791 54137
rect 2741 54013 2833 54065
rect 2885 54013 2957 54065
rect 3009 54013 3081 54065
rect 3133 54013 3205 54065
rect 3257 54013 3329 54065
rect 3381 54013 3453 54065
rect 3505 54013 3577 54065
rect 3629 54013 3701 54065
rect 3753 54013 4340 54065
rect 4392 54013 4464 54065
rect 4516 54013 4588 54065
rect 4640 54013 4712 54065
rect 4764 54013 4791 54065
rect 2741 53941 4791 54013
rect 2741 53889 2833 53941
rect 2885 53889 2957 53941
rect 3009 53889 3081 53941
rect 3133 53889 3205 53941
rect 3257 53889 3329 53941
rect 3381 53889 3453 53941
rect 3505 53889 3577 53941
rect 3629 53889 3701 53941
rect 3753 53889 4340 53941
rect 4392 53889 4464 53941
rect 4516 53889 4588 53941
rect 4640 53889 4712 53941
rect 4764 53889 4791 53941
rect 2741 53817 4791 53889
rect 2741 53765 2833 53817
rect 2885 53765 2957 53817
rect 3009 53765 3081 53817
rect 3133 53765 3205 53817
rect 3257 53765 3329 53817
rect 3381 53765 3453 53817
rect 3505 53765 3577 53817
rect 3629 53765 3701 53817
rect 3753 53765 4340 53817
rect 4392 53765 4464 53817
rect 4516 53765 4588 53817
rect 4640 53765 4712 53817
rect 4764 53765 4791 53817
rect 2741 53693 4791 53765
rect 2741 53641 2833 53693
rect 2885 53641 2957 53693
rect 3009 53641 3081 53693
rect 3133 53641 3205 53693
rect 3257 53641 3329 53693
rect 3381 53641 3453 53693
rect 3505 53641 3577 53693
rect 3629 53641 3701 53693
rect 3753 53641 4340 53693
rect 4392 53641 4464 53693
rect 4516 53641 4588 53693
rect 4640 53641 4712 53693
rect 4764 53641 4791 53693
rect 2741 52588 4791 53641
rect 2741 52536 2810 52588
rect 2862 52536 2934 52588
rect 2986 52536 3058 52588
rect 3110 52536 3182 52588
rect 3234 52536 3306 52588
rect 3358 52536 3430 52588
rect 3482 52536 3554 52588
rect 3606 52536 3678 52588
rect 3730 52536 3802 52588
rect 3854 52536 3926 52588
rect 3978 52536 4050 52588
rect 4102 52536 4174 52588
rect 4226 52536 4298 52588
rect 4350 52536 4422 52588
rect 4474 52536 4546 52588
rect 4598 52536 4670 52588
rect 4722 52536 4791 52588
rect 2741 52464 4791 52536
rect 2741 52412 2810 52464
rect 2862 52412 2934 52464
rect 2986 52412 3058 52464
rect 3110 52412 3182 52464
rect 3234 52412 3306 52464
rect 3358 52412 3430 52464
rect 3482 52412 3554 52464
rect 3606 52412 3678 52464
rect 3730 52412 3802 52464
rect 3854 52412 3926 52464
rect 3978 52412 4050 52464
rect 4102 52412 4174 52464
rect 4226 52412 4298 52464
rect 4350 52412 4422 52464
rect 4474 52412 4546 52464
rect 4598 52412 4670 52464
rect 4722 52412 4791 52464
rect 2741 52340 4791 52412
rect 2741 52288 2810 52340
rect 2862 52288 2934 52340
rect 2986 52288 3058 52340
rect 3110 52288 3182 52340
rect 3234 52288 3306 52340
rect 3358 52288 3430 52340
rect 3482 52288 3554 52340
rect 3606 52288 3678 52340
rect 3730 52288 3802 52340
rect 3854 52288 3926 52340
rect 3978 52288 4050 52340
rect 4102 52288 4174 52340
rect 4226 52288 4298 52340
rect 4350 52288 4422 52340
rect 4474 52288 4546 52340
rect 4598 52288 4670 52340
rect 4722 52288 4791 52340
rect 2741 51627 4791 52288
rect 2741 51575 3559 51627
rect 3611 51575 3683 51627
rect 3735 51575 3807 51627
rect 3859 51575 3931 51627
rect 3983 51575 4055 51627
rect 4107 51575 4179 51627
rect 4231 51575 4303 51627
rect 4355 51575 4427 51627
rect 4479 51575 4551 51627
rect 4603 51575 4675 51627
rect 4727 51575 4791 51627
rect 2741 51503 4791 51575
rect 2741 51451 3559 51503
rect 3611 51451 3683 51503
rect 3735 51451 3807 51503
rect 3859 51451 3931 51503
rect 3983 51451 4055 51503
rect 4107 51451 4179 51503
rect 4231 51451 4303 51503
rect 4355 51451 4427 51503
rect 4479 51451 4551 51503
rect 4603 51451 4675 51503
rect 4727 51451 4791 51503
rect 2741 50948 4791 51451
rect 2741 50892 2808 50948
rect 2864 50892 2932 50948
rect 2988 50892 3056 50948
rect 3112 50892 3180 50948
rect 3236 50892 3304 50948
rect 3360 50892 3428 50948
rect 3484 50892 3552 50948
rect 3608 50892 3676 50948
rect 3732 50892 3800 50948
rect 3856 50892 3924 50948
rect 3980 50892 4048 50948
rect 4104 50892 4172 50948
rect 4228 50892 4296 50948
rect 4352 50892 4420 50948
rect 4476 50892 4544 50948
rect 4600 50892 4668 50948
rect 4724 50892 4791 50948
rect 2741 50824 4791 50892
rect 2741 50768 2808 50824
rect 2864 50768 2932 50824
rect 2988 50768 3056 50824
rect 3112 50768 3180 50824
rect 3236 50768 3304 50824
rect 3360 50768 3428 50824
rect 3484 50768 3552 50824
rect 3608 50768 3676 50824
rect 3732 50768 3800 50824
rect 3856 50768 3924 50824
rect 3980 50768 4048 50824
rect 4104 50768 4172 50824
rect 4228 50768 4296 50824
rect 4352 50768 4420 50824
rect 4476 50768 4544 50824
rect 4600 50768 4668 50824
rect 4724 50768 4791 50824
rect 2741 50700 4791 50768
rect 2741 50644 2808 50700
rect 2864 50644 2932 50700
rect 2988 50644 3056 50700
rect 3112 50644 3180 50700
rect 3236 50644 3304 50700
rect 3360 50644 3428 50700
rect 3484 50644 3552 50700
rect 3608 50693 3676 50700
rect 3732 50693 3800 50700
rect 3856 50693 3924 50700
rect 3980 50693 4048 50700
rect 4104 50693 4172 50700
rect 4228 50693 4296 50700
rect 4352 50693 4420 50700
rect 4476 50693 4544 50700
rect 4600 50693 4668 50700
rect 4724 50693 4791 50700
rect 3611 50644 3676 50693
rect 3735 50644 3800 50693
rect 3859 50644 3924 50693
rect 3983 50644 4048 50693
rect 4107 50644 4172 50693
rect 4231 50644 4296 50693
rect 4355 50644 4420 50693
rect 4479 50644 4544 50693
rect 4603 50644 4668 50693
rect 2741 50641 3559 50644
rect 3611 50641 3683 50644
rect 3735 50641 3807 50644
rect 3859 50641 3931 50644
rect 3983 50641 4055 50644
rect 4107 50641 4179 50644
rect 4231 50641 4303 50644
rect 4355 50641 4427 50644
rect 4479 50641 4551 50644
rect 4603 50641 4675 50644
rect 4727 50641 4791 50693
rect 2741 50576 4791 50641
rect 2741 50520 2808 50576
rect 2864 50520 2932 50576
rect 2988 50520 3056 50576
rect 3112 50520 3180 50576
rect 3236 50520 3304 50576
rect 3360 50520 3428 50576
rect 3484 50520 3552 50576
rect 3608 50569 3676 50576
rect 3732 50569 3800 50576
rect 3856 50569 3924 50576
rect 3980 50569 4048 50576
rect 4104 50569 4172 50576
rect 4228 50569 4296 50576
rect 4352 50569 4420 50576
rect 4476 50569 4544 50576
rect 4600 50569 4668 50576
rect 4724 50569 4791 50576
rect 3611 50520 3676 50569
rect 3735 50520 3800 50569
rect 3859 50520 3924 50569
rect 3983 50520 4048 50569
rect 4107 50520 4172 50569
rect 4231 50520 4296 50569
rect 4355 50520 4420 50569
rect 4479 50520 4544 50569
rect 4603 50520 4668 50569
rect 2741 50517 3559 50520
rect 3611 50517 3683 50520
rect 3735 50517 3807 50520
rect 3859 50517 3931 50520
rect 3983 50517 4055 50520
rect 4107 50517 4179 50520
rect 4231 50517 4303 50520
rect 4355 50517 4427 50520
rect 4479 50517 4551 50520
rect 4603 50517 4675 50520
rect 4727 50517 4791 50569
rect 2741 50452 4791 50517
rect 2741 50396 2808 50452
rect 2864 50396 2932 50452
rect 2988 50396 3056 50452
rect 3112 50396 3180 50452
rect 3236 50396 3304 50452
rect 3360 50396 3428 50452
rect 3484 50396 3552 50452
rect 3608 50396 3676 50452
rect 3732 50396 3800 50452
rect 3856 50396 3924 50452
rect 3980 50396 4048 50452
rect 4104 50396 4172 50452
rect 4228 50396 4296 50452
rect 4352 50396 4420 50452
rect 4476 50396 4544 50452
rect 4600 50396 4668 50452
rect 4724 50396 4791 50452
rect 2741 50328 4791 50396
rect 2741 50272 2808 50328
rect 2864 50272 2932 50328
rect 2988 50272 3056 50328
rect 3112 50272 3180 50328
rect 3236 50272 3304 50328
rect 3360 50272 3428 50328
rect 3484 50272 3552 50328
rect 3608 50272 3676 50328
rect 3732 50272 3800 50328
rect 3856 50272 3924 50328
rect 3980 50272 4048 50328
rect 4104 50272 4172 50328
rect 4228 50272 4296 50328
rect 4352 50272 4420 50328
rect 4476 50272 4544 50328
rect 4600 50272 4668 50328
rect 4724 50272 4791 50328
rect 2741 50204 4791 50272
rect 2741 50148 2808 50204
rect 2864 50148 2932 50204
rect 2988 50148 3056 50204
rect 3112 50148 3180 50204
rect 3236 50148 3304 50204
rect 3360 50148 3428 50204
rect 3484 50148 3552 50204
rect 3608 50148 3676 50204
rect 3732 50148 3800 50204
rect 3856 50148 3924 50204
rect 3980 50148 4048 50204
rect 4104 50148 4172 50204
rect 4228 50148 4296 50204
rect 4352 50148 4420 50204
rect 4476 50148 4544 50204
rect 4600 50148 4668 50204
rect 4724 50148 4791 50204
rect 2741 50080 4791 50148
rect 2741 50024 2808 50080
rect 2864 50024 2932 50080
rect 2988 50024 3056 50080
rect 3112 50024 3180 50080
rect 3236 50024 3304 50080
rect 3360 50024 3428 50080
rect 3484 50024 3552 50080
rect 3608 50024 3676 50080
rect 3732 50024 3800 50080
rect 3856 50024 3924 50080
rect 3980 50024 4048 50080
rect 4104 50024 4172 50080
rect 4228 50024 4296 50080
rect 4352 50024 4420 50080
rect 4476 50024 4544 50080
rect 4600 50024 4668 50080
rect 4724 50024 4791 50080
rect 2741 49956 4791 50024
rect 2741 49900 2808 49956
rect 2864 49900 2932 49956
rect 2988 49900 3056 49956
rect 3112 49900 3180 49956
rect 3236 49900 3304 49956
rect 3360 49900 3428 49956
rect 3484 49900 3552 49956
rect 3608 49900 3676 49956
rect 3732 49900 3800 49956
rect 3856 49900 3924 49956
rect 3980 49900 4048 49956
rect 4104 49900 4172 49956
rect 4228 49900 4296 49956
rect 4352 49900 4420 49956
rect 4476 49900 4544 49956
rect 4600 49900 4668 49956
rect 4724 49900 4791 49956
rect 2741 49832 4791 49900
rect 2741 49776 2808 49832
rect 2864 49776 2932 49832
rect 2988 49776 3056 49832
rect 3112 49776 3180 49832
rect 3236 49776 3304 49832
rect 3360 49776 3428 49832
rect 3484 49776 3552 49832
rect 3608 49776 3676 49832
rect 3732 49776 3800 49832
rect 3856 49776 3924 49832
rect 3980 49776 4048 49832
rect 4104 49776 4172 49832
rect 4228 49776 4296 49832
rect 4352 49776 4420 49832
rect 4476 49776 4544 49832
rect 4600 49776 4668 49832
rect 4724 49776 4791 49832
rect 2741 49759 4791 49776
rect 2741 49708 3559 49759
rect 3611 49708 3683 49759
rect 3735 49708 3807 49759
rect 3859 49708 3931 49759
rect 3983 49708 4055 49759
rect 4107 49708 4179 49759
rect 4231 49708 4303 49759
rect 4355 49708 4427 49759
rect 4479 49708 4551 49759
rect 4603 49708 4675 49759
rect 2741 49652 2808 49708
rect 2864 49652 2932 49708
rect 2988 49652 3056 49708
rect 3112 49652 3180 49708
rect 3236 49652 3304 49708
rect 3360 49652 3428 49708
rect 3484 49652 3552 49708
rect 3611 49707 3676 49708
rect 3735 49707 3800 49708
rect 3859 49707 3924 49708
rect 3983 49707 4048 49708
rect 4107 49707 4172 49708
rect 4231 49707 4296 49708
rect 4355 49707 4420 49708
rect 4479 49707 4544 49708
rect 4603 49707 4668 49708
rect 4727 49707 4791 49759
rect 3608 49652 3676 49707
rect 3732 49652 3800 49707
rect 3856 49652 3924 49707
rect 3980 49652 4048 49707
rect 4104 49652 4172 49707
rect 4228 49652 4296 49707
rect 4352 49652 4420 49707
rect 4476 49652 4544 49707
rect 4600 49652 4668 49707
rect 4724 49652 4791 49707
rect 2741 49635 4791 49652
rect 2741 49583 3559 49635
rect 3611 49583 3683 49635
rect 3735 49583 3807 49635
rect 3859 49583 3931 49635
rect 3983 49583 4055 49635
rect 4107 49583 4179 49635
rect 4231 49583 4303 49635
rect 4355 49583 4427 49635
rect 4479 49583 4551 49635
rect 4603 49583 4675 49635
rect 4727 49583 4791 49635
rect 2741 48825 4791 49583
rect 2741 48773 3559 48825
rect 3611 48773 3683 48825
rect 3735 48773 3807 48825
rect 3859 48773 3931 48825
rect 3983 48773 4055 48825
rect 4107 48773 4179 48825
rect 4231 48773 4303 48825
rect 4355 48773 4427 48825
rect 4479 48773 4551 48825
rect 4603 48773 4675 48825
rect 4727 48773 4791 48825
rect 2741 48701 4791 48773
rect 2741 48649 3559 48701
rect 3611 48649 3683 48701
rect 3735 48649 3807 48701
rect 3859 48649 3931 48701
rect 3983 48649 4055 48701
rect 4107 48649 4179 48701
rect 4231 48649 4303 48701
rect 4355 48649 4427 48701
rect 4479 48649 4551 48701
rect 4603 48649 4675 48701
rect 4727 48649 4791 48701
rect 2741 47988 4791 48649
rect 2741 47936 2810 47988
rect 2862 47936 2934 47988
rect 2986 47936 3058 47988
rect 3110 47936 3182 47988
rect 3234 47936 3306 47988
rect 3358 47936 3430 47988
rect 3482 47936 3554 47988
rect 3606 47936 3678 47988
rect 3730 47936 3802 47988
rect 3854 47936 3926 47988
rect 3978 47936 4050 47988
rect 4102 47936 4174 47988
rect 4226 47936 4298 47988
rect 4350 47936 4422 47988
rect 4474 47936 4546 47988
rect 4598 47936 4670 47988
rect 4722 47936 4791 47988
rect 2741 47864 4791 47936
rect 2741 47812 2810 47864
rect 2862 47812 2934 47864
rect 2986 47812 3058 47864
rect 3110 47812 3182 47864
rect 3234 47812 3306 47864
rect 3358 47812 3430 47864
rect 3482 47812 3554 47864
rect 3606 47812 3678 47864
rect 3730 47812 3802 47864
rect 3854 47812 3926 47864
rect 3978 47812 4050 47864
rect 4102 47812 4174 47864
rect 4226 47812 4298 47864
rect 4350 47812 4422 47864
rect 4474 47812 4546 47864
rect 4598 47812 4670 47864
rect 4722 47812 4791 47864
rect 2741 47740 4791 47812
rect 2741 47688 2810 47740
rect 2862 47688 2934 47740
rect 2986 47688 3058 47740
rect 3110 47688 3182 47740
rect 3234 47688 3306 47740
rect 3358 47688 3430 47740
rect 3482 47688 3554 47740
rect 3606 47688 3678 47740
rect 3730 47688 3802 47740
rect 3854 47688 3926 47740
rect 3978 47688 4050 47740
rect 4102 47688 4174 47740
rect 4226 47688 4298 47740
rect 4350 47688 4422 47740
rect 4474 47688 4546 47740
rect 4598 47688 4670 47740
rect 4722 47688 4791 47740
rect 2741 46430 4791 47688
rect 4851 57108 5051 57278
rect 4851 57056 4871 57108
rect 4923 57056 4979 57108
rect 5031 57056 5051 57108
rect 4851 53484 5051 57056
rect 4851 53432 4871 53484
rect 4923 53432 4979 53484
rect 5031 53432 5051 53484
rect 4851 53376 5051 53432
rect 4851 53324 4871 53376
rect 4923 53324 4979 53376
rect 5031 53324 5051 53376
rect 4851 53268 5051 53324
rect 4851 53216 4871 53268
rect 4923 53216 4979 53268
rect 5031 53216 5051 53268
rect 4851 52548 5051 53216
rect 4851 52492 4861 52548
rect 4917 52492 4985 52548
rect 5041 52492 5051 52548
rect 4851 52424 5051 52492
rect 4851 52368 4861 52424
rect 4917 52368 4985 52424
rect 5041 52368 5051 52424
rect 4851 52300 5051 52368
rect 4851 52244 4861 52300
rect 4917 52244 4985 52300
rect 5041 52244 5051 52300
rect 4851 52176 5051 52244
rect 4851 52120 4861 52176
rect 4917 52120 4985 52176
rect 5041 52120 5051 52176
rect 4851 52052 5051 52120
rect 4851 51996 4861 52052
rect 4917 51996 4985 52052
rect 5041 51996 5051 52052
rect 4851 51965 4863 51996
rect 4915 51965 4987 51996
rect 5039 51965 5051 51996
rect 4851 51928 5051 51965
rect 4851 51872 4861 51928
rect 4917 51872 4985 51928
rect 5041 51872 5051 51928
rect 4851 51841 4863 51872
rect 4915 51841 4987 51872
rect 5039 51841 5051 51872
rect 4851 51804 5051 51841
rect 4851 51748 4861 51804
rect 4917 51748 4985 51804
rect 5041 51748 5051 51804
rect 4851 51680 5051 51748
rect 4851 51624 4861 51680
rect 4917 51624 4985 51680
rect 5041 51624 5051 51680
rect 4851 51556 5051 51624
rect 4851 51500 4861 51556
rect 4917 51500 4985 51556
rect 5041 51500 5051 51556
rect 4851 51432 5051 51500
rect 4851 51376 4861 51432
rect 4917 51376 4985 51432
rect 5041 51376 5051 51432
rect 4851 51308 5051 51376
rect 4851 51252 4861 51308
rect 4917 51252 4985 51308
rect 5041 51252 5051 51308
rect 4851 51222 5051 51252
rect 4851 51170 4863 51222
rect 4915 51170 4987 51222
rect 5039 51170 5051 51222
rect 4851 51098 5051 51170
rect 4851 51046 4863 51098
rect 4915 51046 4987 51098
rect 5039 51046 5051 51098
rect 4851 50974 5051 51046
rect 4851 50922 4863 50974
rect 4915 50922 4987 50974
rect 5039 50922 5051 50974
rect 4851 50288 5051 50922
rect 4851 50236 4863 50288
rect 4915 50236 4987 50288
rect 5039 50236 5051 50288
rect 4851 50164 5051 50236
rect 4851 50112 4863 50164
rect 4915 50112 4987 50164
rect 5039 50112 5051 50164
rect 4851 50040 5051 50112
rect 4851 49988 4863 50040
rect 4915 49988 4987 50040
rect 5039 49988 5051 50040
rect 4851 49354 5051 49988
rect 4851 49302 4863 49354
rect 4915 49302 4987 49354
rect 5039 49302 5051 49354
rect 4851 49230 5051 49302
rect 4851 49178 4863 49230
rect 4915 49178 4987 49230
rect 5039 49178 5051 49230
rect 4851 49106 5051 49178
rect 4851 49054 4863 49106
rect 4915 49054 4987 49106
rect 5039 49054 5051 49106
rect 4851 48435 5051 49054
rect 4851 48383 4863 48435
rect 4915 48383 4987 48435
rect 5039 48383 5051 48435
rect 4851 48311 5051 48383
rect 4851 48259 4863 48311
rect 4915 48259 4987 48311
rect 5039 48259 5051 48311
rect 4851 46430 5051 48259
rect 5111 56669 7161 57600
rect 5111 56617 6297 56669
rect 6349 56617 6421 56669
rect 6473 56617 6545 56669
rect 6597 56617 6669 56669
rect 6721 56617 6793 56669
rect 6845 56617 6917 56669
rect 6969 56617 7041 56669
rect 7093 56617 7161 56669
rect 5111 56545 7161 56617
rect 5111 56493 6297 56545
rect 6349 56493 6421 56545
rect 6473 56493 6545 56545
rect 6597 56493 6669 56545
rect 6721 56493 6793 56545
rect 6845 56493 6917 56545
rect 6969 56493 7041 56545
rect 7093 56493 7161 56545
rect 5111 56421 7161 56493
rect 5111 56369 6297 56421
rect 6349 56369 6421 56421
rect 6473 56369 6545 56421
rect 6597 56369 6669 56421
rect 6721 56369 6793 56421
rect 6845 56369 6917 56421
rect 6969 56369 7041 56421
rect 7093 56369 7161 56421
rect 5111 56297 7161 56369
rect 5111 56245 6297 56297
rect 6349 56245 6421 56297
rect 6473 56245 6545 56297
rect 6597 56245 6669 56297
rect 6721 56245 6793 56297
rect 6845 56245 6917 56297
rect 6969 56245 7041 56297
rect 7093 56245 7161 56297
rect 5111 56173 7161 56245
rect 5111 56121 6297 56173
rect 6349 56121 6421 56173
rect 6473 56121 6545 56173
rect 6597 56121 6669 56173
rect 6721 56121 6793 56173
rect 6845 56121 6917 56173
rect 6969 56121 7041 56173
rect 7093 56121 7161 56173
rect 5111 56049 7161 56121
rect 5111 55997 6297 56049
rect 6349 55997 6421 56049
rect 6473 55997 6545 56049
rect 6597 55997 6669 56049
rect 6721 55997 6793 56049
rect 6845 55997 6917 56049
rect 6969 55997 7041 56049
rect 7093 55997 7161 56049
rect 5111 55925 7161 55997
rect 5111 55873 6297 55925
rect 6349 55873 6421 55925
rect 6473 55873 6545 55925
rect 6597 55873 6669 55925
rect 6721 55873 6793 55925
rect 6845 55873 6917 55925
rect 6969 55873 7041 55925
rect 7093 55873 7161 55925
rect 5111 55801 7161 55873
rect 5111 55749 6297 55801
rect 6349 55749 6421 55801
rect 6473 55749 6545 55801
rect 6597 55749 6669 55801
rect 6721 55749 6793 55801
rect 6845 55749 6917 55801
rect 6969 55749 7041 55801
rect 7093 55749 7161 55801
rect 5111 55677 7161 55749
rect 5111 55625 6297 55677
rect 6349 55625 6421 55677
rect 6473 55625 6545 55677
rect 6597 55625 6669 55677
rect 6721 55625 6793 55677
rect 6845 55625 6917 55677
rect 6969 55625 7041 55677
rect 7093 55625 7161 55677
rect 5111 55553 7161 55625
rect 5111 55501 6297 55553
rect 6349 55501 6421 55553
rect 6473 55501 6545 55553
rect 6597 55501 6669 55553
rect 6721 55501 6793 55553
rect 6845 55501 6917 55553
rect 6969 55501 7041 55553
rect 7093 55501 7161 55553
rect 5111 55429 7161 55501
rect 5111 55377 6297 55429
rect 6349 55377 6421 55429
rect 6473 55377 6545 55429
rect 6597 55377 6669 55429
rect 6721 55377 6793 55429
rect 6845 55377 6917 55429
rect 6969 55377 7041 55429
rect 7093 55377 7161 55429
rect 5111 55305 7161 55377
rect 5111 55253 6297 55305
rect 6349 55253 6421 55305
rect 6473 55253 6545 55305
rect 6597 55253 6669 55305
rect 6721 55253 6793 55305
rect 6845 55253 6917 55305
rect 6969 55253 7041 55305
rect 7093 55253 7161 55305
rect 5111 55181 7161 55253
rect 5111 55129 6297 55181
rect 6349 55129 6421 55181
rect 6473 55129 6545 55181
rect 6597 55129 6669 55181
rect 6721 55129 6793 55181
rect 6845 55129 6917 55181
rect 6969 55129 7041 55181
rect 7093 55129 7161 55181
rect 5111 55057 7161 55129
rect 5111 55005 6297 55057
rect 6349 55005 6421 55057
rect 6473 55005 6545 55057
rect 6597 55005 6669 55057
rect 6721 55005 6793 55057
rect 6845 55005 6917 55057
rect 6969 55005 7041 55057
rect 7093 55005 7161 55057
rect 5111 54933 7161 55005
rect 5111 54881 6297 54933
rect 6349 54881 6421 54933
rect 6473 54881 6545 54933
rect 6597 54881 6669 54933
rect 6721 54881 6793 54933
rect 6845 54881 6917 54933
rect 6969 54881 7041 54933
rect 7093 54881 7161 54933
rect 5111 54809 7161 54881
rect 5111 54757 6297 54809
rect 6349 54757 6421 54809
rect 6473 54757 6545 54809
rect 6597 54757 6669 54809
rect 6721 54757 6793 54809
rect 6845 54757 6917 54809
rect 6969 54757 7041 54809
rect 7093 54757 7161 54809
rect 5111 54685 7161 54757
rect 5111 54633 6297 54685
rect 6349 54633 6421 54685
rect 6473 54633 6545 54685
rect 6597 54633 6669 54685
rect 6721 54633 6793 54685
rect 6845 54633 6917 54685
rect 6969 54633 7041 54685
rect 7093 54633 7161 54685
rect 5111 54561 7161 54633
rect 5111 54509 6297 54561
rect 6349 54509 6421 54561
rect 6473 54509 6545 54561
rect 6597 54509 6669 54561
rect 6721 54509 6793 54561
rect 6845 54509 6917 54561
rect 6969 54509 7041 54561
rect 7093 54509 7161 54561
rect 5111 54437 7161 54509
rect 5111 54385 6297 54437
rect 6349 54385 6421 54437
rect 6473 54385 6545 54437
rect 6597 54385 6669 54437
rect 6721 54385 6793 54437
rect 6845 54385 6917 54437
rect 6969 54385 7041 54437
rect 7093 54385 7161 54437
rect 5111 54313 7161 54385
rect 5111 54261 6297 54313
rect 6349 54261 6421 54313
rect 6473 54261 6545 54313
rect 6597 54261 6669 54313
rect 6721 54261 6793 54313
rect 6845 54261 6917 54313
rect 6969 54261 7041 54313
rect 7093 54261 7161 54313
rect 5111 54189 7161 54261
rect 5111 54137 6297 54189
rect 6349 54137 6421 54189
rect 6473 54137 6545 54189
rect 6597 54137 6669 54189
rect 6721 54137 6793 54189
rect 6845 54137 6917 54189
rect 6969 54137 7041 54189
rect 7093 54137 7161 54189
rect 5111 54065 7161 54137
rect 5111 54013 6297 54065
rect 6349 54013 6421 54065
rect 6473 54013 6545 54065
rect 6597 54013 6669 54065
rect 6721 54013 6793 54065
rect 6845 54013 6917 54065
rect 6969 54013 7041 54065
rect 7093 54013 7161 54065
rect 5111 53941 7161 54013
rect 5111 53889 6297 53941
rect 6349 53889 6421 53941
rect 6473 53889 6545 53941
rect 6597 53889 6669 53941
rect 6721 53889 6793 53941
rect 6845 53889 6917 53941
rect 6969 53889 7041 53941
rect 7093 53889 7161 53941
rect 5111 53817 7161 53889
rect 5111 53765 6297 53817
rect 6349 53765 6421 53817
rect 6473 53765 6545 53817
rect 6597 53765 6669 53817
rect 6721 53765 6793 53817
rect 6845 53765 6917 53817
rect 6969 53765 7041 53817
rect 7093 53765 7161 53817
rect 5111 53693 7161 53765
rect 5111 53641 6297 53693
rect 6349 53641 6421 53693
rect 6473 53641 6545 53693
rect 6597 53641 6669 53693
rect 6721 53641 6793 53693
rect 6845 53641 6917 53693
rect 6969 53641 7041 53693
rect 7093 53641 7161 53693
rect 5111 52588 7161 53641
rect 5111 52536 5180 52588
rect 5232 52536 5304 52588
rect 5356 52536 5428 52588
rect 5480 52536 5552 52588
rect 5604 52536 5676 52588
rect 5728 52536 5800 52588
rect 5852 52536 5924 52588
rect 5976 52536 6048 52588
rect 6100 52536 6172 52588
rect 6224 52536 6296 52588
rect 6348 52536 6420 52588
rect 6472 52536 6544 52588
rect 6596 52536 6668 52588
rect 6720 52536 6792 52588
rect 6844 52536 6916 52588
rect 6968 52536 7040 52588
rect 7092 52536 7161 52588
rect 5111 52464 7161 52536
rect 5111 52412 5180 52464
rect 5232 52412 5304 52464
rect 5356 52412 5428 52464
rect 5480 52412 5552 52464
rect 5604 52412 5676 52464
rect 5728 52412 5800 52464
rect 5852 52412 5924 52464
rect 5976 52412 6048 52464
rect 6100 52412 6172 52464
rect 6224 52412 6296 52464
rect 6348 52412 6420 52464
rect 6472 52412 6544 52464
rect 6596 52412 6668 52464
rect 6720 52412 6792 52464
rect 6844 52412 6916 52464
rect 6968 52412 7040 52464
rect 7092 52412 7161 52464
rect 5111 52340 7161 52412
rect 5111 52288 5180 52340
rect 5232 52288 5304 52340
rect 5356 52288 5428 52340
rect 5480 52288 5552 52340
rect 5604 52288 5676 52340
rect 5728 52288 5800 52340
rect 5852 52288 5924 52340
rect 5976 52288 6048 52340
rect 6100 52288 6172 52340
rect 6224 52288 6296 52340
rect 6348 52288 6420 52340
rect 6472 52288 6544 52340
rect 6596 52288 6668 52340
rect 6720 52288 6792 52340
rect 6844 52288 6916 52340
rect 6968 52288 7040 52340
rect 7092 52288 7161 52340
rect 5111 51627 7161 52288
rect 5111 51575 5180 51627
rect 5232 51575 5304 51627
rect 5356 51575 5428 51627
rect 5480 51575 5552 51627
rect 5604 51575 5676 51627
rect 5728 51575 5800 51627
rect 5852 51575 5924 51627
rect 5976 51575 6048 51627
rect 6100 51575 6172 51627
rect 6224 51575 6296 51627
rect 6348 51575 6420 51627
rect 6472 51575 6544 51627
rect 6596 51575 6668 51627
rect 6720 51575 6792 51627
rect 6844 51575 6916 51627
rect 6968 51575 7040 51627
rect 7092 51575 7161 51627
rect 5111 51503 7161 51575
rect 5111 51451 5180 51503
rect 5232 51451 5304 51503
rect 5356 51451 5428 51503
rect 5480 51451 5552 51503
rect 5604 51451 5676 51503
rect 5728 51451 5800 51503
rect 5852 51451 5924 51503
rect 5976 51451 6048 51503
rect 6100 51451 6172 51503
rect 6224 51451 6296 51503
rect 6348 51451 6420 51503
rect 6472 51451 6544 51503
rect 6596 51451 6668 51503
rect 6720 51451 6792 51503
rect 6844 51451 6916 51503
rect 6968 51451 7040 51503
rect 7092 51451 7161 51503
rect 5111 50948 7161 51451
rect 5111 50892 5178 50948
rect 5234 50892 5302 50948
rect 5358 50892 5426 50948
rect 5482 50892 5550 50948
rect 5606 50892 5674 50948
rect 5730 50892 5798 50948
rect 5854 50892 5922 50948
rect 5978 50892 6046 50948
rect 6102 50892 6170 50948
rect 6226 50892 6294 50948
rect 6350 50892 6418 50948
rect 6474 50892 6542 50948
rect 6598 50892 6666 50948
rect 6722 50892 6790 50948
rect 6846 50892 6914 50948
rect 6970 50892 7038 50948
rect 7094 50892 7161 50948
rect 5111 50824 7161 50892
rect 5111 50768 5178 50824
rect 5234 50768 5302 50824
rect 5358 50768 5426 50824
rect 5482 50768 5550 50824
rect 5606 50768 5674 50824
rect 5730 50768 5798 50824
rect 5854 50768 5922 50824
rect 5978 50768 6046 50824
rect 6102 50768 6170 50824
rect 6226 50768 6294 50824
rect 6350 50768 6418 50824
rect 6474 50768 6542 50824
rect 6598 50768 6666 50824
rect 6722 50768 6790 50824
rect 6846 50768 6914 50824
rect 6970 50768 7038 50824
rect 7094 50768 7161 50824
rect 5111 50700 7161 50768
rect 5111 50644 5178 50700
rect 5234 50644 5302 50700
rect 5358 50644 5426 50700
rect 5482 50644 5550 50700
rect 5606 50644 5674 50700
rect 5730 50644 5798 50700
rect 5854 50644 5922 50700
rect 5978 50644 6046 50700
rect 6102 50644 6170 50700
rect 6226 50644 6294 50700
rect 6350 50644 6418 50700
rect 6474 50644 6542 50700
rect 6598 50644 6666 50700
rect 6722 50644 6790 50700
rect 6846 50644 6914 50700
rect 6970 50644 7038 50700
rect 7094 50644 7161 50700
rect 5111 50641 5180 50644
rect 5232 50641 5304 50644
rect 5356 50641 5428 50644
rect 5480 50641 5552 50644
rect 5604 50641 5676 50644
rect 5728 50641 5800 50644
rect 5852 50641 5924 50644
rect 5976 50641 6048 50644
rect 6100 50641 6172 50644
rect 6224 50641 6296 50644
rect 6348 50641 6420 50644
rect 6472 50641 6544 50644
rect 6596 50641 6668 50644
rect 6720 50641 6792 50644
rect 6844 50641 6916 50644
rect 6968 50641 7040 50644
rect 7092 50641 7161 50644
rect 5111 50576 7161 50641
rect 5111 50520 5178 50576
rect 5234 50520 5302 50576
rect 5358 50520 5426 50576
rect 5482 50520 5550 50576
rect 5606 50520 5674 50576
rect 5730 50520 5798 50576
rect 5854 50520 5922 50576
rect 5978 50520 6046 50576
rect 6102 50520 6170 50576
rect 6226 50520 6294 50576
rect 6350 50520 6418 50576
rect 6474 50520 6542 50576
rect 6598 50520 6666 50576
rect 6722 50520 6790 50576
rect 6846 50520 6914 50576
rect 6970 50520 7038 50576
rect 7094 50520 7161 50576
rect 5111 50517 5180 50520
rect 5232 50517 5304 50520
rect 5356 50517 5428 50520
rect 5480 50517 5552 50520
rect 5604 50517 5676 50520
rect 5728 50517 5800 50520
rect 5852 50517 5924 50520
rect 5976 50517 6048 50520
rect 6100 50517 6172 50520
rect 6224 50517 6296 50520
rect 6348 50517 6420 50520
rect 6472 50517 6544 50520
rect 6596 50517 6668 50520
rect 6720 50517 6792 50520
rect 6844 50517 6916 50520
rect 6968 50517 7040 50520
rect 7092 50517 7161 50520
rect 5111 50452 7161 50517
rect 5111 50396 5178 50452
rect 5234 50396 5302 50452
rect 5358 50396 5426 50452
rect 5482 50396 5550 50452
rect 5606 50396 5674 50452
rect 5730 50396 5798 50452
rect 5854 50396 5922 50452
rect 5978 50396 6046 50452
rect 6102 50396 6170 50452
rect 6226 50396 6294 50452
rect 6350 50396 6418 50452
rect 6474 50396 6542 50452
rect 6598 50396 6666 50452
rect 6722 50396 6790 50452
rect 6846 50396 6914 50452
rect 6970 50396 7038 50452
rect 7094 50396 7161 50452
rect 5111 50328 7161 50396
rect 5111 50272 5178 50328
rect 5234 50272 5302 50328
rect 5358 50272 5426 50328
rect 5482 50272 5550 50328
rect 5606 50272 5674 50328
rect 5730 50272 5798 50328
rect 5854 50272 5922 50328
rect 5978 50272 6046 50328
rect 6102 50272 6170 50328
rect 6226 50272 6294 50328
rect 6350 50272 6418 50328
rect 6474 50272 6542 50328
rect 6598 50272 6666 50328
rect 6722 50272 6790 50328
rect 6846 50272 6914 50328
rect 6970 50272 7038 50328
rect 7094 50272 7161 50328
rect 5111 50204 7161 50272
rect 5111 50148 5178 50204
rect 5234 50148 5302 50204
rect 5358 50148 5426 50204
rect 5482 50148 5550 50204
rect 5606 50148 5674 50204
rect 5730 50148 5798 50204
rect 5854 50148 5922 50204
rect 5978 50148 6046 50204
rect 6102 50148 6170 50204
rect 6226 50148 6294 50204
rect 6350 50148 6418 50204
rect 6474 50148 6542 50204
rect 6598 50148 6666 50204
rect 6722 50148 6790 50204
rect 6846 50148 6914 50204
rect 6970 50148 7038 50204
rect 7094 50148 7161 50204
rect 5111 50080 7161 50148
rect 5111 50024 5178 50080
rect 5234 50024 5302 50080
rect 5358 50024 5426 50080
rect 5482 50024 5550 50080
rect 5606 50024 5674 50080
rect 5730 50024 5798 50080
rect 5854 50024 5922 50080
rect 5978 50024 6046 50080
rect 6102 50024 6170 50080
rect 6226 50024 6294 50080
rect 6350 50024 6418 50080
rect 6474 50024 6542 50080
rect 6598 50024 6666 50080
rect 6722 50024 6790 50080
rect 6846 50024 6914 50080
rect 6970 50024 7038 50080
rect 7094 50024 7161 50080
rect 5111 49956 7161 50024
rect 5111 49900 5178 49956
rect 5234 49900 5302 49956
rect 5358 49900 5426 49956
rect 5482 49900 5550 49956
rect 5606 49900 5674 49956
rect 5730 49900 5798 49956
rect 5854 49900 5922 49956
rect 5978 49900 6046 49956
rect 6102 49900 6170 49956
rect 6226 49900 6294 49956
rect 6350 49900 6418 49956
rect 6474 49900 6542 49956
rect 6598 49900 6666 49956
rect 6722 49900 6790 49956
rect 6846 49900 6914 49956
rect 6970 49900 7038 49956
rect 7094 49900 7161 49956
rect 5111 49832 7161 49900
rect 5111 49776 5178 49832
rect 5234 49776 5302 49832
rect 5358 49776 5426 49832
rect 5482 49776 5550 49832
rect 5606 49776 5674 49832
rect 5730 49776 5798 49832
rect 5854 49776 5922 49832
rect 5978 49776 6046 49832
rect 6102 49776 6170 49832
rect 6226 49776 6294 49832
rect 6350 49776 6418 49832
rect 6474 49776 6542 49832
rect 6598 49776 6666 49832
rect 6722 49776 6790 49832
rect 6846 49776 6914 49832
rect 6970 49776 7038 49832
rect 7094 49776 7161 49832
rect 5111 49759 7161 49776
rect 5111 49708 5180 49759
rect 5232 49708 5304 49759
rect 5356 49708 5428 49759
rect 5480 49708 5552 49759
rect 5604 49708 5676 49759
rect 5728 49708 5800 49759
rect 5852 49708 5924 49759
rect 5976 49708 6048 49759
rect 6100 49708 6172 49759
rect 6224 49708 6296 49759
rect 6348 49708 6420 49759
rect 6472 49708 6544 49759
rect 6596 49708 6668 49759
rect 6720 49708 6792 49759
rect 6844 49708 6916 49759
rect 6968 49708 7040 49759
rect 7092 49708 7161 49759
rect 5111 49652 5178 49708
rect 5234 49652 5302 49708
rect 5358 49652 5426 49708
rect 5482 49652 5550 49708
rect 5606 49652 5674 49708
rect 5730 49652 5798 49708
rect 5854 49652 5922 49708
rect 5978 49652 6046 49708
rect 6102 49652 6170 49708
rect 6226 49652 6294 49708
rect 6350 49652 6418 49708
rect 6474 49652 6542 49708
rect 6598 49652 6666 49708
rect 6722 49652 6790 49708
rect 6846 49652 6914 49708
rect 6970 49652 7038 49708
rect 7094 49652 7161 49708
rect 5111 49635 7161 49652
rect 5111 49583 5180 49635
rect 5232 49583 5304 49635
rect 5356 49583 5428 49635
rect 5480 49583 5552 49635
rect 5604 49583 5676 49635
rect 5728 49583 5800 49635
rect 5852 49583 5924 49635
rect 5976 49583 6048 49635
rect 6100 49583 6172 49635
rect 6224 49583 6296 49635
rect 6348 49583 6420 49635
rect 6472 49583 6544 49635
rect 6596 49583 6668 49635
rect 6720 49583 6792 49635
rect 6844 49583 6916 49635
rect 6968 49583 7040 49635
rect 7092 49583 7161 49635
rect 5111 48825 7161 49583
rect 5111 48773 5180 48825
rect 5232 48773 5304 48825
rect 5356 48773 5428 48825
rect 5480 48773 5552 48825
rect 5604 48773 5676 48825
rect 5728 48773 5800 48825
rect 5852 48773 5924 48825
rect 5976 48773 6048 48825
rect 6100 48773 6172 48825
rect 6224 48773 6296 48825
rect 6348 48773 6420 48825
rect 6472 48773 6544 48825
rect 6596 48773 6668 48825
rect 6720 48773 6792 48825
rect 6844 48773 6916 48825
rect 6968 48773 7040 48825
rect 7092 48773 7161 48825
rect 5111 48701 7161 48773
rect 5111 48649 5180 48701
rect 5232 48649 5304 48701
rect 5356 48649 5428 48701
rect 5480 48649 5552 48701
rect 5604 48649 5676 48701
rect 5728 48649 5800 48701
rect 5852 48649 5924 48701
rect 5976 48649 6048 48701
rect 6100 48649 6172 48701
rect 6224 48649 6296 48701
rect 6348 48649 6420 48701
rect 6472 48649 6544 48701
rect 6596 48649 6668 48701
rect 6720 48649 6792 48701
rect 6844 48649 6916 48701
rect 6968 48649 7040 48701
rect 7092 48649 7161 48701
rect 5111 47988 7161 48649
rect 5111 47936 5180 47988
rect 5232 47936 5304 47988
rect 5356 47936 5428 47988
rect 5480 47936 5552 47988
rect 5604 47936 5676 47988
rect 5728 47936 5800 47988
rect 5852 47936 5924 47988
rect 5976 47936 6048 47988
rect 6100 47936 6172 47988
rect 6224 47936 6296 47988
rect 6348 47936 6420 47988
rect 6472 47936 6544 47988
rect 6596 47936 6668 47988
rect 6720 47936 6792 47988
rect 6844 47936 6916 47988
rect 6968 47936 7040 47988
rect 7092 47936 7161 47988
rect 5111 47864 7161 47936
rect 5111 47812 5180 47864
rect 5232 47812 5304 47864
rect 5356 47812 5428 47864
rect 5480 47812 5552 47864
rect 5604 47812 5676 47864
rect 5728 47812 5800 47864
rect 5852 47812 5924 47864
rect 5976 47812 6048 47864
rect 6100 47812 6172 47864
rect 6224 47812 6296 47864
rect 6348 47812 6420 47864
rect 6472 47812 6544 47864
rect 6596 47812 6668 47864
rect 6720 47812 6792 47864
rect 6844 47812 6916 47864
rect 6968 47812 7040 47864
rect 7092 47812 7161 47864
rect 5111 47740 7161 47812
rect 5111 47688 5180 47740
rect 5232 47688 5304 47740
rect 5356 47688 5428 47740
rect 5480 47688 5552 47740
rect 5604 47688 5676 47740
rect 5728 47688 5800 47740
rect 5852 47688 5924 47740
rect 5976 47688 6048 47740
rect 6100 47688 6172 47740
rect 6224 47688 6296 47740
rect 6348 47688 6420 47740
rect 6472 47688 6544 47740
rect 6596 47688 6668 47740
rect 6720 47688 6792 47740
rect 6844 47688 6916 47740
rect 6968 47688 7040 47740
rect 7092 47688 7161 47740
rect 5111 46430 7161 47688
rect 7221 57108 7757 57278
rect 7221 57056 7247 57108
rect 7299 57056 7355 57108
rect 7407 57056 7463 57108
rect 7515 57056 7571 57108
rect 7623 57056 7679 57108
rect 7731 57056 7757 57108
rect 7221 53484 7757 57056
rect 7221 53432 7247 53484
rect 7299 53432 7355 53484
rect 7407 53432 7463 53484
rect 7515 53432 7571 53484
rect 7623 53432 7679 53484
rect 7731 53432 7757 53484
rect 7221 53376 7757 53432
rect 7221 53324 7247 53376
rect 7299 53324 7355 53376
rect 7407 53324 7463 53376
rect 7515 53324 7571 53376
rect 7623 53324 7679 53376
rect 7731 53324 7757 53376
rect 7221 53268 7757 53324
rect 7221 53216 7247 53268
rect 7299 53216 7355 53268
rect 7407 53216 7463 53268
rect 7515 53216 7571 53268
rect 7623 53216 7679 53268
rect 7731 53216 7757 53268
rect 7221 52548 7757 53216
rect 7221 52492 7275 52548
rect 7331 52492 7399 52548
rect 7455 52492 7523 52548
rect 7579 52492 7647 52548
rect 7703 52492 7757 52548
rect 7221 52424 7757 52492
rect 7221 52368 7275 52424
rect 7331 52368 7399 52424
rect 7455 52368 7523 52424
rect 7579 52368 7647 52424
rect 7703 52368 7757 52424
rect 7221 52300 7757 52368
rect 7221 52244 7275 52300
rect 7331 52244 7399 52300
rect 7455 52244 7523 52300
rect 7579 52244 7647 52300
rect 7703 52244 7757 52300
rect 7221 52176 7757 52244
rect 7221 52120 7275 52176
rect 7331 52120 7399 52176
rect 7455 52120 7523 52176
rect 7579 52120 7647 52176
rect 7703 52120 7757 52176
rect 7221 52052 7757 52120
rect 7221 51996 7275 52052
rect 7331 51996 7399 52052
rect 7455 51996 7523 52052
rect 7579 51996 7647 52052
rect 7703 51996 7757 52052
rect 7221 51965 7277 51996
rect 7329 51965 7401 51996
rect 7453 51965 7525 51996
rect 7577 51965 7649 51996
rect 7701 51965 7757 51996
rect 7221 51928 7757 51965
rect 7221 51872 7275 51928
rect 7331 51872 7399 51928
rect 7455 51872 7523 51928
rect 7579 51872 7647 51928
rect 7703 51872 7757 51928
rect 7221 51841 7277 51872
rect 7329 51841 7401 51872
rect 7453 51841 7525 51872
rect 7577 51841 7649 51872
rect 7701 51841 7757 51872
rect 7221 51804 7757 51841
rect 7221 51748 7275 51804
rect 7331 51748 7399 51804
rect 7455 51748 7523 51804
rect 7579 51748 7647 51804
rect 7703 51748 7757 51804
rect 7221 51680 7757 51748
rect 7221 51624 7275 51680
rect 7331 51624 7399 51680
rect 7455 51624 7523 51680
rect 7579 51624 7647 51680
rect 7703 51624 7757 51680
rect 7221 51556 7757 51624
rect 7221 51500 7275 51556
rect 7331 51500 7399 51556
rect 7455 51500 7523 51556
rect 7579 51500 7647 51556
rect 7703 51500 7757 51556
rect 7221 51432 7757 51500
rect 7221 51376 7275 51432
rect 7331 51376 7399 51432
rect 7455 51376 7523 51432
rect 7579 51376 7647 51432
rect 7703 51376 7757 51432
rect 7221 51308 7757 51376
rect 7221 51252 7275 51308
rect 7331 51252 7399 51308
rect 7455 51252 7523 51308
rect 7579 51252 7647 51308
rect 7703 51252 7757 51308
rect 7221 51222 7757 51252
rect 7221 51170 7277 51222
rect 7329 51170 7401 51222
rect 7453 51170 7525 51222
rect 7577 51170 7649 51222
rect 7701 51170 7757 51222
rect 7221 51098 7757 51170
rect 7221 51046 7277 51098
rect 7329 51046 7401 51098
rect 7453 51046 7525 51098
rect 7577 51046 7649 51098
rect 7701 51046 7757 51098
rect 7221 50974 7757 51046
rect 7221 50922 7277 50974
rect 7329 50922 7401 50974
rect 7453 50922 7525 50974
rect 7577 50922 7649 50974
rect 7701 50922 7757 50974
rect 7221 50288 7757 50922
rect 7221 50236 7277 50288
rect 7329 50236 7401 50288
rect 7453 50236 7525 50288
rect 7577 50236 7649 50288
rect 7701 50236 7757 50288
rect 7221 50164 7757 50236
rect 7221 50112 7277 50164
rect 7329 50112 7401 50164
rect 7453 50112 7525 50164
rect 7577 50112 7649 50164
rect 7701 50112 7757 50164
rect 7221 50040 7757 50112
rect 7221 49988 7277 50040
rect 7329 49988 7401 50040
rect 7453 49988 7525 50040
rect 7577 49988 7649 50040
rect 7701 49988 7757 50040
rect 7221 49354 7757 49988
rect 7221 49302 7277 49354
rect 7329 49302 7401 49354
rect 7453 49302 7525 49354
rect 7577 49302 7649 49354
rect 7701 49302 7757 49354
rect 7221 49230 7757 49302
rect 7221 49178 7277 49230
rect 7329 49178 7401 49230
rect 7453 49178 7525 49230
rect 7577 49178 7649 49230
rect 7701 49178 7757 49230
rect 7221 49106 7757 49178
rect 7221 49054 7277 49106
rect 7329 49054 7401 49106
rect 7453 49054 7525 49106
rect 7577 49054 7649 49106
rect 7701 49054 7757 49106
rect 7221 48435 7757 49054
rect 7221 48383 7277 48435
rect 7329 48383 7401 48435
rect 7453 48383 7525 48435
rect 7577 48383 7649 48435
rect 7701 48383 7757 48435
rect 7221 48311 7757 48383
rect 7221 48259 7277 48311
rect 7329 48259 7401 48311
rect 7453 48259 7525 48311
rect 7577 48259 7649 48311
rect 7701 48259 7757 48311
rect 7221 46430 7757 48259
rect 7817 56669 9867 57600
rect 7817 56617 7885 56669
rect 7937 56617 8009 56669
rect 8061 56617 8133 56669
rect 8185 56617 8257 56669
rect 8309 56617 8381 56669
rect 8433 56617 8505 56669
rect 8557 56617 8629 56669
rect 8681 56617 9867 56669
rect 7817 56545 9867 56617
rect 7817 56493 7885 56545
rect 7937 56493 8009 56545
rect 8061 56493 8133 56545
rect 8185 56493 8257 56545
rect 8309 56493 8381 56545
rect 8433 56493 8505 56545
rect 8557 56493 8629 56545
rect 8681 56493 9867 56545
rect 7817 56421 9867 56493
rect 7817 56369 7885 56421
rect 7937 56369 8009 56421
rect 8061 56369 8133 56421
rect 8185 56369 8257 56421
rect 8309 56369 8381 56421
rect 8433 56369 8505 56421
rect 8557 56369 8629 56421
rect 8681 56369 9867 56421
rect 7817 56297 9867 56369
rect 7817 56245 7885 56297
rect 7937 56245 8009 56297
rect 8061 56245 8133 56297
rect 8185 56245 8257 56297
rect 8309 56245 8381 56297
rect 8433 56245 8505 56297
rect 8557 56245 8629 56297
rect 8681 56245 9867 56297
rect 7817 56173 9867 56245
rect 7817 56121 7885 56173
rect 7937 56121 8009 56173
rect 8061 56121 8133 56173
rect 8185 56121 8257 56173
rect 8309 56121 8381 56173
rect 8433 56121 8505 56173
rect 8557 56121 8629 56173
rect 8681 56121 9867 56173
rect 7817 56049 9867 56121
rect 7817 55997 7885 56049
rect 7937 55997 8009 56049
rect 8061 55997 8133 56049
rect 8185 55997 8257 56049
rect 8309 55997 8381 56049
rect 8433 55997 8505 56049
rect 8557 55997 8629 56049
rect 8681 55997 9867 56049
rect 7817 55925 9867 55997
rect 7817 55873 7885 55925
rect 7937 55873 8009 55925
rect 8061 55873 8133 55925
rect 8185 55873 8257 55925
rect 8309 55873 8381 55925
rect 8433 55873 8505 55925
rect 8557 55873 8629 55925
rect 8681 55873 9867 55925
rect 7817 55801 9867 55873
rect 7817 55749 7885 55801
rect 7937 55749 8009 55801
rect 8061 55749 8133 55801
rect 8185 55749 8257 55801
rect 8309 55749 8381 55801
rect 8433 55749 8505 55801
rect 8557 55749 8629 55801
rect 8681 55749 9867 55801
rect 7817 55677 9867 55749
rect 7817 55625 7885 55677
rect 7937 55625 8009 55677
rect 8061 55625 8133 55677
rect 8185 55625 8257 55677
rect 8309 55625 8381 55677
rect 8433 55625 8505 55677
rect 8557 55625 8629 55677
rect 8681 55625 9867 55677
rect 7817 55553 9867 55625
rect 7817 55501 7885 55553
rect 7937 55501 8009 55553
rect 8061 55501 8133 55553
rect 8185 55501 8257 55553
rect 8309 55501 8381 55553
rect 8433 55501 8505 55553
rect 8557 55501 8629 55553
rect 8681 55501 9867 55553
rect 7817 55429 9867 55501
rect 7817 55377 7885 55429
rect 7937 55377 8009 55429
rect 8061 55377 8133 55429
rect 8185 55377 8257 55429
rect 8309 55377 8381 55429
rect 8433 55377 8505 55429
rect 8557 55377 8629 55429
rect 8681 55377 9867 55429
rect 7817 55305 9867 55377
rect 7817 55253 7885 55305
rect 7937 55253 8009 55305
rect 8061 55253 8133 55305
rect 8185 55253 8257 55305
rect 8309 55253 8381 55305
rect 8433 55253 8505 55305
rect 8557 55253 8629 55305
rect 8681 55253 9867 55305
rect 7817 55181 9867 55253
rect 7817 55129 7885 55181
rect 7937 55129 8009 55181
rect 8061 55129 8133 55181
rect 8185 55129 8257 55181
rect 8309 55129 8381 55181
rect 8433 55129 8505 55181
rect 8557 55129 8629 55181
rect 8681 55129 9867 55181
rect 7817 55057 9867 55129
rect 7817 55005 7885 55057
rect 7937 55005 8009 55057
rect 8061 55005 8133 55057
rect 8185 55005 8257 55057
rect 8309 55005 8381 55057
rect 8433 55005 8505 55057
rect 8557 55005 8629 55057
rect 8681 55005 9867 55057
rect 7817 54933 9867 55005
rect 7817 54881 7885 54933
rect 7937 54881 8009 54933
rect 8061 54881 8133 54933
rect 8185 54881 8257 54933
rect 8309 54881 8381 54933
rect 8433 54881 8505 54933
rect 8557 54881 8629 54933
rect 8681 54881 9867 54933
rect 7817 54809 9867 54881
rect 7817 54757 7885 54809
rect 7937 54757 8009 54809
rect 8061 54757 8133 54809
rect 8185 54757 8257 54809
rect 8309 54757 8381 54809
rect 8433 54757 8505 54809
rect 8557 54757 8629 54809
rect 8681 54757 9867 54809
rect 7817 54685 9867 54757
rect 7817 54633 7885 54685
rect 7937 54633 8009 54685
rect 8061 54633 8133 54685
rect 8185 54633 8257 54685
rect 8309 54633 8381 54685
rect 8433 54633 8505 54685
rect 8557 54633 8629 54685
rect 8681 54633 9867 54685
rect 7817 54561 9867 54633
rect 7817 54509 7885 54561
rect 7937 54509 8009 54561
rect 8061 54509 8133 54561
rect 8185 54509 8257 54561
rect 8309 54509 8381 54561
rect 8433 54509 8505 54561
rect 8557 54509 8629 54561
rect 8681 54509 9867 54561
rect 7817 54437 9867 54509
rect 7817 54385 7885 54437
rect 7937 54385 8009 54437
rect 8061 54385 8133 54437
rect 8185 54385 8257 54437
rect 8309 54385 8381 54437
rect 8433 54385 8505 54437
rect 8557 54385 8629 54437
rect 8681 54385 9867 54437
rect 7817 54313 9867 54385
rect 7817 54261 7885 54313
rect 7937 54261 8009 54313
rect 8061 54261 8133 54313
rect 8185 54261 8257 54313
rect 8309 54261 8381 54313
rect 8433 54261 8505 54313
rect 8557 54261 8629 54313
rect 8681 54261 9867 54313
rect 7817 54189 9867 54261
rect 7817 54137 7885 54189
rect 7937 54137 8009 54189
rect 8061 54137 8133 54189
rect 8185 54137 8257 54189
rect 8309 54137 8381 54189
rect 8433 54137 8505 54189
rect 8557 54137 8629 54189
rect 8681 54137 9867 54189
rect 7817 54065 9867 54137
rect 7817 54013 7885 54065
rect 7937 54013 8009 54065
rect 8061 54013 8133 54065
rect 8185 54013 8257 54065
rect 8309 54013 8381 54065
rect 8433 54013 8505 54065
rect 8557 54013 8629 54065
rect 8681 54013 9867 54065
rect 7817 53941 9867 54013
rect 7817 53889 7885 53941
rect 7937 53889 8009 53941
rect 8061 53889 8133 53941
rect 8185 53889 8257 53941
rect 8309 53889 8381 53941
rect 8433 53889 8505 53941
rect 8557 53889 8629 53941
rect 8681 53889 9867 53941
rect 7817 53817 9867 53889
rect 7817 53765 7885 53817
rect 7937 53765 8009 53817
rect 8061 53765 8133 53817
rect 8185 53765 8257 53817
rect 8309 53765 8381 53817
rect 8433 53765 8505 53817
rect 8557 53765 8629 53817
rect 8681 53765 9867 53817
rect 7817 53693 9867 53765
rect 7817 53641 7885 53693
rect 7937 53641 8009 53693
rect 8061 53641 8133 53693
rect 8185 53641 8257 53693
rect 8309 53641 8381 53693
rect 8433 53641 8505 53693
rect 8557 53641 8629 53693
rect 8681 53641 9867 53693
rect 7817 52588 9867 53641
rect 7817 52536 7886 52588
rect 7938 52536 8010 52588
rect 8062 52536 8134 52588
rect 8186 52536 8258 52588
rect 8310 52536 8382 52588
rect 8434 52536 8506 52588
rect 8558 52536 8630 52588
rect 8682 52536 8754 52588
rect 8806 52536 8878 52588
rect 8930 52536 9002 52588
rect 9054 52536 9126 52588
rect 9178 52536 9250 52588
rect 9302 52536 9374 52588
rect 9426 52536 9498 52588
rect 9550 52536 9622 52588
rect 9674 52536 9746 52588
rect 9798 52536 9867 52588
rect 7817 52464 9867 52536
rect 7817 52412 7886 52464
rect 7938 52412 8010 52464
rect 8062 52412 8134 52464
rect 8186 52412 8258 52464
rect 8310 52412 8382 52464
rect 8434 52412 8506 52464
rect 8558 52412 8630 52464
rect 8682 52412 8754 52464
rect 8806 52412 8878 52464
rect 8930 52412 9002 52464
rect 9054 52412 9126 52464
rect 9178 52412 9250 52464
rect 9302 52412 9374 52464
rect 9426 52412 9498 52464
rect 9550 52412 9622 52464
rect 9674 52412 9746 52464
rect 9798 52412 9867 52464
rect 7817 52340 9867 52412
rect 7817 52288 7886 52340
rect 7938 52288 8010 52340
rect 8062 52288 8134 52340
rect 8186 52288 8258 52340
rect 8310 52288 8382 52340
rect 8434 52288 8506 52340
rect 8558 52288 8630 52340
rect 8682 52288 8754 52340
rect 8806 52288 8878 52340
rect 8930 52288 9002 52340
rect 9054 52288 9126 52340
rect 9178 52288 9250 52340
rect 9302 52288 9374 52340
rect 9426 52288 9498 52340
rect 9550 52288 9622 52340
rect 9674 52288 9746 52340
rect 9798 52288 9867 52340
rect 7817 51627 9867 52288
rect 7817 51575 7886 51627
rect 7938 51575 8010 51627
rect 8062 51575 8134 51627
rect 8186 51575 8258 51627
rect 8310 51575 8382 51627
rect 8434 51575 8506 51627
rect 8558 51575 8630 51627
rect 8682 51575 8754 51627
rect 8806 51575 8878 51627
rect 8930 51575 9002 51627
rect 9054 51575 9126 51627
rect 9178 51575 9250 51627
rect 9302 51575 9374 51627
rect 9426 51575 9498 51627
rect 9550 51575 9622 51627
rect 9674 51575 9746 51627
rect 9798 51575 9867 51627
rect 7817 51503 9867 51575
rect 7817 51451 7886 51503
rect 7938 51451 8010 51503
rect 8062 51451 8134 51503
rect 8186 51451 8258 51503
rect 8310 51451 8382 51503
rect 8434 51451 8506 51503
rect 8558 51451 8630 51503
rect 8682 51451 8754 51503
rect 8806 51451 8878 51503
rect 8930 51451 9002 51503
rect 9054 51451 9126 51503
rect 9178 51451 9250 51503
rect 9302 51451 9374 51503
rect 9426 51451 9498 51503
rect 9550 51451 9622 51503
rect 9674 51451 9746 51503
rect 9798 51451 9867 51503
rect 7817 50948 9867 51451
rect 7817 50892 7884 50948
rect 7940 50892 8008 50948
rect 8064 50892 8132 50948
rect 8188 50892 8256 50948
rect 8312 50892 8380 50948
rect 8436 50892 8504 50948
rect 8560 50892 8628 50948
rect 8684 50892 8752 50948
rect 8808 50892 8876 50948
rect 8932 50892 9000 50948
rect 9056 50892 9124 50948
rect 9180 50892 9248 50948
rect 9304 50892 9372 50948
rect 9428 50892 9496 50948
rect 9552 50892 9620 50948
rect 9676 50892 9744 50948
rect 9800 50892 9867 50948
rect 7817 50824 9867 50892
rect 7817 50768 7884 50824
rect 7940 50768 8008 50824
rect 8064 50768 8132 50824
rect 8188 50768 8256 50824
rect 8312 50768 8380 50824
rect 8436 50768 8504 50824
rect 8560 50768 8628 50824
rect 8684 50768 8752 50824
rect 8808 50768 8876 50824
rect 8932 50768 9000 50824
rect 9056 50768 9124 50824
rect 9180 50768 9248 50824
rect 9304 50768 9372 50824
rect 9428 50768 9496 50824
rect 9552 50768 9620 50824
rect 9676 50768 9744 50824
rect 9800 50768 9867 50824
rect 7817 50700 9867 50768
rect 7817 50644 7884 50700
rect 7940 50644 8008 50700
rect 8064 50644 8132 50700
rect 8188 50644 8256 50700
rect 8312 50644 8380 50700
rect 8436 50644 8504 50700
rect 8560 50644 8628 50700
rect 8684 50644 8752 50700
rect 8808 50644 8876 50700
rect 8932 50644 9000 50700
rect 9056 50644 9124 50700
rect 9180 50644 9248 50700
rect 9304 50644 9372 50700
rect 9428 50644 9496 50700
rect 9552 50644 9620 50700
rect 9676 50644 9744 50700
rect 9800 50644 9867 50700
rect 7817 50641 7886 50644
rect 7938 50641 8010 50644
rect 8062 50641 8134 50644
rect 8186 50641 8258 50644
rect 8310 50641 8382 50644
rect 8434 50641 8506 50644
rect 8558 50641 8630 50644
rect 8682 50641 8754 50644
rect 8806 50641 8878 50644
rect 8930 50641 9002 50644
rect 9054 50641 9126 50644
rect 9178 50641 9250 50644
rect 9302 50641 9374 50644
rect 9426 50641 9498 50644
rect 9550 50641 9622 50644
rect 9674 50641 9746 50644
rect 9798 50641 9867 50644
rect 7817 50576 9867 50641
rect 7817 50520 7884 50576
rect 7940 50520 8008 50576
rect 8064 50520 8132 50576
rect 8188 50520 8256 50576
rect 8312 50520 8380 50576
rect 8436 50520 8504 50576
rect 8560 50520 8628 50576
rect 8684 50520 8752 50576
rect 8808 50520 8876 50576
rect 8932 50520 9000 50576
rect 9056 50520 9124 50576
rect 9180 50520 9248 50576
rect 9304 50520 9372 50576
rect 9428 50520 9496 50576
rect 9552 50520 9620 50576
rect 9676 50520 9744 50576
rect 9800 50520 9867 50576
rect 7817 50517 7886 50520
rect 7938 50517 8010 50520
rect 8062 50517 8134 50520
rect 8186 50517 8258 50520
rect 8310 50517 8382 50520
rect 8434 50517 8506 50520
rect 8558 50517 8630 50520
rect 8682 50517 8754 50520
rect 8806 50517 8878 50520
rect 8930 50517 9002 50520
rect 9054 50517 9126 50520
rect 9178 50517 9250 50520
rect 9302 50517 9374 50520
rect 9426 50517 9498 50520
rect 9550 50517 9622 50520
rect 9674 50517 9746 50520
rect 9798 50517 9867 50520
rect 7817 50452 9867 50517
rect 7817 50396 7884 50452
rect 7940 50396 8008 50452
rect 8064 50396 8132 50452
rect 8188 50396 8256 50452
rect 8312 50396 8380 50452
rect 8436 50396 8504 50452
rect 8560 50396 8628 50452
rect 8684 50396 8752 50452
rect 8808 50396 8876 50452
rect 8932 50396 9000 50452
rect 9056 50396 9124 50452
rect 9180 50396 9248 50452
rect 9304 50396 9372 50452
rect 9428 50396 9496 50452
rect 9552 50396 9620 50452
rect 9676 50396 9744 50452
rect 9800 50396 9867 50452
rect 7817 50328 9867 50396
rect 7817 50272 7884 50328
rect 7940 50272 8008 50328
rect 8064 50272 8132 50328
rect 8188 50272 8256 50328
rect 8312 50272 8380 50328
rect 8436 50272 8504 50328
rect 8560 50272 8628 50328
rect 8684 50272 8752 50328
rect 8808 50272 8876 50328
rect 8932 50272 9000 50328
rect 9056 50272 9124 50328
rect 9180 50272 9248 50328
rect 9304 50272 9372 50328
rect 9428 50272 9496 50328
rect 9552 50272 9620 50328
rect 9676 50272 9744 50328
rect 9800 50272 9867 50328
rect 7817 50204 9867 50272
rect 7817 50148 7884 50204
rect 7940 50148 8008 50204
rect 8064 50148 8132 50204
rect 8188 50148 8256 50204
rect 8312 50148 8380 50204
rect 8436 50148 8504 50204
rect 8560 50148 8628 50204
rect 8684 50148 8752 50204
rect 8808 50148 8876 50204
rect 8932 50148 9000 50204
rect 9056 50148 9124 50204
rect 9180 50148 9248 50204
rect 9304 50148 9372 50204
rect 9428 50148 9496 50204
rect 9552 50148 9620 50204
rect 9676 50148 9744 50204
rect 9800 50148 9867 50204
rect 7817 50080 9867 50148
rect 7817 50024 7884 50080
rect 7940 50024 8008 50080
rect 8064 50024 8132 50080
rect 8188 50024 8256 50080
rect 8312 50024 8380 50080
rect 8436 50024 8504 50080
rect 8560 50024 8628 50080
rect 8684 50024 8752 50080
rect 8808 50024 8876 50080
rect 8932 50024 9000 50080
rect 9056 50024 9124 50080
rect 9180 50024 9248 50080
rect 9304 50024 9372 50080
rect 9428 50024 9496 50080
rect 9552 50024 9620 50080
rect 9676 50024 9744 50080
rect 9800 50024 9867 50080
rect 7817 49956 9867 50024
rect 7817 49900 7884 49956
rect 7940 49900 8008 49956
rect 8064 49900 8132 49956
rect 8188 49900 8256 49956
rect 8312 49900 8380 49956
rect 8436 49900 8504 49956
rect 8560 49900 8628 49956
rect 8684 49900 8752 49956
rect 8808 49900 8876 49956
rect 8932 49900 9000 49956
rect 9056 49900 9124 49956
rect 9180 49900 9248 49956
rect 9304 49900 9372 49956
rect 9428 49900 9496 49956
rect 9552 49900 9620 49956
rect 9676 49900 9744 49956
rect 9800 49900 9867 49956
rect 7817 49832 9867 49900
rect 7817 49776 7884 49832
rect 7940 49776 8008 49832
rect 8064 49776 8132 49832
rect 8188 49776 8256 49832
rect 8312 49776 8380 49832
rect 8436 49776 8504 49832
rect 8560 49776 8628 49832
rect 8684 49776 8752 49832
rect 8808 49776 8876 49832
rect 8932 49776 9000 49832
rect 9056 49776 9124 49832
rect 9180 49776 9248 49832
rect 9304 49776 9372 49832
rect 9428 49776 9496 49832
rect 9552 49776 9620 49832
rect 9676 49776 9744 49832
rect 9800 49776 9867 49832
rect 7817 49759 9867 49776
rect 7817 49708 7886 49759
rect 7938 49708 8010 49759
rect 8062 49708 8134 49759
rect 8186 49708 8258 49759
rect 8310 49708 8382 49759
rect 8434 49708 8506 49759
rect 8558 49708 8630 49759
rect 8682 49708 8754 49759
rect 8806 49708 8878 49759
rect 8930 49708 9002 49759
rect 9054 49708 9126 49759
rect 9178 49708 9250 49759
rect 9302 49708 9374 49759
rect 9426 49708 9498 49759
rect 9550 49708 9622 49759
rect 9674 49708 9746 49759
rect 9798 49708 9867 49759
rect 7817 49652 7884 49708
rect 7940 49652 8008 49708
rect 8064 49652 8132 49708
rect 8188 49652 8256 49708
rect 8312 49652 8380 49708
rect 8436 49652 8504 49708
rect 8560 49652 8628 49708
rect 8684 49652 8752 49708
rect 8808 49652 8876 49708
rect 8932 49652 9000 49708
rect 9056 49652 9124 49708
rect 9180 49652 9248 49708
rect 9304 49652 9372 49708
rect 9428 49652 9496 49708
rect 9552 49652 9620 49708
rect 9676 49652 9744 49708
rect 9800 49652 9867 49708
rect 7817 49635 9867 49652
rect 7817 49583 7886 49635
rect 7938 49583 8010 49635
rect 8062 49583 8134 49635
rect 8186 49583 8258 49635
rect 8310 49583 8382 49635
rect 8434 49583 8506 49635
rect 8558 49583 8630 49635
rect 8682 49583 8754 49635
rect 8806 49583 8878 49635
rect 8930 49583 9002 49635
rect 9054 49583 9126 49635
rect 9178 49583 9250 49635
rect 9302 49583 9374 49635
rect 9426 49583 9498 49635
rect 9550 49583 9622 49635
rect 9674 49583 9746 49635
rect 9798 49583 9867 49635
rect 7817 48825 9867 49583
rect 7817 48773 7886 48825
rect 7938 48773 8010 48825
rect 8062 48773 8134 48825
rect 8186 48773 8258 48825
rect 8310 48773 8382 48825
rect 8434 48773 8506 48825
rect 8558 48773 8630 48825
rect 8682 48773 8754 48825
rect 8806 48773 8878 48825
rect 8930 48773 9002 48825
rect 9054 48773 9126 48825
rect 9178 48773 9250 48825
rect 9302 48773 9374 48825
rect 9426 48773 9498 48825
rect 9550 48773 9622 48825
rect 9674 48773 9746 48825
rect 9798 48773 9867 48825
rect 7817 48701 9867 48773
rect 7817 48649 7886 48701
rect 7938 48649 8010 48701
rect 8062 48649 8134 48701
rect 8186 48649 8258 48701
rect 8310 48649 8382 48701
rect 8434 48649 8506 48701
rect 8558 48649 8630 48701
rect 8682 48649 8754 48701
rect 8806 48649 8878 48701
rect 8930 48649 9002 48701
rect 9054 48649 9126 48701
rect 9178 48649 9250 48701
rect 9302 48649 9374 48701
rect 9426 48649 9498 48701
rect 9550 48649 9622 48701
rect 9674 48649 9746 48701
rect 9798 48649 9867 48701
rect 7817 47988 9867 48649
rect 7817 47936 7886 47988
rect 7938 47936 8010 47988
rect 8062 47936 8134 47988
rect 8186 47936 8258 47988
rect 8310 47936 8382 47988
rect 8434 47936 8506 47988
rect 8558 47936 8630 47988
rect 8682 47936 8754 47988
rect 8806 47936 8878 47988
rect 8930 47936 9002 47988
rect 9054 47936 9126 47988
rect 9178 47936 9250 47988
rect 9302 47936 9374 47988
rect 9426 47936 9498 47988
rect 9550 47936 9622 47988
rect 9674 47936 9746 47988
rect 9798 47936 9867 47988
rect 7817 47864 9867 47936
rect 7817 47812 7886 47864
rect 7938 47812 8010 47864
rect 8062 47812 8134 47864
rect 8186 47812 8258 47864
rect 8310 47812 8382 47864
rect 8434 47812 8506 47864
rect 8558 47812 8630 47864
rect 8682 47812 8754 47864
rect 8806 47812 8878 47864
rect 8930 47812 9002 47864
rect 9054 47812 9126 47864
rect 9178 47812 9250 47864
rect 9302 47812 9374 47864
rect 9426 47812 9498 47864
rect 9550 47812 9622 47864
rect 9674 47812 9746 47864
rect 9798 47812 9867 47864
rect 7817 47740 9867 47812
rect 7817 47688 7886 47740
rect 7938 47688 8010 47740
rect 8062 47688 8134 47740
rect 8186 47688 8258 47740
rect 8310 47688 8382 47740
rect 8434 47688 8506 47740
rect 8558 47688 8630 47740
rect 8682 47688 8754 47740
rect 8806 47688 8878 47740
rect 8930 47688 9002 47740
rect 9054 47688 9126 47740
rect 9178 47688 9250 47740
rect 9302 47688 9374 47740
rect 9426 47688 9498 47740
rect 9550 47688 9622 47740
rect 9674 47688 9746 47740
rect 9798 47688 9867 47740
rect 7817 46430 9867 47688
rect 9927 57108 10127 57278
rect 9927 57056 9947 57108
rect 9999 57056 10055 57108
rect 10107 57056 10127 57108
rect 9927 53484 10127 57056
rect 9927 53432 9947 53484
rect 9999 53432 10055 53484
rect 10107 53432 10127 53484
rect 9927 53376 10127 53432
rect 9927 53324 9947 53376
rect 9999 53324 10055 53376
rect 10107 53324 10127 53376
rect 9927 53268 10127 53324
rect 9927 53216 9947 53268
rect 9999 53216 10055 53268
rect 10107 53216 10127 53268
rect 9927 52548 10127 53216
rect 9927 52492 9937 52548
rect 9993 52492 10061 52548
rect 10117 52492 10127 52548
rect 9927 52424 10127 52492
rect 9927 52368 9937 52424
rect 9993 52368 10061 52424
rect 10117 52368 10127 52424
rect 9927 52300 10127 52368
rect 9927 52244 9937 52300
rect 9993 52244 10061 52300
rect 10117 52244 10127 52300
rect 9927 52176 10127 52244
rect 9927 52120 9937 52176
rect 9993 52120 10061 52176
rect 10117 52120 10127 52176
rect 9927 52052 10127 52120
rect 9927 51996 9937 52052
rect 9993 51996 10061 52052
rect 10117 51996 10127 52052
rect 9927 51965 9939 51996
rect 9991 51965 10063 51996
rect 10115 51965 10127 51996
rect 9927 51928 10127 51965
rect 9927 51872 9937 51928
rect 9993 51872 10061 51928
rect 10117 51872 10127 51928
rect 9927 51841 9939 51872
rect 9991 51841 10063 51872
rect 10115 51841 10127 51872
rect 9927 51804 10127 51841
rect 9927 51748 9937 51804
rect 9993 51748 10061 51804
rect 10117 51748 10127 51804
rect 9927 51680 10127 51748
rect 9927 51624 9937 51680
rect 9993 51624 10061 51680
rect 10117 51624 10127 51680
rect 9927 51556 10127 51624
rect 9927 51500 9937 51556
rect 9993 51500 10061 51556
rect 10117 51500 10127 51556
rect 9927 51432 10127 51500
rect 9927 51376 9937 51432
rect 9993 51376 10061 51432
rect 10117 51376 10127 51432
rect 9927 51308 10127 51376
rect 9927 51252 9937 51308
rect 9993 51252 10061 51308
rect 10117 51252 10127 51308
rect 9927 51222 10127 51252
rect 9927 51170 9939 51222
rect 9991 51170 10063 51222
rect 10115 51170 10127 51222
rect 9927 51098 10127 51170
rect 9927 51046 9939 51098
rect 9991 51046 10063 51098
rect 10115 51046 10127 51098
rect 9927 50974 10127 51046
rect 9927 50922 9939 50974
rect 9991 50922 10063 50974
rect 10115 50922 10127 50974
rect 9927 50288 10127 50922
rect 9927 50236 9939 50288
rect 9991 50236 10063 50288
rect 10115 50236 10127 50288
rect 9927 50164 10127 50236
rect 9927 50112 9939 50164
rect 9991 50112 10063 50164
rect 10115 50112 10127 50164
rect 9927 50040 10127 50112
rect 9927 49988 9939 50040
rect 9991 49988 10063 50040
rect 10115 49988 10127 50040
rect 9927 49354 10127 49988
rect 9927 49302 9939 49354
rect 9991 49302 10063 49354
rect 10115 49302 10127 49354
rect 9927 49230 10127 49302
rect 9927 49178 9939 49230
rect 9991 49178 10063 49230
rect 10115 49178 10127 49230
rect 9927 49106 10127 49178
rect 9927 49054 9939 49106
rect 9991 49054 10063 49106
rect 10115 49054 10127 49106
rect 9927 48435 10127 49054
rect 9927 48383 9939 48435
rect 9991 48383 10063 48435
rect 10115 48383 10127 48435
rect 9927 48311 10127 48383
rect 9927 48259 9939 48311
rect 9991 48259 10063 48311
rect 10115 48259 10127 48311
rect 9927 46430 10127 48259
rect 10187 56669 12237 57600
rect 10187 56617 10214 56669
rect 10266 56617 10338 56669
rect 10390 56617 10462 56669
rect 10514 56617 10586 56669
rect 10638 56617 11225 56669
rect 11277 56617 11349 56669
rect 11401 56617 11473 56669
rect 11525 56617 11597 56669
rect 11649 56617 11721 56669
rect 11773 56617 11845 56669
rect 11897 56617 11969 56669
rect 12021 56617 12093 56669
rect 12145 56617 12237 56669
rect 10187 56545 12237 56617
rect 10187 56493 10214 56545
rect 10266 56493 10338 56545
rect 10390 56493 10462 56545
rect 10514 56493 10586 56545
rect 10638 56493 11225 56545
rect 11277 56493 11349 56545
rect 11401 56493 11473 56545
rect 11525 56493 11597 56545
rect 11649 56493 11721 56545
rect 11773 56493 11845 56545
rect 11897 56493 11969 56545
rect 12021 56493 12093 56545
rect 12145 56493 12237 56545
rect 10187 56421 12237 56493
rect 10187 56369 10214 56421
rect 10266 56369 10338 56421
rect 10390 56369 10462 56421
rect 10514 56369 10586 56421
rect 10638 56369 11225 56421
rect 11277 56369 11349 56421
rect 11401 56369 11473 56421
rect 11525 56369 11597 56421
rect 11649 56369 11721 56421
rect 11773 56369 11845 56421
rect 11897 56369 11969 56421
rect 12021 56369 12093 56421
rect 12145 56369 12237 56421
rect 10187 56297 12237 56369
rect 10187 56245 10214 56297
rect 10266 56245 10338 56297
rect 10390 56245 10462 56297
rect 10514 56245 10586 56297
rect 10638 56245 11225 56297
rect 11277 56245 11349 56297
rect 11401 56245 11473 56297
rect 11525 56245 11597 56297
rect 11649 56245 11721 56297
rect 11773 56245 11845 56297
rect 11897 56245 11969 56297
rect 12021 56245 12093 56297
rect 12145 56245 12237 56297
rect 10187 56173 12237 56245
rect 10187 56121 10214 56173
rect 10266 56121 10338 56173
rect 10390 56121 10462 56173
rect 10514 56121 10586 56173
rect 10638 56121 11225 56173
rect 11277 56121 11349 56173
rect 11401 56121 11473 56173
rect 11525 56121 11597 56173
rect 11649 56121 11721 56173
rect 11773 56121 11845 56173
rect 11897 56121 11969 56173
rect 12021 56121 12093 56173
rect 12145 56121 12237 56173
rect 10187 56049 12237 56121
rect 10187 55997 10214 56049
rect 10266 55997 10338 56049
rect 10390 55997 10462 56049
rect 10514 55997 10586 56049
rect 10638 55997 11225 56049
rect 11277 55997 11349 56049
rect 11401 55997 11473 56049
rect 11525 55997 11597 56049
rect 11649 55997 11721 56049
rect 11773 55997 11845 56049
rect 11897 55997 11969 56049
rect 12021 55997 12093 56049
rect 12145 55997 12237 56049
rect 10187 55925 12237 55997
rect 10187 55873 10214 55925
rect 10266 55873 10338 55925
rect 10390 55873 10462 55925
rect 10514 55873 10586 55925
rect 10638 55873 11225 55925
rect 11277 55873 11349 55925
rect 11401 55873 11473 55925
rect 11525 55873 11597 55925
rect 11649 55873 11721 55925
rect 11773 55873 11845 55925
rect 11897 55873 11969 55925
rect 12021 55873 12093 55925
rect 12145 55873 12237 55925
rect 10187 55801 12237 55873
rect 10187 55749 10214 55801
rect 10266 55749 10338 55801
rect 10390 55749 10462 55801
rect 10514 55749 10586 55801
rect 10638 55749 11225 55801
rect 11277 55749 11349 55801
rect 11401 55749 11473 55801
rect 11525 55749 11597 55801
rect 11649 55749 11721 55801
rect 11773 55749 11845 55801
rect 11897 55749 11969 55801
rect 12021 55749 12093 55801
rect 12145 55749 12237 55801
rect 10187 55677 12237 55749
rect 10187 55625 10214 55677
rect 10266 55625 10338 55677
rect 10390 55625 10462 55677
rect 10514 55625 10586 55677
rect 10638 55625 11225 55677
rect 11277 55625 11349 55677
rect 11401 55625 11473 55677
rect 11525 55625 11597 55677
rect 11649 55625 11721 55677
rect 11773 55625 11845 55677
rect 11897 55625 11969 55677
rect 12021 55625 12093 55677
rect 12145 55625 12237 55677
rect 10187 55553 12237 55625
rect 10187 55501 10214 55553
rect 10266 55501 10338 55553
rect 10390 55501 10462 55553
rect 10514 55501 10586 55553
rect 10638 55501 11225 55553
rect 11277 55501 11349 55553
rect 11401 55501 11473 55553
rect 11525 55501 11597 55553
rect 11649 55501 11721 55553
rect 11773 55501 11845 55553
rect 11897 55501 11969 55553
rect 12021 55501 12093 55553
rect 12145 55501 12237 55553
rect 10187 55429 12237 55501
rect 10187 55377 10214 55429
rect 10266 55377 10338 55429
rect 10390 55377 10462 55429
rect 10514 55377 10586 55429
rect 10638 55377 11225 55429
rect 11277 55377 11349 55429
rect 11401 55377 11473 55429
rect 11525 55377 11597 55429
rect 11649 55377 11721 55429
rect 11773 55377 11845 55429
rect 11897 55377 11969 55429
rect 12021 55377 12093 55429
rect 12145 55377 12237 55429
rect 10187 55305 12237 55377
rect 10187 55253 10214 55305
rect 10266 55253 10338 55305
rect 10390 55253 10462 55305
rect 10514 55253 10586 55305
rect 10638 55253 11225 55305
rect 11277 55253 11349 55305
rect 11401 55253 11473 55305
rect 11525 55253 11597 55305
rect 11649 55253 11721 55305
rect 11773 55253 11845 55305
rect 11897 55253 11969 55305
rect 12021 55253 12093 55305
rect 12145 55253 12237 55305
rect 10187 55181 12237 55253
rect 10187 55129 10214 55181
rect 10266 55129 10338 55181
rect 10390 55129 10462 55181
rect 10514 55129 10586 55181
rect 10638 55129 11225 55181
rect 11277 55129 11349 55181
rect 11401 55129 11473 55181
rect 11525 55129 11597 55181
rect 11649 55129 11721 55181
rect 11773 55129 11845 55181
rect 11897 55129 11969 55181
rect 12021 55129 12093 55181
rect 12145 55129 12237 55181
rect 10187 55057 12237 55129
rect 10187 55005 10214 55057
rect 10266 55005 10338 55057
rect 10390 55005 10462 55057
rect 10514 55005 10586 55057
rect 10638 55005 11225 55057
rect 11277 55005 11349 55057
rect 11401 55005 11473 55057
rect 11525 55005 11597 55057
rect 11649 55005 11721 55057
rect 11773 55005 11845 55057
rect 11897 55005 11969 55057
rect 12021 55005 12093 55057
rect 12145 55005 12237 55057
rect 10187 54933 12237 55005
rect 10187 54881 10214 54933
rect 10266 54881 10338 54933
rect 10390 54881 10462 54933
rect 10514 54881 10586 54933
rect 10638 54881 11225 54933
rect 11277 54881 11349 54933
rect 11401 54881 11473 54933
rect 11525 54881 11597 54933
rect 11649 54881 11721 54933
rect 11773 54881 11845 54933
rect 11897 54881 11969 54933
rect 12021 54881 12093 54933
rect 12145 54881 12237 54933
rect 10187 54809 12237 54881
rect 10187 54757 10214 54809
rect 10266 54757 10338 54809
rect 10390 54757 10462 54809
rect 10514 54757 10586 54809
rect 10638 54757 11225 54809
rect 11277 54757 11349 54809
rect 11401 54757 11473 54809
rect 11525 54757 11597 54809
rect 11649 54757 11721 54809
rect 11773 54757 11845 54809
rect 11897 54757 11969 54809
rect 12021 54757 12093 54809
rect 12145 54757 12237 54809
rect 10187 54685 12237 54757
rect 10187 54633 10214 54685
rect 10266 54633 10338 54685
rect 10390 54633 10462 54685
rect 10514 54633 10586 54685
rect 10638 54633 11225 54685
rect 11277 54633 11349 54685
rect 11401 54633 11473 54685
rect 11525 54633 11597 54685
rect 11649 54633 11721 54685
rect 11773 54633 11845 54685
rect 11897 54633 11969 54685
rect 12021 54633 12093 54685
rect 12145 54633 12237 54685
rect 10187 54561 12237 54633
rect 10187 54509 10214 54561
rect 10266 54509 10338 54561
rect 10390 54509 10462 54561
rect 10514 54509 10586 54561
rect 10638 54509 11225 54561
rect 11277 54509 11349 54561
rect 11401 54509 11473 54561
rect 11525 54509 11597 54561
rect 11649 54509 11721 54561
rect 11773 54509 11845 54561
rect 11897 54509 11969 54561
rect 12021 54509 12093 54561
rect 12145 54509 12237 54561
rect 10187 54437 12237 54509
rect 10187 54385 10214 54437
rect 10266 54385 10338 54437
rect 10390 54385 10462 54437
rect 10514 54385 10586 54437
rect 10638 54385 11225 54437
rect 11277 54385 11349 54437
rect 11401 54385 11473 54437
rect 11525 54385 11597 54437
rect 11649 54385 11721 54437
rect 11773 54385 11845 54437
rect 11897 54385 11969 54437
rect 12021 54385 12093 54437
rect 12145 54385 12237 54437
rect 10187 54313 12237 54385
rect 10187 54261 10214 54313
rect 10266 54261 10338 54313
rect 10390 54261 10462 54313
rect 10514 54261 10586 54313
rect 10638 54261 11225 54313
rect 11277 54261 11349 54313
rect 11401 54261 11473 54313
rect 11525 54261 11597 54313
rect 11649 54261 11721 54313
rect 11773 54261 11845 54313
rect 11897 54261 11969 54313
rect 12021 54261 12093 54313
rect 12145 54261 12237 54313
rect 10187 54189 12237 54261
rect 10187 54137 10214 54189
rect 10266 54137 10338 54189
rect 10390 54137 10462 54189
rect 10514 54137 10586 54189
rect 10638 54137 11225 54189
rect 11277 54137 11349 54189
rect 11401 54137 11473 54189
rect 11525 54137 11597 54189
rect 11649 54137 11721 54189
rect 11773 54137 11845 54189
rect 11897 54137 11969 54189
rect 12021 54137 12093 54189
rect 12145 54137 12237 54189
rect 10187 54065 12237 54137
rect 10187 54013 10214 54065
rect 10266 54013 10338 54065
rect 10390 54013 10462 54065
rect 10514 54013 10586 54065
rect 10638 54013 11225 54065
rect 11277 54013 11349 54065
rect 11401 54013 11473 54065
rect 11525 54013 11597 54065
rect 11649 54013 11721 54065
rect 11773 54013 11845 54065
rect 11897 54013 11969 54065
rect 12021 54013 12093 54065
rect 12145 54013 12237 54065
rect 10187 53941 12237 54013
rect 10187 53889 10214 53941
rect 10266 53889 10338 53941
rect 10390 53889 10462 53941
rect 10514 53889 10586 53941
rect 10638 53889 11225 53941
rect 11277 53889 11349 53941
rect 11401 53889 11473 53941
rect 11525 53889 11597 53941
rect 11649 53889 11721 53941
rect 11773 53889 11845 53941
rect 11897 53889 11969 53941
rect 12021 53889 12093 53941
rect 12145 53889 12237 53941
rect 10187 53817 12237 53889
rect 10187 53765 10214 53817
rect 10266 53765 10338 53817
rect 10390 53765 10462 53817
rect 10514 53765 10586 53817
rect 10638 53765 11225 53817
rect 11277 53765 11349 53817
rect 11401 53765 11473 53817
rect 11525 53765 11597 53817
rect 11649 53765 11721 53817
rect 11773 53765 11845 53817
rect 11897 53765 11969 53817
rect 12021 53765 12093 53817
rect 12145 53765 12237 53817
rect 10187 53693 12237 53765
rect 10187 53641 10214 53693
rect 10266 53641 10338 53693
rect 10390 53641 10462 53693
rect 10514 53641 10586 53693
rect 10638 53641 11225 53693
rect 11277 53641 11349 53693
rect 11401 53641 11473 53693
rect 11525 53641 11597 53693
rect 11649 53641 11721 53693
rect 11773 53641 11845 53693
rect 11897 53641 11969 53693
rect 12021 53641 12093 53693
rect 12145 53641 12237 53693
rect 10187 52588 12237 53641
rect 10187 52536 10256 52588
rect 10308 52536 10380 52588
rect 10432 52536 10504 52588
rect 10556 52536 10628 52588
rect 10680 52536 10752 52588
rect 10804 52536 10876 52588
rect 10928 52536 11000 52588
rect 11052 52536 11124 52588
rect 11176 52536 11248 52588
rect 11300 52536 11372 52588
rect 11424 52536 11496 52588
rect 11548 52536 11620 52588
rect 11672 52536 11744 52588
rect 11796 52536 11868 52588
rect 11920 52536 11992 52588
rect 12044 52536 12116 52588
rect 12168 52536 12237 52588
rect 10187 52464 12237 52536
rect 10187 52412 10256 52464
rect 10308 52412 10380 52464
rect 10432 52412 10504 52464
rect 10556 52412 10628 52464
rect 10680 52412 10752 52464
rect 10804 52412 10876 52464
rect 10928 52412 11000 52464
rect 11052 52412 11124 52464
rect 11176 52412 11248 52464
rect 11300 52412 11372 52464
rect 11424 52412 11496 52464
rect 11548 52412 11620 52464
rect 11672 52412 11744 52464
rect 11796 52412 11868 52464
rect 11920 52412 11992 52464
rect 12044 52412 12116 52464
rect 12168 52412 12237 52464
rect 10187 52340 12237 52412
rect 10187 52288 10256 52340
rect 10308 52288 10380 52340
rect 10432 52288 10504 52340
rect 10556 52288 10628 52340
rect 10680 52288 10752 52340
rect 10804 52288 10876 52340
rect 10928 52288 11000 52340
rect 11052 52288 11124 52340
rect 11176 52288 11248 52340
rect 11300 52288 11372 52340
rect 11424 52288 11496 52340
rect 11548 52288 11620 52340
rect 11672 52288 11744 52340
rect 11796 52288 11868 52340
rect 11920 52288 11992 52340
rect 12044 52288 12116 52340
rect 12168 52288 12237 52340
rect 10187 51627 12237 52288
rect 10187 51575 10251 51627
rect 10303 51575 10375 51627
rect 10427 51575 10499 51627
rect 10551 51575 10623 51627
rect 10675 51575 10747 51627
rect 10799 51575 10871 51627
rect 10923 51575 10995 51627
rect 11047 51575 11119 51627
rect 11171 51575 11243 51627
rect 11295 51575 11367 51627
rect 11419 51575 12237 51627
rect 10187 51503 12237 51575
rect 10187 51451 10251 51503
rect 10303 51451 10375 51503
rect 10427 51451 10499 51503
rect 10551 51451 10623 51503
rect 10675 51451 10747 51503
rect 10799 51451 10871 51503
rect 10923 51451 10995 51503
rect 11047 51451 11119 51503
rect 11171 51451 11243 51503
rect 11295 51451 11367 51503
rect 11419 51451 12237 51503
rect 10187 50948 12237 51451
rect 10187 50892 10254 50948
rect 10310 50892 10378 50948
rect 10434 50892 10502 50948
rect 10558 50892 10626 50948
rect 10682 50892 10750 50948
rect 10806 50892 10874 50948
rect 10930 50892 10998 50948
rect 11054 50892 11122 50948
rect 11178 50892 11246 50948
rect 11302 50892 11370 50948
rect 11426 50892 11494 50948
rect 11550 50892 11618 50948
rect 11674 50892 11742 50948
rect 11798 50892 11866 50948
rect 11922 50892 11990 50948
rect 12046 50892 12114 50948
rect 12170 50892 12237 50948
rect 10187 50824 12237 50892
rect 10187 50768 10254 50824
rect 10310 50768 10378 50824
rect 10434 50768 10502 50824
rect 10558 50768 10626 50824
rect 10682 50768 10750 50824
rect 10806 50768 10874 50824
rect 10930 50768 10998 50824
rect 11054 50768 11122 50824
rect 11178 50768 11246 50824
rect 11302 50768 11370 50824
rect 11426 50768 11494 50824
rect 11550 50768 11618 50824
rect 11674 50768 11742 50824
rect 11798 50768 11866 50824
rect 11922 50768 11990 50824
rect 12046 50768 12114 50824
rect 12170 50768 12237 50824
rect 10187 50700 12237 50768
rect 10187 50693 10254 50700
rect 10310 50693 10378 50700
rect 10434 50693 10502 50700
rect 10558 50693 10626 50700
rect 10682 50693 10750 50700
rect 10806 50693 10874 50700
rect 10930 50693 10998 50700
rect 11054 50693 11122 50700
rect 11178 50693 11246 50700
rect 11302 50693 11370 50700
rect 10187 50641 10251 50693
rect 10310 50644 10375 50693
rect 10434 50644 10499 50693
rect 10558 50644 10623 50693
rect 10682 50644 10747 50693
rect 10806 50644 10871 50693
rect 10930 50644 10995 50693
rect 11054 50644 11119 50693
rect 11178 50644 11243 50693
rect 11302 50644 11367 50693
rect 11426 50644 11494 50700
rect 11550 50644 11618 50700
rect 11674 50644 11742 50700
rect 11798 50644 11866 50700
rect 11922 50644 11990 50700
rect 12046 50644 12114 50700
rect 12170 50644 12237 50700
rect 10303 50641 10375 50644
rect 10427 50641 10499 50644
rect 10551 50641 10623 50644
rect 10675 50641 10747 50644
rect 10799 50641 10871 50644
rect 10923 50641 10995 50644
rect 11047 50641 11119 50644
rect 11171 50641 11243 50644
rect 11295 50641 11367 50644
rect 11419 50641 12237 50644
rect 10187 50576 12237 50641
rect 10187 50569 10254 50576
rect 10310 50569 10378 50576
rect 10434 50569 10502 50576
rect 10558 50569 10626 50576
rect 10682 50569 10750 50576
rect 10806 50569 10874 50576
rect 10930 50569 10998 50576
rect 11054 50569 11122 50576
rect 11178 50569 11246 50576
rect 11302 50569 11370 50576
rect 10187 50517 10251 50569
rect 10310 50520 10375 50569
rect 10434 50520 10499 50569
rect 10558 50520 10623 50569
rect 10682 50520 10747 50569
rect 10806 50520 10871 50569
rect 10930 50520 10995 50569
rect 11054 50520 11119 50569
rect 11178 50520 11243 50569
rect 11302 50520 11367 50569
rect 11426 50520 11494 50576
rect 11550 50520 11618 50576
rect 11674 50520 11742 50576
rect 11798 50520 11866 50576
rect 11922 50520 11990 50576
rect 12046 50520 12114 50576
rect 12170 50520 12237 50576
rect 10303 50517 10375 50520
rect 10427 50517 10499 50520
rect 10551 50517 10623 50520
rect 10675 50517 10747 50520
rect 10799 50517 10871 50520
rect 10923 50517 10995 50520
rect 11047 50517 11119 50520
rect 11171 50517 11243 50520
rect 11295 50517 11367 50520
rect 11419 50517 12237 50520
rect 10187 50452 12237 50517
rect 10187 50396 10254 50452
rect 10310 50396 10378 50452
rect 10434 50396 10502 50452
rect 10558 50396 10626 50452
rect 10682 50396 10750 50452
rect 10806 50396 10874 50452
rect 10930 50396 10998 50452
rect 11054 50396 11122 50452
rect 11178 50396 11246 50452
rect 11302 50396 11370 50452
rect 11426 50396 11494 50452
rect 11550 50396 11618 50452
rect 11674 50396 11742 50452
rect 11798 50396 11866 50452
rect 11922 50396 11990 50452
rect 12046 50396 12114 50452
rect 12170 50396 12237 50452
rect 10187 50328 12237 50396
rect 10187 50272 10254 50328
rect 10310 50272 10378 50328
rect 10434 50272 10502 50328
rect 10558 50272 10626 50328
rect 10682 50272 10750 50328
rect 10806 50272 10874 50328
rect 10930 50272 10998 50328
rect 11054 50272 11122 50328
rect 11178 50272 11246 50328
rect 11302 50272 11370 50328
rect 11426 50272 11494 50328
rect 11550 50272 11618 50328
rect 11674 50272 11742 50328
rect 11798 50272 11866 50328
rect 11922 50272 11990 50328
rect 12046 50272 12114 50328
rect 12170 50272 12237 50328
rect 10187 50204 12237 50272
rect 10187 50148 10254 50204
rect 10310 50148 10378 50204
rect 10434 50148 10502 50204
rect 10558 50148 10626 50204
rect 10682 50148 10750 50204
rect 10806 50148 10874 50204
rect 10930 50148 10998 50204
rect 11054 50148 11122 50204
rect 11178 50148 11246 50204
rect 11302 50148 11370 50204
rect 11426 50148 11494 50204
rect 11550 50148 11618 50204
rect 11674 50148 11742 50204
rect 11798 50148 11866 50204
rect 11922 50148 11990 50204
rect 12046 50148 12114 50204
rect 12170 50148 12237 50204
rect 10187 50080 12237 50148
rect 10187 50024 10254 50080
rect 10310 50024 10378 50080
rect 10434 50024 10502 50080
rect 10558 50024 10626 50080
rect 10682 50024 10750 50080
rect 10806 50024 10874 50080
rect 10930 50024 10998 50080
rect 11054 50024 11122 50080
rect 11178 50024 11246 50080
rect 11302 50024 11370 50080
rect 11426 50024 11494 50080
rect 11550 50024 11618 50080
rect 11674 50024 11742 50080
rect 11798 50024 11866 50080
rect 11922 50024 11990 50080
rect 12046 50024 12114 50080
rect 12170 50024 12237 50080
rect 10187 49956 12237 50024
rect 10187 49900 10254 49956
rect 10310 49900 10378 49956
rect 10434 49900 10502 49956
rect 10558 49900 10626 49956
rect 10682 49900 10750 49956
rect 10806 49900 10874 49956
rect 10930 49900 10998 49956
rect 11054 49900 11122 49956
rect 11178 49900 11246 49956
rect 11302 49900 11370 49956
rect 11426 49900 11494 49956
rect 11550 49900 11618 49956
rect 11674 49900 11742 49956
rect 11798 49900 11866 49956
rect 11922 49900 11990 49956
rect 12046 49900 12114 49956
rect 12170 49900 12237 49956
rect 10187 49832 12237 49900
rect 10187 49776 10254 49832
rect 10310 49776 10378 49832
rect 10434 49776 10502 49832
rect 10558 49776 10626 49832
rect 10682 49776 10750 49832
rect 10806 49776 10874 49832
rect 10930 49776 10998 49832
rect 11054 49776 11122 49832
rect 11178 49776 11246 49832
rect 11302 49776 11370 49832
rect 11426 49776 11494 49832
rect 11550 49776 11618 49832
rect 11674 49776 11742 49832
rect 11798 49776 11866 49832
rect 11922 49776 11990 49832
rect 12046 49776 12114 49832
rect 12170 49776 12237 49832
rect 10187 49759 12237 49776
rect 10187 49707 10251 49759
rect 10303 49708 10375 49759
rect 10427 49708 10499 49759
rect 10551 49708 10623 49759
rect 10675 49708 10747 49759
rect 10799 49708 10871 49759
rect 10923 49708 10995 49759
rect 11047 49708 11119 49759
rect 11171 49708 11243 49759
rect 11295 49708 11367 49759
rect 11419 49708 12237 49759
rect 10310 49707 10375 49708
rect 10434 49707 10499 49708
rect 10558 49707 10623 49708
rect 10682 49707 10747 49708
rect 10806 49707 10871 49708
rect 10930 49707 10995 49708
rect 11054 49707 11119 49708
rect 11178 49707 11243 49708
rect 11302 49707 11367 49708
rect 10187 49652 10254 49707
rect 10310 49652 10378 49707
rect 10434 49652 10502 49707
rect 10558 49652 10626 49707
rect 10682 49652 10750 49707
rect 10806 49652 10874 49707
rect 10930 49652 10998 49707
rect 11054 49652 11122 49707
rect 11178 49652 11246 49707
rect 11302 49652 11370 49707
rect 11426 49652 11494 49708
rect 11550 49652 11618 49708
rect 11674 49652 11742 49708
rect 11798 49652 11866 49708
rect 11922 49652 11990 49708
rect 12046 49652 12114 49708
rect 12170 49652 12237 49708
rect 10187 49635 12237 49652
rect 10187 49583 10251 49635
rect 10303 49583 10375 49635
rect 10427 49583 10499 49635
rect 10551 49583 10623 49635
rect 10675 49583 10747 49635
rect 10799 49583 10871 49635
rect 10923 49583 10995 49635
rect 11047 49583 11119 49635
rect 11171 49583 11243 49635
rect 11295 49583 11367 49635
rect 11419 49583 12237 49635
rect 10187 48825 12237 49583
rect 10187 48773 10251 48825
rect 10303 48773 10375 48825
rect 10427 48773 10499 48825
rect 10551 48773 10623 48825
rect 10675 48773 10747 48825
rect 10799 48773 10871 48825
rect 10923 48773 10995 48825
rect 11047 48773 11119 48825
rect 11171 48773 11243 48825
rect 11295 48773 11367 48825
rect 11419 48773 12237 48825
rect 10187 48701 12237 48773
rect 10187 48649 10251 48701
rect 10303 48649 10375 48701
rect 10427 48649 10499 48701
rect 10551 48649 10623 48701
rect 10675 48649 10747 48701
rect 10799 48649 10871 48701
rect 10923 48649 10995 48701
rect 11047 48649 11119 48701
rect 11171 48649 11243 48701
rect 11295 48649 11367 48701
rect 11419 48649 12237 48701
rect 10187 47988 12237 48649
rect 10187 47936 10256 47988
rect 10308 47936 10380 47988
rect 10432 47936 10504 47988
rect 10556 47936 10628 47988
rect 10680 47936 10752 47988
rect 10804 47936 10876 47988
rect 10928 47936 11000 47988
rect 11052 47936 11124 47988
rect 11176 47936 11248 47988
rect 11300 47936 11372 47988
rect 11424 47936 11496 47988
rect 11548 47936 11620 47988
rect 11672 47936 11744 47988
rect 11796 47936 11868 47988
rect 11920 47936 11992 47988
rect 12044 47936 12116 47988
rect 12168 47936 12237 47988
rect 10187 47864 12237 47936
rect 10187 47812 10256 47864
rect 10308 47812 10380 47864
rect 10432 47812 10504 47864
rect 10556 47812 10628 47864
rect 10680 47812 10752 47864
rect 10804 47812 10876 47864
rect 10928 47812 11000 47864
rect 11052 47812 11124 47864
rect 11176 47812 11248 47864
rect 11300 47812 11372 47864
rect 11424 47812 11496 47864
rect 11548 47812 11620 47864
rect 11672 47812 11744 47864
rect 11796 47812 11868 47864
rect 11920 47812 11992 47864
rect 12044 47812 12116 47864
rect 12168 47812 12237 47864
rect 10187 47740 12237 47812
rect 10187 47688 10256 47740
rect 10308 47688 10380 47740
rect 10432 47688 10504 47740
rect 10556 47688 10628 47740
rect 10680 47688 10752 47740
rect 10804 47688 10876 47740
rect 10928 47688 11000 47740
rect 11052 47688 11124 47740
rect 11176 47688 11248 47740
rect 11300 47688 11372 47740
rect 11424 47688 11496 47740
rect 11548 47688 11620 47740
rect 11672 47688 11744 47740
rect 11796 47688 11868 47740
rect 11920 47688 11992 47740
rect 12044 47688 12116 47740
rect 12168 47688 12237 47740
rect 10187 46430 12237 47688
rect 12297 57108 12497 57278
rect 12297 57056 12317 57108
rect 12369 57056 12425 57108
rect 12477 57056 12497 57108
rect 12297 53484 12497 57056
rect 12297 53432 12317 53484
rect 12369 53432 12425 53484
rect 12477 53432 12497 53484
rect 12297 53376 12497 53432
rect 12297 53324 12317 53376
rect 12369 53324 12425 53376
rect 12477 53324 12497 53376
rect 12297 53268 12497 53324
rect 12297 53216 12317 53268
rect 12369 53216 12425 53268
rect 12477 53216 12497 53268
rect 12297 52548 12497 53216
rect 12297 52492 12307 52548
rect 12363 52492 12431 52548
rect 12487 52492 12497 52548
rect 12297 52424 12497 52492
rect 12297 52368 12307 52424
rect 12363 52368 12431 52424
rect 12487 52368 12497 52424
rect 12297 52300 12497 52368
rect 12297 52244 12307 52300
rect 12363 52244 12431 52300
rect 12487 52244 12497 52300
rect 12297 52176 12497 52244
rect 12297 52120 12307 52176
rect 12363 52120 12431 52176
rect 12487 52120 12497 52176
rect 12297 52052 12497 52120
rect 12297 51996 12307 52052
rect 12363 51996 12431 52052
rect 12487 51996 12497 52052
rect 12297 51928 12497 51996
rect 12297 51872 12307 51928
rect 12363 51872 12431 51928
rect 12487 51872 12497 51928
rect 12297 51804 12497 51872
rect 12297 51748 12307 51804
rect 12363 51748 12431 51804
rect 12487 51748 12497 51804
rect 12297 51680 12497 51748
rect 12297 51624 12307 51680
rect 12363 51624 12431 51680
rect 12487 51624 12497 51680
rect 12297 51556 12497 51624
rect 12297 51500 12307 51556
rect 12363 51500 12431 51556
rect 12487 51500 12497 51556
rect 12297 51432 12497 51500
rect 12297 51376 12307 51432
rect 12363 51376 12431 51432
rect 12487 51376 12497 51432
rect 12297 51308 12497 51376
rect 12297 51252 12307 51308
rect 12363 51252 12431 51308
rect 12487 51252 12497 51308
rect 12297 46430 12497 51252
rect 12817 56669 14717 57600
rect 12817 56617 13141 56669
rect 13193 56617 13265 56669
rect 13317 56617 13389 56669
rect 13441 56617 13513 56669
rect 13565 56617 13637 56669
rect 13689 56617 13761 56669
rect 13813 56617 13885 56669
rect 13937 56617 14009 56669
rect 14061 56617 14717 56669
rect 12817 56545 14717 56617
rect 12817 56493 13141 56545
rect 13193 56493 13265 56545
rect 13317 56493 13389 56545
rect 13441 56493 13513 56545
rect 13565 56493 13637 56545
rect 13689 56493 13761 56545
rect 13813 56493 13885 56545
rect 13937 56493 14009 56545
rect 14061 56493 14717 56545
rect 12817 56421 14717 56493
rect 12817 56369 13141 56421
rect 13193 56369 13265 56421
rect 13317 56369 13389 56421
rect 13441 56369 13513 56421
rect 13565 56369 13637 56421
rect 13689 56369 13761 56421
rect 13813 56369 13885 56421
rect 13937 56369 14009 56421
rect 14061 56369 14717 56421
rect 12817 56297 14717 56369
rect 12817 56245 13141 56297
rect 13193 56245 13265 56297
rect 13317 56245 13389 56297
rect 13441 56245 13513 56297
rect 13565 56245 13637 56297
rect 13689 56245 13761 56297
rect 13813 56245 13885 56297
rect 13937 56245 14009 56297
rect 14061 56245 14717 56297
rect 12817 56173 14717 56245
rect 12817 56121 13141 56173
rect 13193 56121 13265 56173
rect 13317 56121 13389 56173
rect 13441 56121 13513 56173
rect 13565 56121 13637 56173
rect 13689 56121 13761 56173
rect 13813 56121 13885 56173
rect 13937 56121 14009 56173
rect 14061 56121 14717 56173
rect 12817 56049 14717 56121
rect 12817 55997 13141 56049
rect 13193 55997 13265 56049
rect 13317 55997 13389 56049
rect 13441 55997 13513 56049
rect 13565 55997 13637 56049
rect 13689 55997 13761 56049
rect 13813 55997 13885 56049
rect 13937 55997 14009 56049
rect 14061 55997 14717 56049
rect 12817 55925 14717 55997
rect 12817 55873 13141 55925
rect 13193 55873 13265 55925
rect 13317 55873 13389 55925
rect 13441 55873 13513 55925
rect 13565 55873 13637 55925
rect 13689 55873 13761 55925
rect 13813 55873 13885 55925
rect 13937 55873 14009 55925
rect 14061 55873 14717 55925
rect 12817 55801 14717 55873
rect 12817 55749 13141 55801
rect 13193 55749 13265 55801
rect 13317 55749 13389 55801
rect 13441 55749 13513 55801
rect 13565 55749 13637 55801
rect 13689 55749 13761 55801
rect 13813 55749 13885 55801
rect 13937 55749 14009 55801
rect 14061 55749 14717 55801
rect 12817 55677 14717 55749
rect 12817 55625 13141 55677
rect 13193 55625 13265 55677
rect 13317 55625 13389 55677
rect 13441 55625 13513 55677
rect 13565 55625 13637 55677
rect 13689 55625 13761 55677
rect 13813 55625 13885 55677
rect 13937 55625 14009 55677
rect 14061 55625 14717 55677
rect 12817 55553 14717 55625
rect 12817 55501 13141 55553
rect 13193 55501 13265 55553
rect 13317 55501 13389 55553
rect 13441 55501 13513 55553
rect 13565 55501 13637 55553
rect 13689 55501 13761 55553
rect 13813 55501 13885 55553
rect 13937 55501 14009 55553
rect 14061 55501 14717 55553
rect 12817 55429 14717 55501
rect 12817 55377 13141 55429
rect 13193 55377 13265 55429
rect 13317 55377 13389 55429
rect 13441 55377 13513 55429
rect 13565 55377 13637 55429
rect 13689 55377 13761 55429
rect 13813 55377 13885 55429
rect 13937 55377 14009 55429
rect 14061 55377 14717 55429
rect 12817 55305 14717 55377
rect 12817 55253 13141 55305
rect 13193 55253 13265 55305
rect 13317 55253 13389 55305
rect 13441 55253 13513 55305
rect 13565 55253 13637 55305
rect 13689 55253 13761 55305
rect 13813 55253 13885 55305
rect 13937 55253 14009 55305
rect 14061 55253 14717 55305
rect 12817 55181 14717 55253
rect 12817 55129 13141 55181
rect 13193 55129 13265 55181
rect 13317 55129 13389 55181
rect 13441 55129 13513 55181
rect 13565 55129 13637 55181
rect 13689 55129 13761 55181
rect 13813 55129 13885 55181
rect 13937 55129 14009 55181
rect 14061 55129 14717 55181
rect 12817 55057 14717 55129
rect 12817 55005 13141 55057
rect 13193 55005 13265 55057
rect 13317 55005 13389 55057
rect 13441 55005 13513 55057
rect 13565 55005 13637 55057
rect 13689 55005 13761 55057
rect 13813 55005 13885 55057
rect 13937 55005 14009 55057
rect 14061 55005 14717 55057
rect 12817 54933 14717 55005
rect 12817 54881 13141 54933
rect 13193 54881 13265 54933
rect 13317 54881 13389 54933
rect 13441 54881 13513 54933
rect 13565 54881 13637 54933
rect 13689 54881 13761 54933
rect 13813 54881 13885 54933
rect 13937 54881 14009 54933
rect 14061 54881 14717 54933
rect 12817 54809 14717 54881
rect 12817 54757 13141 54809
rect 13193 54757 13265 54809
rect 13317 54757 13389 54809
rect 13441 54757 13513 54809
rect 13565 54757 13637 54809
rect 13689 54757 13761 54809
rect 13813 54757 13885 54809
rect 13937 54757 14009 54809
rect 14061 54757 14717 54809
rect 12817 54685 14717 54757
rect 12817 54633 13141 54685
rect 13193 54633 13265 54685
rect 13317 54633 13389 54685
rect 13441 54633 13513 54685
rect 13565 54633 13637 54685
rect 13689 54633 13761 54685
rect 13813 54633 13885 54685
rect 13937 54633 14009 54685
rect 14061 54633 14717 54685
rect 12817 54561 14717 54633
rect 12817 54509 13141 54561
rect 13193 54509 13265 54561
rect 13317 54509 13389 54561
rect 13441 54509 13513 54561
rect 13565 54509 13637 54561
rect 13689 54509 13761 54561
rect 13813 54509 13885 54561
rect 13937 54509 14009 54561
rect 14061 54509 14717 54561
rect 12817 54437 14717 54509
rect 12817 54385 13141 54437
rect 13193 54385 13265 54437
rect 13317 54385 13389 54437
rect 13441 54385 13513 54437
rect 13565 54385 13637 54437
rect 13689 54385 13761 54437
rect 13813 54385 13885 54437
rect 13937 54385 14009 54437
rect 14061 54385 14717 54437
rect 12817 54313 14717 54385
rect 12817 54261 13141 54313
rect 13193 54261 13265 54313
rect 13317 54261 13389 54313
rect 13441 54261 13513 54313
rect 13565 54261 13637 54313
rect 13689 54261 13761 54313
rect 13813 54261 13885 54313
rect 13937 54261 14009 54313
rect 14061 54261 14717 54313
rect 12817 54189 14717 54261
rect 12817 54137 13141 54189
rect 13193 54137 13265 54189
rect 13317 54137 13389 54189
rect 13441 54137 13513 54189
rect 13565 54137 13637 54189
rect 13689 54137 13761 54189
rect 13813 54137 13885 54189
rect 13937 54137 14009 54189
rect 14061 54137 14717 54189
rect 12817 54065 14717 54137
rect 12817 54013 13141 54065
rect 13193 54013 13265 54065
rect 13317 54013 13389 54065
rect 13441 54013 13513 54065
rect 13565 54013 13637 54065
rect 13689 54013 13761 54065
rect 13813 54013 13885 54065
rect 13937 54013 14009 54065
rect 14061 54013 14717 54065
rect 12817 53941 14717 54013
rect 12817 53889 13141 53941
rect 13193 53889 13265 53941
rect 13317 53889 13389 53941
rect 13441 53889 13513 53941
rect 13565 53889 13637 53941
rect 13689 53889 13761 53941
rect 13813 53889 13885 53941
rect 13937 53889 14009 53941
rect 14061 53889 14717 53941
rect 12817 53817 14717 53889
rect 12817 53765 13141 53817
rect 13193 53765 13265 53817
rect 13317 53765 13389 53817
rect 13441 53765 13513 53817
rect 13565 53765 13637 53817
rect 13689 53765 13761 53817
rect 13813 53765 13885 53817
rect 13937 53765 14009 53817
rect 14061 53765 14717 53817
rect 12817 53693 14717 53765
rect 12817 53641 13141 53693
rect 13193 53641 13265 53693
rect 13317 53641 13389 53693
rect 13441 53641 13513 53693
rect 13565 53641 13637 53693
rect 13689 53641 13761 53693
rect 13813 53641 13885 53693
rect 13937 53641 14009 53693
rect 14061 53641 14717 53693
rect 12817 50948 14717 53641
rect 14892 52576 14989 52600
rect 14892 51224 14902 52576
rect 14958 51224 14989 52576
rect 14892 51200 14989 51224
rect 12817 50892 12871 50948
rect 12927 50892 12995 50948
rect 13051 50892 13119 50948
rect 13175 50892 13243 50948
rect 13299 50892 13367 50948
rect 13423 50892 13491 50948
rect 13547 50892 13615 50948
rect 13671 50892 13739 50948
rect 13795 50892 13863 50948
rect 13919 50892 13987 50948
rect 14043 50892 14111 50948
rect 14167 50892 14235 50948
rect 14291 50892 14359 50948
rect 14415 50892 14483 50948
rect 14539 50892 14607 50948
rect 14663 50892 14717 50948
rect 12817 50824 14717 50892
rect 12817 50768 12871 50824
rect 12927 50768 12995 50824
rect 13051 50768 13119 50824
rect 13175 50768 13243 50824
rect 13299 50768 13367 50824
rect 13423 50768 13491 50824
rect 13547 50768 13615 50824
rect 13671 50768 13739 50824
rect 13795 50768 13863 50824
rect 13919 50768 13987 50824
rect 14043 50768 14111 50824
rect 14167 50768 14235 50824
rect 14291 50768 14359 50824
rect 14415 50768 14483 50824
rect 14539 50768 14607 50824
rect 14663 50768 14717 50824
rect 12817 50700 14717 50768
rect 12817 50644 12871 50700
rect 12927 50644 12995 50700
rect 13051 50644 13119 50700
rect 13175 50644 13243 50700
rect 13299 50644 13367 50700
rect 13423 50644 13491 50700
rect 13547 50644 13615 50700
rect 13671 50644 13739 50700
rect 13795 50644 13863 50700
rect 13919 50644 13987 50700
rect 14043 50644 14111 50700
rect 14167 50644 14235 50700
rect 14291 50644 14359 50700
rect 14415 50644 14483 50700
rect 14539 50644 14607 50700
rect 14663 50644 14717 50700
rect 12817 50576 14717 50644
rect 12817 50520 12871 50576
rect 12927 50520 12995 50576
rect 13051 50520 13119 50576
rect 13175 50520 13243 50576
rect 13299 50520 13367 50576
rect 13423 50520 13491 50576
rect 13547 50520 13615 50576
rect 13671 50520 13739 50576
rect 13795 50520 13863 50576
rect 13919 50520 13987 50576
rect 14043 50520 14111 50576
rect 14167 50520 14235 50576
rect 14291 50520 14359 50576
rect 14415 50520 14483 50576
rect 14539 50520 14607 50576
rect 14663 50520 14717 50576
rect 12817 50452 14717 50520
rect 12817 50396 12871 50452
rect 12927 50396 12995 50452
rect 13051 50396 13119 50452
rect 13175 50396 13243 50452
rect 13299 50396 13367 50452
rect 13423 50396 13491 50452
rect 13547 50396 13615 50452
rect 13671 50396 13739 50452
rect 13795 50396 13863 50452
rect 13919 50396 13987 50452
rect 14043 50396 14111 50452
rect 14167 50396 14235 50452
rect 14291 50396 14359 50452
rect 14415 50396 14483 50452
rect 14539 50396 14607 50452
rect 14663 50396 14717 50452
rect 12817 50328 14717 50396
rect 12817 50272 12871 50328
rect 12927 50272 12995 50328
rect 13051 50272 13119 50328
rect 13175 50272 13243 50328
rect 13299 50272 13367 50328
rect 13423 50272 13491 50328
rect 13547 50272 13615 50328
rect 13671 50272 13739 50328
rect 13795 50272 13863 50328
rect 13919 50272 13987 50328
rect 14043 50272 14111 50328
rect 14167 50272 14235 50328
rect 14291 50272 14359 50328
rect 14415 50272 14483 50328
rect 14539 50272 14607 50328
rect 14663 50272 14717 50328
rect 12817 50204 14717 50272
rect 12817 50148 12871 50204
rect 12927 50148 12995 50204
rect 13051 50148 13119 50204
rect 13175 50148 13243 50204
rect 13299 50148 13367 50204
rect 13423 50148 13491 50204
rect 13547 50148 13615 50204
rect 13671 50148 13739 50204
rect 13795 50148 13863 50204
rect 13919 50148 13987 50204
rect 14043 50148 14111 50204
rect 14167 50148 14235 50204
rect 14291 50148 14359 50204
rect 14415 50148 14483 50204
rect 14539 50148 14607 50204
rect 14663 50148 14717 50204
rect 12817 50080 14717 50148
rect 12817 50024 12871 50080
rect 12927 50024 12995 50080
rect 13051 50024 13119 50080
rect 13175 50024 13243 50080
rect 13299 50024 13367 50080
rect 13423 50024 13491 50080
rect 13547 50024 13615 50080
rect 13671 50024 13739 50080
rect 13795 50024 13863 50080
rect 13919 50024 13987 50080
rect 14043 50024 14111 50080
rect 14167 50024 14235 50080
rect 14291 50024 14359 50080
rect 14415 50024 14483 50080
rect 14539 50024 14607 50080
rect 14663 50024 14717 50080
rect 12817 49956 14717 50024
rect 12817 49900 12871 49956
rect 12927 49900 12995 49956
rect 13051 49900 13119 49956
rect 13175 49900 13243 49956
rect 13299 49900 13367 49956
rect 13423 49900 13491 49956
rect 13547 49900 13615 49956
rect 13671 49900 13739 49956
rect 13795 49900 13863 49956
rect 13919 49900 13987 49956
rect 14043 49900 14111 49956
rect 14167 49900 14235 49956
rect 14291 49900 14359 49956
rect 14415 49900 14483 49956
rect 14539 49900 14607 49956
rect 14663 49900 14717 49956
rect 12817 49832 14717 49900
rect 12817 49776 12871 49832
rect 12927 49776 12995 49832
rect 13051 49776 13119 49832
rect 13175 49776 13243 49832
rect 13299 49776 13367 49832
rect 13423 49776 13491 49832
rect 13547 49776 13615 49832
rect 13671 49776 13739 49832
rect 13795 49776 13863 49832
rect 13919 49776 13987 49832
rect 14043 49776 14111 49832
rect 14167 49776 14235 49832
rect 14291 49776 14359 49832
rect 14415 49776 14483 49832
rect 14539 49776 14607 49832
rect 14663 49776 14717 49832
rect 12817 49708 14717 49776
rect 12817 49652 12871 49708
rect 12927 49652 12995 49708
rect 13051 49652 13119 49708
rect 13175 49652 13243 49708
rect 13299 49652 13367 49708
rect 13423 49652 13491 49708
rect 13547 49652 13615 49708
rect 13671 49652 13739 49708
rect 13795 49652 13863 49708
rect 13919 49652 13987 49708
rect 14043 49652 14111 49708
rect 14167 49652 14235 49708
rect 14291 49652 14359 49708
rect 14415 49652 14483 49708
rect 14539 49652 14607 49708
rect 14663 49652 14717 49708
rect 12817 46430 14717 49652
rect 2481 44842 2681 46158
rect 4851 44842 5051 46158
rect 7265 44842 7713 46158
rect 9927 44842 10127 46158
rect 12297 44842 12497 46158
rect 2798 43242 4734 44558
rect 5168 43242 7104 44558
rect 7874 43242 9810 44558
rect 10244 43242 12180 44558
rect 12861 43242 14673 44558
rect 2798 41642 4734 42958
rect 5168 41642 7104 42958
rect 7874 41642 9810 42958
rect 10244 41642 12180 42958
rect 12861 41642 14673 42958
rect 2481 40050 2681 41360
rect 2741 40050 4791 41360
rect 4851 40050 5051 41360
rect 5111 40050 7161 41360
rect 7221 40050 7757 41360
rect 7817 40050 9867 41360
rect 9927 40050 10127 41360
rect 10187 40050 12237 41360
rect 12297 40050 12497 41360
rect 12817 41358 14669 41360
rect 12817 40050 14673 41358
rect 2798 40042 4734 40050
rect 5168 40042 7104 40050
rect 7874 40042 9810 40050
rect 10244 40042 12180 40050
rect 12861 40042 14673 40050
rect 2798 39748 4734 39758
rect 2798 39692 2808 39748
rect 2864 39692 2932 39748
rect 2988 39692 3056 39748
rect 3112 39692 3180 39748
rect 3236 39692 3304 39748
rect 3360 39692 3428 39748
rect 3484 39692 3552 39748
rect 3608 39692 3676 39748
rect 3732 39692 3800 39748
rect 3856 39692 3924 39748
rect 3980 39692 4048 39748
rect 4104 39692 4172 39748
rect 4228 39692 4296 39748
rect 4352 39692 4420 39748
rect 4476 39692 4544 39748
rect 4600 39692 4668 39748
rect 4724 39692 4734 39748
rect 2798 39624 4734 39692
rect 2798 39568 2808 39624
rect 2864 39568 2932 39624
rect 2988 39568 3056 39624
rect 3112 39568 3180 39624
rect 3236 39568 3304 39624
rect 3360 39568 3428 39624
rect 3484 39568 3552 39624
rect 3608 39568 3676 39624
rect 3732 39568 3800 39624
rect 3856 39568 3924 39624
rect 3980 39568 4048 39624
rect 4104 39568 4172 39624
rect 4228 39568 4296 39624
rect 4352 39568 4420 39624
rect 4476 39568 4544 39624
rect 4600 39568 4668 39624
rect 4724 39568 4734 39624
rect 2798 39500 4734 39568
rect 2798 39444 2808 39500
rect 2864 39444 2932 39500
rect 2988 39444 3056 39500
rect 3112 39444 3180 39500
rect 3236 39444 3304 39500
rect 3360 39444 3428 39500
rect 3484 39444 3552 39500
rect 3608 39444 3676 39500
rect 3732 39444 3800 39500
rect 3856 39444 3924 39500
rect 3980 39444 4048 39500
rect 4104 39444 4172 39500
rect 4228 39444 4296 39500
rect 4352 39444 4420 39500
rect 4476 39444 4544 39500
rect 4600 39444 4668 39500
rect 4724 39444 4734 39500
rect 2798 39376 4734 39444
rect 2798 39320 2808 39376
rect 2864 39320 2932 39376
rect 2988 39320 3056 39376
rect 3112 39320 3180 39376
rect 3236 39320 3304 39376
rect 3360 39320 3428 39376
rect 3484 39320 3552 39376
rect 3608 39320 3676 39376
rect 3732 39320 3800 39376
rect 3856 39320 3924 39376
rect 3980 39320 4048 39376
rect 4104 39320 4172 39376
rect 4228 39320 4296 39376
rect 4352 39320 4420 39376
rect 4476 39320 4544 39376
rect 4600 39320 4668 39376
rect 4724 39320 4734 39376
rect 2798 39252 4734 39320
rect 2798 39196 2808 39252
rect 2864 39196 2932 39252
rect 2988 39196 3056 39252
rect 3112 39196 3180 39252
rect 3236 39196 3304 39252
rect 3360 39196 3428 39252
rect 3484 39196 3552 39252
rect 3608 39196 3676 39252
rect 3732 39196 3800 39252
rect 3856 39196 3924 39252
rect 3980 39196 4048 39252
rect 4104 39196 4172 39252
rect 4228 39196 4296 39252
rect 4352 39196 4420 39252
rect 4476 39196 4544 39252
rect 4600 39196 4668 39252
rect 4724 39196 4734 39252
rect 2798 39128 4734 39196
rect 2798 39072 2808 39128
rect 2864 39072 2932 39128
rect 2988 39072 3056 39128
rect 3112 39072 3180 39128
rect 3236 39072 3304 39128
rect 3360 39072 3428 39128
rect 3484 39072 3552 39128
rect 3608 39072 3676 39128
rect 3732 39072 3800 39128
rect 3856 39072 3924 39128
rect 3980 39072 4048 39128
rect 4104 39072 4172 39128
rect 4228 39072 4296 39128
rect 4352 39072 4420 39128
rect 4476 39072 4544 39128
rect 4600 39072 4668 39128
rect 4724 39072 4734 39128
rect 2798 39004 4734 39072
rect 2798 38948 2808 39004
rect 2864 38948 2932 39004
rect 2988 38948 3056 39004
rect 3112 38948 3180 39004
rect 3236 38948 3304 39004
rect 3360 38948 3428 39004
rect 3484 38948 3552 39004
rect 3608 38948 3676 39004
rect 3732 38948 3800 39004
rect 3856 38948 3924 39004
rect 3980 38948 4048 39004
rect 4104 38948 4172 39004
rect 4228 38948 4296 39004
rect 4352 38948 4420 39004
rect 4476 38948 4544 39004
rect 4600 38948 4668 39004
rect 4724 38948 4734 39004
rect 2798 38880 4734 38948
rect 2798 38824 2808 38880
rect 2864 38824 2932 38880
rect 2988 38824 3056 38880
rect 3112 38824 3180 38880
rect 3236 38824 3304 38880
rect 3360 38824 3428 38880
rect 3484 38824 3552 38880
rect 3608 38824 3676 38880
rect 3732 38824 3800 38880
rect 3856 38824 3924 38880
rect 3980 38824 4048 38880
rect 4104 38824 4172 38880
rect 4228 38824 4296 38880
rect 4352 38824 4420 38880
rect 4476 38824 4544 38880
rect 4600 38824 4668 38880
rect 4724 38824 4734 38880
rect 2798 38756 4734 38824
rect 2798 38700 2808 38756
rect 2864 38700 2932 38756
rect 2988 38700 3056 38756
rect 3112 38700 3180 38756
rect 3236 38700 3304 38756
rect 3360 38700 3428 38756
rect 3484 38700 3552 38756
rect 3608 38700 3676 38756
rect 3732 38700 3800 38756
rect 3856 38700 3924 38756
rect 3980 38700 4048 38756
rect 4104 38700 4172 38756
rect 4228 38700 4296 38756
rect 4352 38700 4420 38756
rect 4476 38700 4544 38756
rect 4600 38700 4668 38756
rect 4724 38700 4734 38756
rect 2798 38632 4734 38700
rect 2798 38576 2808 38632
rect 2864 38576 2932 38632
rect 2988 38576 3056 38632
rect 3112 38576 3180 38632
rect 3236 38576 3304 38632
rect 3360 38576 3428 38632
rect 3484 38576 3552 38632
rect 3608 38576 3676 38632
rect 3732 38576 3800 38632
rect 3856 38576 3924 38632
rect 3980 38576 4048 38632
rect 4104 38576 4172 38632
rect 4228 38576 4296 38632
rect 4352 38576 4420 38632
rect 4476 38576 4544 38632
rect 4600 38576 4668 38632
rect 4724 38576 4734 38632
rect 2798 38508 4734 38576
rect 2798 38452 2808 38508
rect 2864 38452 2932 38508
rect 2988 38452 3056 38508
rect 3112 38452 3180 38508
rect 3236 38452 3304 38508
rect 3360 38452 3428 38508
rect 3484 38452 3552 38508
rect 3608 38452 3676 38508
rect 3732 38452 3800 38508
rect 3856 38452 3924 38508
rect 3980 38452 4048 38508
rect 4104 38452 4172 38508
rect 4228 38452 4296 38508
rect 4352 38452 4420 38508
rect 4476 38452 4544 38508
rect 4600 38452 4668 38508
rect 4724 38452 4734 38508
rect 2798 38442 4734 38452
rect 5168 39748 7104 39758
rect 5168 39692 5178 39748
rect 5234 39692 5302 39748
rect 5358 39692 5426 39748
rect 5482 39692 5550 39748
rect 5606 39692 5674 39748
rect 5730 39692 5798 39748
rect 5854 39692 5922 39748
rect 5978 39692 6046 39748
rect 6102 39692 6170 39748
rect 6226 39692 6294 39748
rect 6350 39692 6418 39748
rect 6474 39692 6542 39748
rect 6598 39692 6666 39748
rect 6722 39692 6790 39748
rect 6846 39692 6914 39748
rect 6970 39692 7038 39748
rect 7094 39692 7104 39748
rect 5168 39624 7104 39692
rect 5168 39568 5178 39624
rect 5234 39568 5302 39624
rect 5358 39568 5426 39624
rect 5482 39568 5550 39624
rect 5606 39568 5674 39624
rect 5730 39568 5798 39624
rect 5854 39568 5922 39624
rect 5978 39568 6046 39624
rect 6102 39568 6170 39624
rect 6226 39568 6294 39624
rect 6350 39568 6418 39624
rect 6474 39568 6542 39624
rect 6598 39568 6666 39624
rect 6722 39568 6790 39624
rect 6846 39568 6914 39624
rect 6970 39568 7038 39624
rect 7094 39568 7104 39624
rect 5168 39500 7104 39568
rect 5168 39444 5178 39500
rect 5234 39444 5302 39500
rect 5358 39444 5426 39500
rect 5482 39444 5550 39500
rect 5606 39444 5674 39500
rect 5730 39444 5798 39500
rect 5854 39444 5922 39500
rect 5978 39444 6046 39500
rect 6102 39444 6170 39500
rect 6226 39444 6294 39500
rect 6350 39444 6418 39500
rect 6474 39444 6542 39500
rect 6598 39444 6666 39500
rect 6722 39444 6790 39500
rect 6846 39444 6914 39500
rect 6970 39444 7038 39500
rect 7094 39444 7104 39500
rect 5168 39376 7104 39444
rect 5168 39320 5178 39376
rect 5234 39320 5302 39376
rect 5358 39320 5426 39376
rect 5482 39320 5550 39376
rect 5606 39320 5674 39376
rect 5730 39320 5798 39376
rect 5854 39320 5922 39376
rect 5978 39320 6046 39376
rect 6102 39320 6170 39376
rect 6226 39320 6294 39376
rect 6350 39320 6418 39376
rect 6474 39320 6542 39376
rect 6598 39320 6666 39376
rect 6722 39320 6790 39376
rect 6846 39320 6914 39376
rect 6970 39320 7038 39376
rect 7094 39320 7104 39376
rect 5168 39252 7104 39320
rect 5168 39196 5178 39252
rect 5234 39196 5302 39252
rect 5358 39196 5426 39252
rect 5482 39196 5550 39252
rect 5606 39196 5674 39252
rect 5730 39196 5798 39252
rect 5854 39196 5922 39252
rect 5978 39196 6046 39252
rect 6102 39196 6170 39252
rect 6226 39196 6294 39252
rect 6350 39196 6418 39252
rect 6474 39196 6542 39252
rect 6598 39196 6666 39252
rect 6722 39196 6790 39252
rect 6846 39196 6914 39252
rect 6970 39196 7038 39252
rect 7094 39196 7104 39252
rect 5168 39128 7104 39196
rect 5168 39072 5178 39128
rect 5234 39072 5302 39128
rect 5358 39072 5426 39128
rect 5482 39072 5550 39128
rect 5606 39072 5674 39128
rect 5730 39072 5798 39128
rect 5854 39072 5922 39128
rect 5978 39072 6046 39128
rect 6102 39072 6170 39128
rect 6226 39072 6294 39128
rect 6350 39072 6418 39128
rect 6474 39072 6542 39128
rect 6598 39072 6666 39128
rect 6722 39072 6790 39128
rect 6846 39072 6914 39128
rect 6970 39072 7038 39128
rect 7094 39072 7104 39128
rect 5168 39004 7104 39072
rect 5168 38948 5178 39004
rect 5234 38948 5302 39004
rect 5358 38948 5426 39004
rect 5482 38948 5550 39004
rect 5606 38948 5674 39004
rect 5730 38948 5798 39004
rect 5854 38948 5922 39004
rect 5978 38948 6046 39004
rect 6102 38948 6170 39004
rect 6226 38948 6294 39004
rect 6350 38948 6418 39004
rect 6474 38948 6542 39004
rect 6598 38948 6666 39004
rect 6722 38948 6790 39004
rect 6846 38948 6914 39004
rect 6970 38948 7038 39004
rect 7094 38948 7104 39004
rect 5168 38880 7104 38948
rect 5168 38824 5178 38880
rect 5234 38824 5302 38880
rect 5358 38824 5426 38880
rect 5482 38824 5550 38880
rect 5606 38824 5674 38880
rect 5730 38824 5798 38880
rect 5854 38824 5922 38880
rect 5978 38824 6046 38880
rect 6102 38824 6170 38880
rect 6226 38824 6294 38880
rect 6350 38824 6418 38880
rect 6474 38824 6542 38880
rect 6598 38824 6666 38880
rect 6722 38824 6790 38880
rect 6846 38824 6914 38880
rect 6970 38824 7038 38880
rect 7094 38824 7104 38880
rect 5168 38756 7104 38824
rect 5168 38700 5178 38756
rect 5234 38700 5302 38756
rect 5358 38700 5426 38756
rect 5482 38700 5550 38756
rect 5606 38700 5674 38756
rect 5730 38700 5798 38756
rect 5854 38700 5922 38756
rect 5978 38700 6046 38756
rect 6102 38700 6170 38756
rect 6226 38700 6294 38756
rect 6350 38700 6418 38756
rect 6474 38700 6542 38756
rect 6598 38700 6666 38756
rect 6722 38700 6790 38756
rect 6846 38700 6914 38756
rect 6970 38700 7038 38756
rect 7094 38700 7104 38756
rect 5168 38632 7104 38700
rect 5168 38576 5178 38632
rect 5234 38576 5302 38632
rect 5358 38576 5426 38632
rect 5482 38576 5550 38632
rect 5606 38576 5674 38632
rect 5730 38576 5798 38632
rect 5854 38576 5922 38632
rect 5978 38576 6046 38632
rect 6102 38576 6170 38632
rect 6226 38576 6294 38632
rect 6350 38576 6418 38632
rect 6474 38576 6542 38632
rect 6598 38576 6666 38632
rect 6722 38576 6790 38632
rect 6846 38576 6914 38632
rect 6970 38576 7038 38632
rect 7094 38576 7104 38632
rect 5168 38508 7104 38576
rect 5168 38452 5178 38508
rect 5234 38452 5302 38508
rect 5358 38452 5426 38508
rect 5482 38452 5550 38508
rect 5606 38452 5674 38508
rect 5730 38452 5798 38508
rect 5854 38452 5922 38508
rect 5978 38452 6046 38508
rect 6102 38452 6170 38508
rect 6226 38452 6294 38508
rect 6350 38452 6418 38508
rect 6474 38452 6542 38508
rect 6598 38452 6666 38508
rect 6722 38452 6790 38508
rect 6846 38452 6914 38508
rect 6970 38452 7038 38508
rect 7094 38452 7104 38508
rect 5168 38442 7104 38452
rect 7874 39748 9810 39758
rect 7874 39692 7884 39748
rect 7940 39692 8008 39748
rect 8064 39692 8132 39748
rect 8188 39692 8256 39748
rect 8312 39692 8380 39748
rect 8436 39692 8504 39748
rect 8560 39692 8628 39748
rect 8684 39692 8752 39748
rect 8808 39692 8876 39748
rect 8932 39692 9000 39748
rect 9056 39692 9124 39748
rect 9180 39692 9248 39748
rect 9304 39692 9372 39748
rect 9428 39692 9496 39748
rect 9552 39692 9620 39748
rect 9676 39692 9744 39748
rect 9800 39692 9810 39748
rect 7874 39624 9810 39692
rect 7874 39568 7884 39624
rect 7940 39568 8008 39624
rect 8064 39568 8132 39624
rect 8188 39568 8256 39624
rect 8312 39568 8380 39624
rect 8436 39568 8504 39624
rect 8560 39568 8628 39624
rect 8684 39568 8752 39624
rect 8808 39568 8876 39624
rect 8932 39568 9000 39624
rect 9056 39568 9124 39624
rect 9180 39568 9248 39624
rect 9304 39568 9372 39624
rect 9428 39568 9496 39624
rect 9552 39568 9620 39624
rect 9676 39568 9744 39624
rect 9800 39568 9810 39624
rect 7874 39500 9810 39568
rect 7874 39444 7884 39500
rect 7940 39444 8008 39500
rect 8064 39444 8132 39500
rect 8188 39444 8256 39500
rect 8312 39444 8380 39500
rect 8436 39444 8504 39500
rect 8560 39444 8628 39500
rect 8684 39444 8752 39500
rect 8808 39444 8876 39500
rect 8932 39444 9000 39500
rect 9056 39444 9124 39500
rect 9180 39444 9248 39500
rect 9304 39444 9372 39500
rect 9428 39444 9496 39500
rect 9552 39444 9620 39500
rect 9676 39444 9744 39500
rect 9800 39444 9810 39500
rect 7874 39376 9810 39444
rect 7874 39320 7884 39376
rect 7940 39320 8008 39376
rect 8064 39320 8132 39376
rect 8188 39320 8256 39376
rect 8312 39320 8380 39376
rect 8436 39320 8504 39376
rect 8560 39320 8628 39376
rect 8684 39320 8752 39376
rect 8808 39320 8876 39376
rect 8932 39320 9000 39376
rect 9056 39320 9124 39376
rect 9180 39320 9248 39376
rect 9304 39320 9372 39376
rect 9428 39320 9496 39376
rect 9552 39320 9620 39376
rect 9676 39320 9744 39376
rect 9800 39320 9810 39376
rect 7874 39252 9810 39320
rect 7874 39196 7884 39252
rect 7940 39196 8008 39252
rect 8064 39196 8132 39252
rect 8188 39196 8256 39252
rect 8312 39196 8380 39252
rect 8436 39196 8504 39252
rect 8560 39196 8628 39252
rect 8684 39196 8752 39252
rect 8808 39196 8876 39252
rect 8932 39196 9000 39252
rect 9056 39196 9124 39252
rect 9180 39196 9248 39252
rect 9304 39196 9372 39252
rect 9428 39196 9496 39252
rect 9552 39196 9620 39252
rect 9676 39196 9744 39252
rect 9800 39196 9810 39252
rect 7874 39128 9810 39196
rect 7874 39072 7884 39128
rect 7940 39072 8008 39128
rect 8064 39072 8132 39128
rect 8188 39072 8256 39128
rect 8312 39072 8380 39128
rect 8436 39072 8504 39128
rect 8560 39072 8628 39128
rect 8684 39072 8752 39128
rect 8808 39072 8876 39128
rect 8932 39072 9000 39128
rect 9056 39072 9124 39128
rect 9180 39072 9248 39128
rect 9304 39072 9372 39128
rect 9428 39072 9496 39128
rect 9552 39072 9620 39128
rect 9676 39072 9744 39128
rect 9800 39072 9810 39128
rect 7874 39004 9810 39072
rect 7874 38948 7884 39004
rect 7940 38948 8008 39004
rect 8064 38948 8132 39004
rect 8188 38948 8256 39004
rect 8312 38948 8380 39004
rect 8436 38948 8504 39004
rect 8560 38948 8628 39004
rect 8684 38948 8752 39004
rect 8808 38948 8876 39004
rect 8932 38948 9000 39004
rect 9056 38948 9124 39004
rect 9180 38948 9248 39004
rect 9304 38948 9372 39004
rect 9428 38948 9496 39004
rect 9552 38948 9620 39004
rect 9676 38948 9744 39004
rect 9800 38948 9810 39004
rect 7874 38880 9810 38948
rect 7874 38824 7884 38880
rect 7940 38824 8008 38880
rect 8064 38824 8132 38880
rect 8188 38824 8256 38880
rect 8312 38824 8380 38880
rect 8436 38824 8504 38880
rect 8560 38824 8628 38880
rect 8684 38824 8752 38880
rect 8808 38824 8876 38880
rect 8932 38824 9000 38880
rect 9056 38824 9124 38880
rect 9180 38824 9248 38880
rect 9304 38824 9372 38880
rect 9428 38824 9496 38880
rect 9552 38824 9620 38880
rect 9676 38824 9744 38880
rect 9800 38824 9810 38880
rect 7874 38756 9810 38824
rect 7874 38700 7884 38756
rect 7940 38700 8008 38756
rect 8064 38700 8132 38756
rect 8188 38700 8256 38756
rect 8312 38700 8380 38756
rect 8436 38700 8504 38756
rect 8560 38700 8628 38756
rect 8684 38700 8752 38756
rect 8808 38700 8876 38756
rect 8932 38700 9000 38756
rect 9056 38700 9124 38756
rect 9180 38700 9248 38756
rect 9304 38700 9372 38756
rect 9428 38700 9496 38756
rect 9552 38700 9620 38756
rect 9676 38700 9744 38756
rect 9800 38700 9810 38756
rect 7874 38632 9810 38700
rect 7874 38576 7884 38632
rect 7940 38576 8008 38632
rect 8064 38576 8132 38632
rect 8188 38576 8256 38632
rect 8312 38576 8380 38632
rect 8436 38576 8504 38632
rect 8560 38576 8628 38632
rect 8684 38576 8752 38632
rect 8808 38576 8876 38632
rect 8932 38576 9000 38632
rect 9056 38576 9124 38632
rect 9180 38576 9248 38632
rect 9304 38576 9372 38632
rect 9428 38576 9496 38632
rect 9552 38576 9620 38632
rect 9676 38576 9744 38632
rect 9800 38576 9810 38632
rect 7874 38508 9810 38576
rect 7874 38452 7884 38508
rect 7940 38452 8008 38508
rect 8064 38452 8132 38508
rect 8188 38452 8256 38508
rect 8312 38452 8380 38508
rect 8436 38452 8504 38508
rect 8560 38452 8628 38508
rect 8684 38452 8752 38508
rect 8808 38452 8876 38508
rect 8932 38452 9000 38508
rect 9056 38452 9124 38508
rect 9180 38452 9248 38508
rect 9304 38452 9372 38508
rect 9428 38452 9496 38508
rect 9552 38452 9620 38508
rect 9676 38452 9744 38508
rect 9800 38452 9810 38508
rect 7874 38442 9810 38452
rect 10244 39748 12180 39758
rect 10244 39692 10254 39748
rect 10310 39692 10378 39748
rect 10434 39692 10502 39748
rect 10558 39692 10626 39748
rect 10682 39692 10750 39748
rect 10806 39692 10874 39748
rect 10930 39692 10998 39748
rect 11054 39692 11122 39748
rect 11178 39692 11246 39748
rect 11302 39692 11370 39748
rect 11426 39692 11494 39748
rect 11550 39692 11618 39748
rect 11674 39692 11742 39748
rect 11798 39692 11866 39748
rect 11922 39692 11990 39748
rect 12046 39692 12114 39748
rect 12170 39692 12180 39748
rect 10244 39624 12180 39692
rect 10244 39568 10254 39624
rect 10310 39568 10378 39624
rect 10434 39568 10502 39624
rect 10558 39568 10626 39624
rect 10682 39568 10750 39624
rect 10806 39568 10874 39624
rect 10930 39568 10998 39624
rect 11054 39568 11122 39624
rect 11178 39568 11246 39624
rect 11302 39568 11370 39624
rect 11426 39568 11494 39624
rect 11550 39568 11618 39624
rect 11674 39568 11742 39624
rect 11798 39568 11866 39624
rect 11922 39568 11990 39624
rect 12046 39568 12114 39624
rect 12170 39568 12180 39624
rect 10244 39500 12180 39568
rect 10244 39444 10254 39500
rect 10310 39444 10378 39500
rect 10434 39444 10502 39500
rect 10558 39444 10626 39500
rect 10682 39444 10750 39500
rect 10806 39444 10874 39500
rect 10930 39444 10998 39500
rect 11054 39444 11122 39500
rect 11178 39444 11246 39500
rect 11302 39444 11370 39500
rect 11426 39444 11494 39500
rect 11550 39444 11618 39500
rect 11674 39444 11742 39500
rect 11798 39444 11866 39500
rect 11922 39444 11990 39500
rect 12046 39444 12114 39500
rect 12170 39444 12180 39500
rect 10244 39376 12180 39444
rect 10244 39320 10254 39376
rect 10310 39320 10378 39376
rect 10434 39320 10502 39376
rect 10558 39320 10626 39376
rect 10682 39320 10750 39376
rect 10806 39320 10874 39376
rect 10930 39320 10998 39376
rect 11054 39320 11122 39376
rect 11178 39320 11246 39376
rect 11302 39320 11370 39376
rect 11426 39320 11494 39376
rect 11550 39320 11618 39376
rect 11674 39320 11742 39376
rect 11798 39320 11866 39376
rect 11922 39320 11990 39376
rect 12046 39320 12114 39376
rect 12170 39320 12180 39376
rect 10244 39252 12180 39320
rect 10244 39196 10254 39252
rect 10310 39196 10378 39252
rect 10434 39196 10502 39252
rect 10558 39196 10626 39252
rect 10682 39196 10750 39252
rect 10806 39196 10874 39252
rect 10930 39196 10998 39252
rect 11054 39196 11122 39252
rect 11178 39196 11246 39252
rect 11302 39196 11370 39252
rect 11426 39196 11494 39252
rect 11550 39196 11618 39252
rect 11674 39196 11742 39252
rect 11798 39196 11866 39252
rect 11922 39196 11990 39252
rect 12046 39196 12114 39252
rect 12170 39196 12180 39252
rect 10244 39128 12180 39196
rect 10244 39072 10254 39128
rect 10310 39072 10378 39128
rect 10434 39072 10502 39128
rect 10558 39072 10626 39128
rect 10682 39072 10750 39128
rect 10806 39072 10874 39128
rect 10930 39072 10998 39128
rect 11054 39072 11122 39128
rect 11178 39072 11246 39128
rect 11302 39072 11370 39128
rect 11426 39072 11494 39128
rect 11550 39072 11618 39128
rect 11674 39072 11742 39128
rect 11798 39072 11866 39128
rect 11922 39072 11990 39128
rect 12046 39072 12114 39128
rect 12170 39072 12180 39128
rect 10244 39004 12180 39072
rect 10244 38948 10254 39004
rect 10310 38948 10378 39004
rect 10434 38948 10502 39004
rect 10558 38948 10626 39004
rect 10682 38948 10750 39004
rect 10806 38948 10874 39004
rect 10930 38948 10998 39004
rect 11054 38948 11122 39004
rect 11178 38948 11246 39004
rect 11302 38948 11370 39004
rect 11426 38948 11494 39004
rect 11550 38948 11618 39004
rect 11674 38948 11742 39004
rect 11798 38948 11866 39004
rect 11922 38948 11990 39004
rect 12046 38948 12114 39004
rect 12170 38948 12180 39004
rect 10244 38880 12180 38948
rect 10244 38824 10254 38880
rect 10310 38824 10378 38880
rect 10434 38824 10502 38880
rect 10558 38824 10626 38880
rect 10682 38824 10750 38880
rect 10806 38824 10874 38880
rect 10930 38824 10998 38880
rect 11054 38824 11122 38880
rect 11178 38824 11246 38880
rect 11302 38824 11370 38880
rect 11426 38824 11494 38880
rect 11550 38824 11618 38880
rect 11674 38824 11742 38880
rect 11798 38824 11866 38880
rect 11922 38824 11990 38880
rect 12046 38824 12114 38880
rect 12170 38824 12180 38880
rect 10244 38756 12180 38824
rect 10244 38700 10254 38756
rect 10310 38700 10378 38756
rect 10434 38700 10502 38756
rect 10558 38700 10626 38756
rect 10682 38700 10750 38756
rect 10806 38700 10874 38756
rect 10930 38700 10998 38756
rect 11054 38700 11122 38756
rect 11178 38700 11246 38756
rect 11302 38700 11370 38756
rect 11426 38700 11494 38756
rect 11550 38700 11618 38756
rect 11674 38700 11742 38756
rect 11798 38700 11866 38756
rect 11922 38700 11990 38756
rect 12046 38700 12114 38756
rect 12170 38700 12180 38756
rect 10244 38632 12180 38700
rect 10244 38576 10254 38632
rect 10310 38576 10378 38632
rect 10434 38576 10502 38632
rect 10558 38576 10626 38632
rect 10682 38576 10750 38632
rect 10806 38576 10874 38632
rect 10930 38576 10998 38632
rect 11054 38576 11122 38632
rect 11178 38576 11246 38632
rect 11302 38576 11370 38632
rect 11426 38576 11494 38632
rect 11550 38576 11618 38632
rect 11674 38576 11742 38632
rect 11798 38576 11866 38632
rect 11922 38576 11990 38632
rect 12046 38576 12114 38632
rect 12170 38576 12180 38632
rect 10244 38508 12180 38576
rect 10244 38452 10254 38508
rect 10310 38452 10378 38508
rect 10434 38452 10502 38508
rect 10558 38452 10626 38508
rect 10682 38452 10750 38508
rect 10806 38452 10874 38508
rect 10930 38452 10998 38508
rect 11054 38452 11122 38508
rect 11178 38452 11246 38508
rect 11302 38452 11370 38508
rect 11426 38452 11494 38508
rect 11550 38452 11618 38508
rect 11674 38452 11742 38508
rect 11798 38452 11866 38508
rect 11922 38452 11990 38508
rect 12046 38452 12114 38508
rect 12170 38452 12180 38508
rect 10244 38442 12180 38452
rect 12861 39748 14673 39758
rect 12861 39692 12871 39748
rect 12927 39692 12995 39748
rect 13051 39692 13119 39748
rect 13175 39692 13243 39748
rect 13299 39692 13367 39748
rect 13423 39692 13491 39748
rect 13547 39692 13615 39748
rect 13671 39692 13739 39748
rect 13795 39692 13863 39748
rect 13919 39692 13987 39748
rect 14043 39692 14111 39748
rect 14167 39692 14235 39748
rect 14291 39692 14359 39748
rect 14415 39692 14483 39748
rect 14539 39692 14607 39748
rect 14663 39692 14673 39748
rect 12861 39624 14673 39692
rect 12861 39568 12871 39624
rect 12927 39568 12995 39624
rect 13051 39568 13119 39624
rect 13175 39568 13243 39624
rect 13299 39568 13367 39624
rect 13423 39568 13491 39624
rect 13547 39568 13615 39624
rect 13671 39568 13739 39624
rect 13795 39568 13863 39624
rect 13919 39568 13987 39624
rect 14043 39568 14111 39624
rect 14167 39568 14235 39624
rect 14291 39568 14359 39624
rect 14415 39568 14483 39624
rect 14539 39568 14607 39624
rect 14663 39568 14673 39624
rect 12861 39500 14673 39568
rect 12861 39444 12871 39500
rect 12927 39444 12995 39500
rect 13051 39444 13119 39500
rect 13175 39444 13243 39500
rect 13299 39444 13367 39500
rect 13423 39444 13491 39500
rect 13547 39444 13615 39500
rect 13671 39444 13739 39500
rect 13795 39444 13863 39500
rect 13919 39444 13987 39500
rect 14043 39444 14111 39500
rect 14167 39444 14235 39500
rect 14291 39444 14359 39500
rect 14415 39444 14483 39500
rect 14539 39444 14607 39500
rect 14663 39444 14673 39500
rect 12861 39376 14673 39444
rect 12861 39320 12871 39376
rect 12927 39320 12995 39376
rect 13051 39320 13119 39376
rect 13175 39320 13243 39376
rect 13299 39320 13367 39376
rect 13423 39320 13491 39376
rect 13547 39320 13615 39376
rect 13671 39320 13739 39376
rect 13795 39320 13863 39376
rect 13919 39320 13987 39376
rect 14043 39320 14111 39376
rect 14167 39320 14235 39376
rect 14291 39320 14359 39376
rect 14415 39320 14483 39376
rect 14539 39320 14607 39376
rect 14663 39320 14673 39376
rect 12861 39252 14673 39320
rect 12861 39196 12871 39252
rect 12927 39196 12995 39252
rect 13051 39196 13119 39252
rect 13175 39196 13243 39252
rect 13299 39196 13367 39252
rect 13423 39196 13491 39252
rect 13547 39196 13615 39252
rect 13671 39196 13739 39252
rect 13795 39196 13863 39252
rect 13919 39196 13987 39252
rect 14043 39196 14111 39252
rect 14167 39196 14235 39252
rect 14291 39196 14359 39252
rect 14415 39196 14483 39252
rect 14539 39196 14607 39252
rect 14663 39196 14673 39252
rect 12861 39128 14673 39196
rect 12861 39072 12871 39128
rect 12927 39072 12995 39128
rect 13051 39072 13119 39128
rect 13175 39072 13243 39128
rect 13299 39072 13367 39128
rect 13423 39072 13491 39128
rect 13547 39072 13615 39128
rect 13671 39072 13739 39128
rect 13795 39072 13863 39128
rect 13919 39072 13987 39128
rect 14043 39072 14111 39128
rect 14167 39072 14235 39128
rect 14291 39072 14359 39128
rect 14415 39072 14483 39128
rect 14539 39072 14607 39128
rect 14663 39072 14673 39128
rect 12861 39004 14673 39072
rect 12861 38948 12871 39004
rect 12927 38948 12995 39004
rect 13051 38948 13119 39004
rect 13175 38948 13243 39004
rect 13299 38948 13367 39004
rect 13423 38948 13491 39004
rect 13547 38948 13615 39004
rect 13671 38948 13739 39004
rect 13795 38948 13863 39004
rect 13919 38948 13987 39004
rect 14043 38948 14111 39004
rect 14167 38948 14235 39004
rect 14291 38948 14359 39004
rect 14415 38948 14483 39004
rect 14539 38948 14607 39004
rect 14663 38948 14673 39004
rect 12861 38880 14673 38948
rect 12861 38824 12871 38880
rect 12927 38824 12995 38880
rect 13051 38824 13119 38880
rect 13175 38824 13243 38880
rect 13299 38824 13367 38880
rect 13423 38824 13491 38880
rect 13547 38824 13615 38880
rect 13671 38824 13739 38880
rect 13795 38824 13863 38880
rect 13919 38824 13987 38880
rect 14043 38824 14111 38880
rect 14167 38824 14235 38880
rect 14291 38824 14359 38880
rect 14415 38824 14483 38880
rect 14539 38824 14607 38880
rect 14663 38824 14673 38880
rect 12861 38756 14673 38824
rect 12861 38700 12871 38756
rect 12927 38700 12995 38756
rect 13051 38700 13119 38756
rect 13175 38700 13243 38756
rect 13299 38700 13367 38756
rect 13423 38700 13491 38756
rect 13547 38700 13615 38756
rect 13671 38700 13739 38756
rect 13795 38700 13863 38756
rect 13919 38700 13987 38756
rect 14043 38700 14111 38756
rect 14167 38700 14235 38756
rect 14291 38700 14359 38756
rect 14415 38700 14483 38756
rect 14539 38700 14607 38756
rect 14663 38700 14673 38756
rect 12861 38632 14673 38700
rect 12861 38576 12871 38632
rect 12927 38576 12995 38632
rect 13051 38576 13119 38632
rect 13175 38576 13243 38632
rect 13299 38576 13367 38632
rect 13423 38576 13491 38632
rect 13547 38576 13615 38632
rect 13671 38576 13739 38632
rect 13795 38576 13863 38632
rect 13919 38576 13987 38632
rect 14043 38576 14111 38632
rect 14167 38576 14235 38632
rect 14291 38576 14359 38632
rect 14415 38576 14483 38632
rect 14539 38576 14607 38632
rect 14663 38576 14673 38632
rect 12861 38508 14673 38576
rect 12861 38452 12871 38508
rect 12927 38452 12995 38508
rect 13051 38452 13119 38508
rect 13175 38452 13243 38508
rect 13299 38452 13367 38508
rect 13423 38452 13491 38508
rect 13547 38452 13615 38508
rect 13671 38452 13739 38508
rect 13795 38452 13863 38508
rect 13919 38452 13987 38508
rect 14043 38452 14111 38508
rect 14167 38452 14235 38508
rect 14291 38452 14359 38508
rect 14415 38452 14483 38508
rect 14539 38452 14607 38508
rect 14663 38452 14673 38508
rect 12861 38442 14673 38452
rect 14892 38176 14989 38200
rect 2279 38079 2289 38135
rect 2345 38079 2355 38135
rect 2279 38003 2355 38079
rect 2279 37947 2289 38003
rect 2345 37947 2355 38003
rect 2279 37871 2355 37947
rect 2279 37815 2289 37871
rect 2345 37815 2355 37871
rect 2279 37739 2355 37815
rect 2279 37683 2289 37739
rect 2345 37683 2355 37739
rect 2279 37607 2355 37683
rect 2279 37551 2289 37607
rect 2345 37551 2355 37607
rect 2279 37475 2355 37551
rect 2279 37419 2289 37475
rect 2345 37419 2355 37475
rect 2279 37343 2355 37419
rect 2279 37287 2289 37343
rect 2345 37287 2355 37343
rect 2279 37211 2355 37287
rect 2279 37155 2289 37211
rect 2345 37155 2355 37211
rect 2279 37079 2355 37155
rect 2279 37023 2289 37079
rect 2345 37023 2355 37079
rect 2279 36947 2355 37023
rect 2279 36891 2289 36947
rect 2345 36891 2355 36947
rect 2279 36800 2355 36891
rect 14892 36824 14902 38176
rect 14958 36824 14989 38176
rect 14892 36800 14989 36824
rect 2481 33636 2681 36564
rect 4851 33636 5051 36564
rect 7265 33636 7713 36564
rect 9927 33636 10127 36564
rect 12297 33636 12497 36564
rect 305 30436 2117 33364
rect 2798 30436 4734 33364
rect 5168 30436 7104 33364
rect 7874 30436 9810 33364
rect 10244 30436 12180 33364
rect 12861 30436 14673 33364
rect 305 28842 2117 30158
rect 2798 28842 4734 30158
rect 5168 28842 7104 30158
rect 7874 28842 9810 30158
rect 10244 28842 12180 30158
rect 12861 28842 14673 30158
rect 2481 27242 2681 28558
rect 4851 27242 5051 28558
rect 7265 27242 7713 28558
rect 9927 27242 10127 28558
rect 12297 27242 12497 28558
rect 305 24036 2117 26964
rect 2798 24036 4734 26964
rect 5168 24036 7104 26964
rect 7874 24036 9810 26964
rect 10244 24036 12180 26964
rect 12861 24036 14673 26964
rect 305 20836 2117 23764
rect 2798 20836 4734 23764
rect 5168 20836 7104 23764
rect 7874 20836 9810 23764
rect 10244 20836 12180 23764
rect 12861 20836 14673 23764
rect 305 17636 2117 20564
rect 2798 17636 4734 20564
rect 5168 17636 7104 20564
rect 7874 17636 9810 20564
rect 10244 17636 12180 20564
rect 12861 17636 14673 20564
rect 305 14436 2117 17364
rect 2798 14436 4734 17364
rect 5168 14436 7104 17364
rect 7874 14436 9810 17364
rect 10244 14436 12180 17364
rect 12861 14436 14673 17364
rect 2481 12842 2681 14158
rect 4851 12842 5051 14158
rect 7265 12842 7713 14158
rect 9927 12842 10127 14158
rect 12297 12842 12497 14158
rect 305 11242 2117 12558
rect 2798 11242 4734 12558
rect 5168 11242 7104 12558
rect 7874 11242 9810 12558
rect 10244 11242 12180 12558
rect 12861 11242 14673 12558
rect 2481 8036 2681 10964
rect 4851 8036 5051 10964
rect 7265 8036 7713 10964
rect 9927 8036 10127 10964
rect 12297 8036 12497 10964
rect 2481 4836 2681 7764
rect 4851 4836 5051 7764
rect 7265 4836 7713 7764
rect 9927 4836 10127 7764
rect 12297 4836 12497 7764
rect 2481 1636 2681 4564
rect 4851 1636 5051 4564
rect 7265 1636 7713 4564
rect 9927 1636 10127 4564
rect 12297 1636 12497 4564
rect 261 0 2161 1190
rect 2741 0 4791 1190
rect 5111 0 7161 1190
rect 7817 0 9867 1190
rect 10187 0 12237 1190
rect 12817 0 14717 1190
<< via2 >>
rect 20 52574 76 52576
rect 20 52522 22 52574
rect 22 52522 74 52574
rect 74 52522 76 52574
rect 20 52466 76 52522
rect 20 52414 22 52466
rect 22 52414 74 52466
rect 74 52414 76 52466
rect 20 52358 76 52414
rect 20 52306 22 52358
rect 22 52306 74 52358
rect 74 52306 76 52358
rect 20 52250 76 52306
rect 20 52198 22 52250
rect 22 52198 74 52250
rect 74 52198 76 52250
rect 20 52142 76 52198
rect 20 52090 22 52142
rect 22 52090 74 52142
rect 74 52090 76 52142
rect 20 52034 76 52090
rect 20 51982 22 52034
rect 22 51982 74 52034
rect 74 51982 76 52034
rect 20 51926 76 51982
rect 20 51874 22 51926
rect 22 51874 74 51926
rect 74 51874 76 51926
rect 20 51818 76 51874
rect 20 51766 22 51818
rect 22 51766 74 51818
rect 74 51766 76 51818
rect 20 51710 76 51766
rect 20 51658 22 51710
rect 22 51658 74 51710
rect 74 51658 76 51710
rect 20 51602 76 51658
rect 20 51550 22 51602
rect 22 51550 74 51602
rect 74 51550 76 51602
rect 20 51494 76 51550
rect 20 51442 22 51494
rect 22 51442 74 51494
rect 74 51442 76 51494
rect 20 51386 76 51442
rect 20 51334 22 51386
rect 22 51334 74 51386
rect 74 51334 76 51386
rect 20 51278 76 51334
rect 20 51226 22 51278
rect 22 51226 74 51278
rect 74 51226 76 51278
rect 20 51224 76 51226
rect 315 50892 371 50948
rect 439 50892 495 50948
rect 563 50892 619 50948
rect 687 50892 743 50948
rect 811 50892 867 50948
rect 935 50892 991 50948
rect 1059 50892 1115 50948
rect 1183 50892 1239 50948
rect 1307 50892 1363 50948
rect 1431 50892 1487 50948
rect 1555 50892 1611 50948
rect 1679 50892 1735 50948
rect 1803 50892 1859 50948
rect 1927 50892 1983 50948
rect 2051 50892 2107 50948
rect 315 50768 371 50824
rect 439 50768 495 50824
rect 563 50768 619 50824
rect 687 50768 743 50824
rect 811 50768 867 50824
rect 935 50768 991 50824
rect 1059 50768 1115 50824
rect 1183 50768 1239 50824
rect 1307 50768 1363 50824
rect 1431 50768 1487 50824
rect 1555 50768 1611 50824
rect 1679 50768 1735 50824
rect 1803 50768 1859 50824
rect 1927 50768 1983 50824
rect 2051 50768 2107 50824
rect 315 50644 371 50700
rect 439 50644 495 50700
rect 563 50644 619 50700
rect 687 50644 743 50700
rect 811 50644 867 50700
rect 935 50644 991 50700
rect 1059 50644 1115 50700
rect 1183 50644 1239 50700
rect 1307 50644 1363 50700
rect 1431 50644 1487 50700
rect 1555 50644 1611 50700
rect 1679 50644 1735 50700
rect 1803 50644 1859 50700
rect 1927 50644 1983 50700
rect 2051 50644 2107 50700
rect 315 50520 371 50576
rect 439 50520 495 50576
rect 563 50520 619 50576
rect 687 50520 743 50576
rect 811 50520 867 50576
rect 935 50520 991 50576
rect 1059 50520 1115 50576
rect 1183 50520 1239 50576
rect 1307 50520 1363 50576
rect 1431 50520 1487 50576
rect 1555 50520 1611 50576
rect 1679 50520 1735 50576
rect 1803 50520 1859 50576
rect 1927 50520 1983 50576
rect 2051 50520 2107 50576
rect 315 50396 371 50452
rect 439 50396 495 50452
rect 563 50396 619 50452
rect 687 50396 743 50452
rect 811 50396 867 50452
rect 935 50396 991 50452
rect 1059 50396 1115 50452
rect 1183 50396 1239 50452
rect 1307 50396 1363 50452
rect 1431 50396 1487 50452
rect 1555 50396 1611 50452
rect 1679 50396 1735 50452
rect 1803 50396 1859 50452
rect 1927 50396 1983 50452
rect 2051 50396 2107 50452
rect 315 50272 371 50328
rect 439 50272 495 50328
rect 563 50272 619 50328
rect 687 50272 743 50328
rect 811 50272 867 50328
rect 935 50272 991 50328
rect 1059 50272 1115 50328
rect 1183 50272 1239 50328
rect 1307 50272 1363 50328
rect 1431 50272 1487 50328
rect 1555 50272 1611 50328
rect 1679 50272 1735 50328
rect 1803 50272 1859 50328
rect 1927 50272 1983 50328
rect 2051 50272 2107 50328
rect 315 50148 371 50204
rect 439 50148 495 50204
rect 563 50148 619 50204
rect 687 50148 743 50204
rect 811 50148 867 50204
rect 935 50148 991 50204
rect 1059 50148 1115 50204
rect 1183 50148 1239 50204
rect 1307 50148 1363 50204
rect 1431 50148 1487 50204
rect 1555 50148 1611 50204
rect 1679 50148 1735 50204
rect 1803 50148 1859 50204
rect 1927 50148 1983 50204
rect 2051 50148 2107 50204
rect 315 50024 371 50080
rect 439 50024 495 50080
rect 563 50024 619 50080
rect 687 50024 743 50080
rect 811 50024 867 50080
rect 935 50024 991 50080
rect 1059 50024 1115 50080
rect 1183 50024 1239 50080
rect 1307 50024 1363 50080
rect 1431 50024 1487 50080
rect 1555 50024 1611 50080
rect 1679 50024 1735 50080
rect 1803 50024 1859 50080
rect 1927 50024 1983 50080
rect 2051 50024 2107 50080
rect 315 49900 371 49956
rect 439 49900 495 49956
rect 563 49900 619 49956
rect 687 49900 743 49956
rect 811 49900 867 49956
rect 935 49900 991 49956
rect 1059 49900 1115 49956
rect 1183 49900 1239 49956
rect 1307 49900 1363 49956
rect 1431 49900 1487 49956
rect 1555 49900 1611 49956
rect 1679 49900 1735 49956
rect 1803 49900 1859 49956
rect 1927 49900 1983 49956
rect 2051 49900 2107 49956
rect 315 49776 371 49832
rect 439 49776 495 49832
rect 563 49776 619 49832
rect 687 49776 743 49832
rect 811 49776 867 49832
rect 935 49776 991 49832
rect 1059 49776 1115 49832
rect 1183 49776 1239 49832
rect 1307 49776 1363 49832
rect 1431 49776 1487 49832
rect 1555 49776 1611 49832
rect 1679 49776 1735 49832
rect 1803 49776 1859 49832
rect 1927 49776 1983 49832
rect 2051 49776 2107 49832
rect 315 49652 371 49708
rect 439 49652 495 49708
rect 563 49652 619 49708
rect 687 49652 743 49708
rect 811 49652 867 49708
rect 935 49652 991 49708
rect 1059 49652 1115 49708
rect 1183 49652 1239 49708
rect 1307 49652 1363 49708
rect 1431 49652 1487 49708
rect 1555 49652 1611 49708
rect 1679 49652 1735 49708
rect 1803 49652 1859 49708
rect 1927 49652 1983 49708
rect 2051 49652 2107 49708
rect 2289 52465 2345 52521
rect 2289 52333 2345 52389
rect 2289 52201 2345 52257
rect 2289 52069 2345 52125
rect 2289 51937 2345 51993
rect 2289 51805 2345 51861
rect 2289 51673 2345 51729
rect 2289 51541 2345 51597
rect 2289 51409 2345 51465
rect 2289 51277 2345 51333
rect 315 39692 371 39748
rect 439 39692 495 39748
rect 563 39692 619 39748
rect 687 39692 743 39748
rect 811 39692 867 39748
rect 935 39692 991 39748
rect 1059 39692 1115 39748
rect 1183 39692 1239 39748
rect 1307 39692 1363 39748
rect 1431 39692 1487 39748
rect 1555 39692 1611 39748
rect 1679 39692 1735 39748
rect 1803 39692 1859 39748
rect 1927 39692 1983 39748
rect 2051 39692 2107 39748
rect 315 39568 371 39624
rect 439 39568 495 39624
rect 563 39568 619 39624
rect 687 39568 743 39624
rect 811 39568 867 39624
rect 935 39568 991 39624
rect 1059 39568 1115 39624
rect 1183 39568 1239 39624
rect 1307 39568 1363 39624
rect 1431 39568 1487 39624
rect 1555 39568 1611 39624
rect 1679 39568 1735 39624
rect 1803 39568 1859 39624
rect 1927 39568 1983 39624
rect 2051 39568 2107 39624
rect 315 39444 371 39500
rect 439 39444 495 39500
rect 563 39444 619 39500
rect 687 39444 743 39500
rect 811 39444 867 39500
rect 935 39444 991 39500
rect 1059 39444 1115 39500
rect 1183 39444 1239 39500
rect 1307 39444 1363 39500
rect 1431 39444 1487 39500
rect 1555 39444 1611 39500
rect 1679 39444 1735 39500
rect 1803 39444 1859 39500
rect 1927 39444 1983 39500
rect 2051 39444 2107 39500
rect 315 39320 371 39376
rect 439 39320 495 39376
rect 563 39320 619 39376
rect 687 39320 743 39376
rect 811 39320 867 39376
rect 935 39320 991 39376
rect 1059 39320 1115 39376
rect 1183 39320 1239 39376
rect 1307 39320 1363 39376
rect 1431 39320 1487 39376
rect 1555 39320 1611 39376
rect 1679 39320 1735 39376
rect 1803 39320 1859 39376
rect 1927 39320 1983 39376
rect 2051 39320 2107 39376
rect 315 39196 371 39252
rect 439 39196 495 39252
rect 563 39196 619 39252
rect 687 39196 743 39252
rect 811 39196 867 39252
rect 935 39196 991 39252
rect 1059 39196 1115 39252
rect 1183 39196 1239 39252
rect 1307 39196 1363 39252
rect 1431 39196 1487 39252
rect 1555 39196 1611 39252
rect 1679 39196 1735 39252
rect 1803 39196 1859 39252
rect 1927 39196 1983 39252
rect 2051 39196 2107 39252
rect 315 39072 371 39128
rect 439 39072 495 39128
rect 563 39072 619 39128
rect 687 39072 743 39128
rect 811 39072 867 39128
rect 935 39072 991 39128
rect 1059 39072 1115 39128
rect 1183 39072 1239 39128
rect 1307 39072 1363 39128
rect 1431 39072 1487 39128
rect 1555 39072 1611 39128
rect 1679 39072 1735 39128
rect 1803 39072 1859 39128
rect 1927 39072 1983 39128
rect 2051 39072 2107 39128
rect 315 38948 371 39004
rect 439 38948 495 39004
rect 563 38948 619 39004
rect 687 38948 743 39004
rect 811 38948 867 39004
rect 935 38948 991 39004
rect 1059 38948 1115 39004
rect 1183 38948 1239 39004
rect 1307 38948 1363 39004
rect 1431 38948 1487 39004
rect 1555 38948 1611 39004
rect 1679 38948 1735 39004
rect 1803 38948 1859 39004
rect 1927 38948 1983 39004
rect 2051 38948 2107 39004
rect 315 38824 371 38880
rect 439 38824 495 38880
rect 563 38824 619 38880
rect 687 38824 743 38880
rect 811 38824 867 38880
rect 935 38824 991 38880
rect 1059 38824 1115 38880
rect 1183 38824 1239 38880
rect 1307 38824 1363 38880
rect 1431 38824 1487 38880
rect 1555 38824 1611 38880
rect 1679 38824 1735 38880
rect 1803 38824 1859 38880
rect 1927 38824 1983 38880
rect 2051 38824 2107 38880
rect 315 38700 371 38756
rect 439 38700 495 38756
rect 563 38700 619 38756
rect 687 38700 743 38756
rect 811 38700 867 38756
rect 935 38700 991 38756
rect 1059 38700 1115 38756
rect 1183 38700 1239 38756
rect 1307 38700 1363 38756
rect 1431 38700 1487 38756
rect 1555 38700 1611 38756
rect 1679 38700 1735 38756
rect 1803 38700 1859 38756
rect 1927 38700 1983 38756
rect 2051 38700 2107 38756
rect 315 38576 371 38632
rect 439 38576 495 38632
rect 563 38576 619 38632
rect 687 38576 743 38632
rect 811 38576 867 38632
rect 935 38576 991 38632
rect 1059 38576 1115 38632
rect 1183 38576 1239 38632
rect 1307 38576 1363 38632
rect 1431 38576 1487 38632
rect 1555 38576 1611 38632
rect 1679 38576 1735 38632
rect 1803 38576 1859 38632
rect 1927 38576 1983 38632
rect 2051 38576 2107 38632
rect 315 38452 371 38508
rect 439 38452 495 38508
rect 563 38452 619 38508
rect 687 38452 743 38508
rect 811 38452 867 38508
rect 935 38452 991 38508
rect 1059 38452 1115 38508
rect 1183 38452 1239 38508
rect 1307 38452 1363 38508
rect 1431 38452 1487 38508
rect 1555 38452 1611 38508
rect 1679 38452 1735 38508
rect 1803 38452 1859 38508
rect 1927 38452 1983 38508
rect 2051 38452 2107 38508
rect 20 38174 76 38176
rect 20 38122 22 38174
rect 22 38122 74 38174
rect 74 38122 76 38174
rect 20 38066 76 38122
rect 20 38014 22 38066
rect 22 38014 74 38066
rect 74 38014 76 38066
rect 20 37958 76 38014
rect 20 37906 22 37958
rect 22 37906 74 37958
rect 74 37906 76 37958
rect 20 37850 76 37906
rect 20 37798 22 37850
rect 22 37798 74 37850
rect 74 37798 76 37850
rect 20 37742 76 37798
rect 20 37690 22 37742
rect 22 37690 74 37742
rect 74 37690 76 37742
rect 20 37634 76 37690
rect 20 37582 22 37634
rect 22 37582 74 37634
rect 74 37582 76 37634
rect 20 37526 76 37582
rect 20 37474 22 37526
rect 22 37474 74 37526
rect 74 37474 76 37526
rect 20 37418 76 37474
rect 20 37366 22 37418
rect 22 37366 74 37418
rect 74 37366 76 37418
rect 20 37310 76 37366
rect 20 37258 22 37310
rect 22 37258 74 37310
rect 74 37258 76 37310
rect 20 37202 76 37258
rect 20 37150 22 37202
rect 22 37150 74 37202
rect 74 37150 76 37202
rect 20 37094 76 37150
rect 20 37042 22 37094
rect 22 37042 74 37094
rect 74 37042 76 37094
rect 20 36986 76 37042
rect 20 36934 22 36986
rect 22 36934 74 36986
rect 74 36934 76 36986
rect 20 36878 76 36934
rect 20 36826 22 36878
rect 22 36826 74 36878
rect 74 36826 76 36878
rect 20 36824 76 36826
rect 2491 52492 2547 52548
rect 2615 52492 2671 52548
rect 2491 52368 2547 52424
rect 2615 52368 2671 52424
rect 2491 52244 2547 52300
rect 2615 52244 2671 52300
rect 2491 52120 2547 52176
rect 2615 52120 2671 52176
rect 2491 51996 2547 52052
rect 2615 51996 2671 52052
rect 2491 51872 2547 51928
rect 2615 51872 2671 51928
rect 2491 51748 2547 51804
rect 2615 51748 2671 51804
rect 2491 51624 2547 51680
rect 2615 51624 2671 51680
rect 2491 51500 2547 51556
rect 2615 51500 2671 51556
rect 2491 51376 2547 51432
rect 2615 51376 2671 51432
rect 2491 51252 2547 51308
rect 2615 51252 2671 51308
rect 2808 50892 2864 50948
rect 2932 50892 2988 50948
rect 3056 50892 3112 50948
rect 3180 50892 3236 50948
rect 3304 50892 3360 50948
rect 3428 50892 3484 50948
rect 3552 50892 3608 50948
rect 3676 50892 3732 50948
rect 3800 50892 3856 50948
rect 3924 50892 3980 50948
rect 4048 50892 4104 50948
rect 4172 50892 4228 50948
rect 4296 50892 4352 50948
rect 4420 50892 4476 50948
rect 4544 50892 4600 50948
rect 4668 50892 4724 50948
rect 2808 50768 2864 50824
rect 2932 50768 2988 50824
rect 3056 50768 3112 50824
rect 3180 50768 3236 50824
rect 3304 50768 3360 50824
rect 3428 50768 3484 50824
rect 3552 50768 3608 50824
rect 3676 50768 3732 50824
rect 3800 50768 3856 50824
rect 3924 50768 3980 50824
rect 4048 50768 4104 50824
rect 4172 50768 4228 50824
rect 4296 50768 4352 50824
rect 4420 50768 4476 50824
rect 4544 50768 4600 50824
rect 4668 50768 4724 50824
rect 2808 50644 2864 50700
rect 2932 50644 2988 50700
rect 3056 50644 3112 50700
rect 3180 50644 3236 50700
rect 3304 50644 3360 50700
rect 3428 50644 3484 50700
rect 3552 50693 3608 50700
rect 3676 50693 3732 50700
rect 3800 50693 3856 50700
rect 3924 50693 3980 50700
rect 4048 50693 4104 50700
rect 4172 50693 4228 50700
rect 4296 50693 4352 50700
rect 4420 50693 4476 50700
rect 4544 50693 4600 50700
rect 4668 50693 4724 50700
rect 3552 50644 3559 50693
rect 3559 50644 3608 50693
rect 3676 50644 3683 50693
rect 3683 50644 3732 50693
rect 3800 50644 3807 50693
rect 3807 50644 3856 50693
rect 3924 50644 3931 50693
rect 3931 50644 3980 50693
rect 4048 50644 4055 50693
rect 4055 50644 4104 50693
rect 4172 50644 4179 50693
rect 4179 50644 4228 50693
rect 4296 50644 4303 50693
rect 4303 50644 4352 50693
rect 4420 50644 4427 50693
rect 4427 50644 4476 50693
rect 4544 50644 4551 50693
rect 4551 50644 4600 50693
rect 4668 50644 4675 50693
rect 4675 50644 4724 50693
rect 2808 50520 2864 50576
rect 2932 50520 2988 50576
rect 3056 50520 3112 50576
rect 3180 50520 3236 50576
rect 3304 50520 3360 50576
rect 3428 50520 3484 50576
rect 3552 50569 3608 50576
rect 3676 50569 3732 50576
rect 3800 50569 3856 50576
rect 3924 50569 3980 50576
rect 4048 50569 4104 50576
rect 4172 50569 4228 50576
rect 4296 50569 4352 50576
rect 4420 50569 4476 50576
rect 4544 50569 4600 50576
rect 4668 50569 4724 50576
rect 3552 50520 3559 50569
rect 3559 50520 3608 50569
rect 3676 50520 3683 50569
rect 3683 50520 3732 50569
rect 3800 50520 3807 50569
rect 3807 50520 3856 50569
rect 3924 50520 3931 50569
rect 3931 50520 3980 50569
rect 4048 50520 4055 50569
rect 4055 50520 4104 50569
rect 4172 50520 4179 50569
rect 4179 50520 4228 50569
rect 4296 50520 4303 50569
rect 4303 50520 4352 50569
rect 4420 50520 4427 50569
rect 4427 50520 4476 50569
rect 4544 50520 4551 50569
rect 4551 50520 4600 50569
rect 4668 50520 4675 50569
rect 4675 50520 4724 50569
rect 2808 50396 2864 50452
rect 2932 50396 2988 50452
rect 3056 50396 3112 50452
rect 3180 50396 3236 50452
rect 3304 50396 3360 50452
rect 3428 50396 3484 50452
rect 3552 50396 3608 50452
rect 3676 50396 3732 50452
rect 3800 50396 3856 50452
rect 3924 50396 3980 50452
rect 4048 50396 4104 50452
rect 4172 50396 4228 50452
rect 4296 50396 4352 50452
rect 4420 50396 4476 50452
rect 4544 50396 4600 50452
rect 4668 50396 4724 50452
rect 2808 50272 2864 50328
rect 2932 50272 2988 50328
rect 3056 50272 3112 50328
rect 3180 50272 3236 50328
rect 3304 50272 3360 50328
rect 3428 50272 3484 50328
rect 3552 50272 3608 50328
rect 3676 50272 3732 50328
rect 3800 50272 3856 50328
rect 3924 50272 3980 50328
rect 4048 50272 4104 50328
rect 4172 50272 4228 50328
rect 4296 50272 4352 50328
rect 4420 50272 4476 50328
rect 4544 50272 4600 50328
rect 4668 50272 4724 50328
rect 2808 50148 2864 50204
rect 2932 50148 2988 50204
rect 3056 50148 3112 50204
rect 3180 50148 3236 50204
rect 3304 50148 3360 50204
rect 3428 50148 3484 50204
rect 3552 50148 3608 50204
rect 3676 50148 3732 50204
rect 3800 50148 3856 50204
rect 3924 50148 3980 50204
rect 4048 50148 4104 50204
rect 4172 50148 4228 50204
rect 4296 50148 4352 50204
rect 4420 50148 4476 50204
rect 4544 50148 4600 50204
rect 4668 50148 4724 50204
rect 2808 50024 2864 50080
rect 2932 50024 2988 50080
rect 3056 50024 3112 50080
rect 3180 50024 3236 50080
rect 3304 50024 3360 50080
rect 3428 50024 3484 50080
rect 3552 50024 3608 50080
rect 3676 50024 3732 50080
rect 3800 50024 3856 50080
rect 3924 50024 3980 50080
rect 4048 50024 4104 50080
rect 4172 50024 4228 50080
rect 4296 50024 4352 50080
rect 4420 50024 4476 50080
rect 4544 50024 4600 50080
rect 4668 50024 4724 50080
rect 2808 49900 2864 49956
rect 2932 49900 2988 49956
rect 3056 49900 3112 49956
rect 3180 49900 3236 49956
rect 3304 49900 3360 49956
rect 3428 49900 3484 49956
rect 3552 49900 3608 49956
rect 3676 49900 3732 49956
rect 3800 49900 3856 49956
rect 3924 49900 3980 49956
rect 4048 49900 4104 49956
rect 4172 49900 4228 49956
rect 4296 49900 4352 49956
rect 4420 49900 4476 49956
rect 4544 49900 4600 49956
rect 4668 49900 4724 49956
rect 2808 49776 2864 49832
rect 2932 49776 2988 49832
rect 3056 49776 3112 49832
rect 3180 49776 3236 49832
rect 3304 49776 3360 49832
rect 3428 49776 3484 49832
rect 3552 49776 3608 49832
rect 3676 49776 3732 49832
rect 3800 49776 3856 49832
rect 3924 49776 3980 49832
rect 4048 49776 4104 49832
rect 4172 49776 4228 49832
rect 4296 49776 4352 49832
rect 4420 49776 4476 49832
rect 4544 49776 4600 49832
rect 4668 49776 4724 49832
rect 2808 49652 2864 49708
rect 2932 49652 2988 49708
rect 3056 49652 3112 49708
rect 3180 49652 3236 49708
rect 3304 49652 3360 49708
rect 3428 49652 3484 49708
rect 3552 49707 3559 49708
rect 3559 49707 3608 49708
rect 3676 49707 3683 49708
rect 3683 49707 3732 49708
rect 3800 49707 3807 49708
rect 3807 49707 3856 49708
rect 3924 49707 3931 49708
rect 3931 49707 3980 49708
rect 4048 49707 4055 49708
rect 4055 49707 4104 49708
rect 4172 49707 4179 49708
rect 4179 49707 4228 49708
rect 4296 49707 4303 49708
rect 4303 49707 4352 49708
rect 4420 49707 4427 49708
rect 4427 49707 4476 49708
rect 4544 49707 4551 49708
rect 4551 49707 4600 49708
rect 4668 49707 4675 49708
rect 4675 49707 4724 49708
rect 3552 49652 3608 49707
rect 3676 49652 3732 49707
rect 3800 49652 3856 49707
rect 3924 49652 3980 49707
rect 4048 49652 4104 49707
rect 4172 49652 4228 49707
rect 4296 49652 4352 49707
rect 4420 49652 4476 49707
rect 4544 49652 4600 49707
rect 4668 49652 4724 49707
rect 4861 52492 4917 52548
rect 4985 52492 5041 52548
rect 4861 52368 4917 52424
rect 4985 52368 5041 52424
rect 4861 52244 4917 52300
rect 4985 52244 5041 52300
rect 4861 52120 4917 52176
rect 4985 52120 5041 52176
rect 4861 52017 4917 52052
rect 4861 51996 4863 52017
rect 4863 51996 4915 52017
rect 4915 51996 4917 52017
rect 4985 52017 5041 52052
rect 4985 51996 4987 52017
rect 4987 51996 5039 52017
rect 5039 51996 5041 52017
rect 4861 51893 4917 51928
rect 4861 51872 4863 51893
rect 4863 51872 4915 51893
rect 4915 51872 4917 51893
rect 4985 51893 5041 51928
rect 4985 51872 4987 51893
rect 4987 51872 5039 51893
rect 5039 51872 5041 51893
rect 4861 51748 4917 51804
rect 4985 51748 5041 51804
rect 4861 51624 4917 51680
rect 4985 51624 5041 51680
rect 4861 51500 4917 51556
rect 4985 51500 5041 51556
rect 4861 51376 4917 51432
rect 4985 51376 5041 51432
rect 4861 51252 4917 51308
rect 4985 51252 5041 51308
rect 5178 50892 5234 50948
rect 5302 50892 5358 50948
rect 5426 50892 5482 50948
rect 5550 50892 5606 50948
rect 5674 50892 5730 50948
rect 5798 50892 5854 50948
rect 5922 50892 5978 50948
rect 6046 50892 6102 50948
rect 6170 50892 6226 50948
rect 6294 50892 6350 50948
rect 6418 50892 6474 50948
rect 6542 50892 6598 50948
rect 6666 50892 6722 50948
rect 6790 50892 6846 50948
rect 6914 50892 6970 50948
rect 7038 50892 7094 50948
rect 5178 50768 5234 50824
rect 5302 50768 5358 50824
rect 5426 50768 5482 50824
rect 5550 50768 5606 50824
rect 5674 50768 5730 50824
rect 5798 50768 5854 50824
rect 5922 50768 5978 50824
rect 6046 50768 6102 50824
rect 6170 50768 6226 50824
rect 6294 50768 6350 50824
rect 6418 50768 6474 50824
rect 6542 50768 6598 50824
rect 6666 50768 6722 50824
rect 6790 50768 6846 50824
rect 6914 50768 6970 50824
rect 7038 50768 7094 50824
rect 5178 50693 5234 50700
rect 5178 50644 5180 50693
rect 5180 50644 5232 50693
rect 5232 50644 5234 50693
rect 5302 50693 5358 50700
rect 5302 50644 5304 50693
rect 5304 50644 5356 50693
rect 5356 50644 5358 50693
rect 5426 50693 5482 50700
rect 5426 50644 5428 50693
rect 5428 50644 5480 50693
rect 5480 50644 5482 50693
rect 5550 50693 5606 50700
rect 5550 50644 5552 50693
rect 5552 50644 5604 50693
rect 5604 50644 5606 50693
rect 5674 50693 5730 50700
rect 5674 50644 5676 50693
rect 5676 50644 5728 50693
rect 5728 50644 5730 50693
rect 5798 50693 5854 50700
rect 5798 50644 5800 50693
rect 5800 50644 5852 50693
rect 5852 50644 5854 50693
rect 5922 50693 5978 50700
rect 5922 50644 5924 50693
rect 5924 50644 5976 50693
rect 5976 50644 5978 50693
rect 6046 50693 6102 50700
rect 6046 50644 6048 50693
rect 6048 50644 6100 50693
rect 6100 50644 6102 50693
rect 6170 50693 6226 50700
rect 6170 50644 6172 50693
rect 6172 50644 6224 50693
rect 6224 50644 6226 50693
rect 6294 50693 6350 50700
rect 6294 50644 6296 50693
rect 6296 50644 6348 50693
rect 6348 50644 6350 50693
rect 6418 50693 6474 50700
rect 6418 50644 6420 50693
rect 6420 50644 6472 50693
rect 6472 50644 6474 50693
rect 6542 50693 6598 50700
rect 6542 50644 6544 50693
rect 6544 50644 6596 50693
rect 6596 50644 6598 50693
rect 6666 50693 6722 50700
rect 6666 50644 6668 50693
rect 6668 50644 6720 50693
rect 6720 50644 6722 50693
rect 6790 50693 6846 50700
rect 6790 50644 6792 50693
rect 6792 50644 6844 50693
rect 6844 50644 6846 50693
rect 6914 50693 6970 50700
rect 6914 50644 6916 50693
rect 6916 50644 6968 50693
rect 6968 50644 6970 50693
rect 7038 50693 7094 50700
rect 7038 50644 7040 50693
rect 7040 50644 7092 50693
rect 7092 50644 7094 50693
rect 5178 50569 5234 50576
rect 5178 50520 5180 50569
rect 5180 50520 5232 50569
rect 5232 50520 5234 50569
rect 5302 50569 5358 50576
rect 5302 50520 5304 50569
rect 5304 50520 5356 50569
rect 5356 50520 5358 50569
rect 5426 50569 5482 50576
rect 5426 50520 5428 50569
rect 5428 50520 5480 50569
rect 5480 50520 5482 50569
rect 5550 50569 5606 50576
rect 5550 50520 5552 50569
rect 5552 50520 5604 50569
rect 5604 50520 5606 50569
rect 5674 50569 5730 50576
rect 5674 50520 5676 50569
rect 5676 50520 5728 50569
rect 5728 50520 5730 50569
rect 5798 50569 5854 50576
rect 5798 50520 5800 50569
rect 5800 50520 5852 50569
rect 5852 50520 5854 50569
rect 5922 50569 5978 50576
rect 5922 50520 5924 50569
rect 5924 50520 5976 50569
rect 5976 50520 5978 50569
rect 6046 50569 6102 50576
rect 6046 50520 6048 50569
rect 6048 50520 6100 50569
rect 6100 50520 6102 50569
rect 6170 50569 6226 50576
rect 6170 50520 6172 50569
rect 6172 50520 6224 50569
rect 6224 50520 6226 50569
rect 6294 50569 6350 50576
rect 6294 50520 6296 50569
rect 6296 50520 6348 50569
rect 6348 50520 6350 50569
rect 6418 50569 6474 50576
rect 6418 50520 6420 50569
rect 6420 50520 6472 50569
rect 6472 50520 6474 50569
rect 6542 50569 6598 50576
rect 6542 50520 6544 50569
rect 6544 50520 6596 50569
rect 6596 50520 6598 50569
rect 6666 50569 6722 50576
rect 6666 50520 6668 50569
rect 6668 50520 6720 50569
rect 6720 50520 6722 50569
rect 6790 50569 6846 50576
rect 6790 50520 6792 50569
rect 6792 50520 6844 50569
rect 6844 50520 6846 50569
rect 6914 50569 6970 50576
rect 6914 50520 6916 50569
rect 6916 50520 6968 50569
rect 6968 50520 6970 50569
rect 7038 50569 7094 50576
rect 7038 50520 7040 50569
rect 7040 50520 7092 50569
rect 7092 50520 7094 50569
rect 5178 50396 5234 50452
rect 5302 50396 5358 50452
rect 5426 50396 5482 50452
rect 5550 50396 5606 50452
rect 5674 50396 5730 50452
rect 5798 50396 5854 50452
rect 5922 50396 5978 50452
rect 6046 50396 6102 50452
rect 6170 50396 6226 50452
rect 6294 50396 6350 50452
rect 6418 50396 6474 50452
rect 6542 50396 6598 50452
rect 6666 50396 6722 50452
rect 6790 50396 6846 50452
rect 6914 50396 6970 50452
rect 7038 50396 7094 50452
rect 5178 50272 5234 50328
rect 5302 50272 5358 50328
rect 5426 50272 5482 50328
rect 5550 50272 5606 50328
rect 5674 50272 5730 50328
rect 5798 50272 5854 50328
rect 5922 50272 5978 50328
rect 6046 50272 6102 50328
rect 6170 50272 6226 50328
rect 6294 50272 6350 50328
rect 6418 50272 6474 50328
rect 6542 50272 6598 50328
rect 6666 50272 6722 50328
rect 6790 50272 6846 50328
rect 6914 50272 6970 50328
rect 7038 50272 7094 50328
rect 5178 50148 5234 50204
rect 5302 50148 5358 50204
rect 5426 50148 5482 50204
rect 5550 50148 5606 50204
rect 5674 50148 5730 50204
rect 5798 50148 5854 50204
rect 5922 50148 5978 50204
rect 6046 50148 6102 50204
rect 6170 50148 6226 50204
rect 6294 50148 6350 50204
rect 6418 50148 6474 50204
rect 6542 50148 6598 50204
rect 6666 50148 6722 50204
rect 6790 50148 6846 50204
rect 6914 50148 6970 50204
rect 7038 50148 7094 50204
rect 5178 50024 5234 50080
rect 5302 50024 5358 50080
rect 5426 50024 5482 50080
rect 5550 50024 5606 50080
rect 5674 50024 5730 50080
rect 5798 50024 5854 50080
rect 5922 50024 5978 50080
rect 6046 50024 6102 50080
rect 6170 50024 6226 50080
rect 6294 50024 6350 50080
rect 6418 50024 6474 50080
rect 6542 50024 6598 50080
rect 6666 50024 6722 50080
rect 6790 50024 6846 50080
rect 6914 50024 6970 50080
rect 7038 50024 7094 50080
rect 5178 49900 5234 49956
rect 5302 49900 5358 49956
rect 5426 49900 5482 49956
rect 5550 49900 5606 49956
rect 5674 49900 5730 49956
rect 5798 49900 5854 49956
rect 5922 49900 5978 49956
rect 6046 49900 6102 49956
rect 6170 49900 6226 49956
rect 6294 49900 6350 49956
rect 6418 49900 6474 49956
rect 6542 49900 6598 49956
rect 6666 49900 6722 49956
rect 6790 49900 6846 49956
rect 6914 49900 6970 49956
rect 7038 49900 7094 49956
rect 5178 49776 5234 49832
rect 5302 49776 5358 49832
rect 5426 49776 5482 49832
rect 5550 49776 5606 49832
rect 5674 49776 5730 49832
rect 5798 49776 5854 49832
rect 5922 49776 5978 49832
rect 6046 49776 6102 49832
rect 6170 49776 6226 49832
rect 6294 49776 6350 49832
rect 6418 49776 6474 49832
rect 6542 49776 6598 49832
rect 6666 49776 6722 49832
rect 6790 49776 6846 49832
rect 6914 49776 6970 49832
rect 7038 49776 7094 49832
rect 5178 49707 5180 49708
rect 5180 49707 5232 49708
rect 5232 49707 5234 49708
rect 5178 49652 5234 49707
rect 5302 49707 5304 49708
rect 5304 49707 5356 49708
rect 5356 49707 5358 49708
rect 5302 49652 5358 49707
rect 5426 49707 5428 49708
rect 5428 49707 5480 49708
rect 5480 49707 5482 49708
rect 5426 49652 5482 49707
rect 5550 49707 5552 49708
rect 5552 49707 5604 49708
rect 5604 49707 5606 49708
rect 5550 49652 5606 49707
rect 5674 49707 5676 49708
rect 5676 49707 5728 49708
rect 5728 49707 5730 49708
rect 5674 49652 5730 49707
rect 5798 49707 5800 49708
rect 5800 49707 5852 49708
rect 5852 49707 5854 49708
rect 5798 49652 5854 49707
rect 5922 49707 5924 49708
rect 5924 49707 5976 49708
rect 5976 49707 5978 49708
rect 5922 49652 5978 49707
rect 6046 49707 6048 49708
rect 6048 49707 6100 49708
rect 6100 49707 6102 49708
rect 6046 49652 6102 49707
rect 6170 49707 6172 49708
rect 6172 49707 6224 49708
rect 6224 49707 6226 49708
rect 6170 49652 6226 49707
rect 6294 49707 6296 49708
rect 6296 49707 6348 49708
rect 6348 49707 6350 49708
rect 6294 49652 6350 49707
rect 6418 49707 6420 49708
rect 6420 49707 6472 49708
rect 6472 49707 6474 49708
rect 6418 49652 6474 49707
rect 6542 49707 6544 49708
rect 6544 49707 6596 49708
rect 6596 49707 6598 49708
rect 6542 49652 6598 49707
rect 6666 49707 6668 49708
rect 6668 49707 6720 49708
rect 6720 49707 6722 49708
rect 6666 49652 6722 49707
rect 6790 49707 6792 49708
rect 6792 49707 6844 49708
rect 6844 49707 6846 49708
rect 6790 49652 6846 49707
rect 6914 49707 6916 49708
rect 6916 49707 6968 49708
rect 6968 49707 6970 49708
rect 6914 49652 6970 49707
rect 7038 49707 7040 49708
rect 7040 49707 7092 49708
rect 7092 49707 7094 49708
rect 7038 49652 7094 49707
rect 7275 52492 7331 52548
rect 7399 52492 7455 52548
rect 7523 52492 7579 52548
rect 7647 52492 7703 52548
rect 7275 52368 7331 52424
rect 7399 52368 7455 52424
rect 7523 52368 7579 52424
rect 7647 52368 7703 52424
rect 7275 52244 7331 52300
rect 7399 52244 7455 52300
rect 7523 52244 7579 52300
rect 7647 52244 7703 52300
rect 7275 52120 7331 52176
rect 7399 52120 7455 52176
rect 7523 52120 7579 52176
rect 7647 52120 7703 52176
rect 7275 52017 7331 52052
rect 7275 51996 7277 52017
rect 7277 51996 7329 52017
rect 7329 51996 7331 52017
rect 7399 52017 7455 52052
rect 7399 51996 7401 52017
rect 7401 51996 7453 52017
rect 7453 51996 7455 52017
rect 7523 52017 7579 52052
rect 7523 51996 7525 52017
rect 7525 51996 7577 52017
rect 7577 51996 7579 52017
rect 7647 52017 7703 52052
rect 7647 51996 7649 52017
rect 7649 51996 7701 52017
rect 7701 51996 7703 52017
rect 7275 51893 7331 51928
rect 7275 51872 7277 51893
rect 7277 51872 7329 51893
rect 7329 51872 7331 51893
rect 7399 51893 7455 51928
rect 7399 51872 7401 51893
rect 7401 51872 7453 51893
rect 7453 51872 7455 51893
rect 7523 51893 7579 51928
rect 7523 51872 7525 51893
rect 7525 51872 7577 51893
rect 7577 51872 7579 51893
rect 7647 51893 7703 51928
rect 7647 51872 7649 51893
rect 7649 51872 7701 51893
rect 7701 51872 7703 51893
rect 7275 51748 7331 51804
rect 7399 51748 7455 51804
rect 7523 51748 7579 51804
rect 7647 51748 7703 51804
rect 7275 51624 7331 51680
rect 7399 51624 7455 51680
rect 7523 51624 7579 51680
rect 7647 51624 7703 51680
rect 7275 51500 7331 51556
rect 7399 51500 7455 51556
rect 7523 51500 7579 51556
rect 7647 51500 7703 51556
rect 7275 51376 7331 51432
rect 7399 51376 7455 51432
rect 7523 51376 7579 51432
rect 7647 51376 7703 51432
rect 7275 51252 7331 51308
rect 7399 51252 7455 51308
rect 7523 51252 7579 51308
rect 7647 51252 7703 51308
rect 7884 50892 7940 50948
rect 8008 50892 8064 50948
rect 8132 50892 8188 50948
rect 8256 50892 8312 50948
rect 8380 50892 8436 50948
rect 8504 50892 8560 50948
rect 8628 50892 8684 50948
rect 8752 50892 8808 50948
rect 8876 50892 8932 50948
rect 9000 50892 9056 50948
rect 9124 50892 9180 50948
rect 9248 50892 9304 50948
rect 9372 50892 9428 50948
rect 9496 50892 9552 50948
rect 9620 50892 9676 50948
rect 9744 50892 9800 50948
rect 7884 50768 7940 50824
rect 8008 50768 8064 50824
rect 8132 50768 8188 50824
rect 8256 50768 8312 50824
rect 8380 50768 8436 50824
rect 8504 50768 8560 50824
rect 8628 50768 8684 50824
rect 8752 50768 8808 50824
rect 8876 50768 8932 50824
rect 9000 50768 9056 50824
rect 9124 50768 9180 50824
rect 9248 50768 9304 50824
rect 9372 50768 9428 50824
rect 9496 50768 9552 50824
rect 9620 50768 9676 50824
rect 9744 50768 9800 50824
rect 7884 50693 7940 50700
rect 7884 50644 7886 50693
rect 7886 50644 7938 50693
rect 7938 50644 7940 50693
rect 8008 50693 8064 50700
rect 8008 50644 8010 50693
rect 8010 50644 8062 50693
rect 8062 50644 8064 50693
rect 8132 50693 8188 50700
rect 8132 50644 8134 50693
rect 8134 50644 8186 50693
rect 8186 50644 8188 50693
rect 8256 50693 8312 50700
rect 8256 50644 8258 50693
rect 8258 50644 8310 50693
rect 8310 50644 8312 50693
rect 8380 50693 8436 50700
rect 8380 50644 8382 50693
rect 8382 50644 8434 50693
rect 8434 50644 8436 50693
rect 8504 50693 8560 50700
rect 8504 50644 8506 50693
rect 8506 50644 8558 50693
rect 8558 50644 8560 50693
rect 8628 50693 8684 50700
rect 8628 50644 8630 50693
rect 8630 50644 8682 50693
rect 8682 50644 8684 50693
rect 8752 50693 8808 50700
rect 8752 50644 8754 50693
rect 8754 50644 8806 50693
rect 8806 50644 8808 50693
rect 8876 50693 8932 50700
rect 8876 50644 8878 50693
rect 8878 50644 8930 50693
rect 8930 50644 8932 50693
rect 9000 50693 9056 50700
rect 9000 50644 9002 50693
rect 9002 50644 9054 50693
rect 9054 50644 9056 50693
rect 9124 50693 9180 50700
rect 9124 50644 9126 50693
rect 9126 50644 9178 50693
rect 9178 50644 9180 50693
rect 9248 50693 9304 50700
rect 9248 50644 9250 50693
rect 9250 50644 9302 50693
rect 9302 50644 9304 50693
rect 9372 50693 9428 50700
rect 9372 50644 9374 50693
rect 9374 50644 9426 50693
rect 9426 50644 9428 50693
rect 9496 50693 9552 50700
rect 9496 50644 9498 50693
rect 9498 50644 9550 50693
rect 9550 50644 9552 50693
rect 9620 50693 9676 50700
rect 9620 50644 9622 50693
rect 9622 50644 9674 50693
rect 9674 50644 9676 50693
rect 9744 50693 9800 50700
rect 9744 50644 9746 50693
rect 9746 50644 9798 50693
rect 9798 50644 9800 50693
rect 7884 50569 7940 50576
rect 7884 50520 7886 50569
rect 7886 50520 7938 50569
rect 7938 50520 7940 50569
rect 8008 50569 8064 50576
rect 8008 50520 8010 50569
rect 8010 50520 8062 50569
rect 8062 50520 8064 50569
rect 8132 50569 8188 50576
rect 8132 50520 8134 50569
rect 8134 50520 8186 50569
rect 8186 50520 8188 50569
rect 8256 50569 8312 50576
rect 8256 50520 8258 50569
rect 8258 50520 8310 50569
rect 8310 50520 8312 50569
rect 8380 50569 8436 50576
rect 8380 50520 8382 50569
rect 8382 50520 8434 50569
rect 8434 50520 8436 50569
rect 8504 50569 8560 50576
rect 8504 50520 8506 50569
rect 8506 50520 8558 50569
rect 8558 50520 8560 50569
rect 8628 50569 8684 50576
rect 8628 50520 8630 50569
rect 8630 50520 8682 50569
rect 8682 50520 8684 50569
rect 8752 50569 8808 50576
rect 8752 50520 8754 50569
rect 8754 50520 8806 50569
rect 8806 50520 8808 50569
rect 8876 50569 8932 50576
rect 8876 50520 8878 50569
rect 8878 50520 8930 50569
rect 8930 50520 8932 50569
rect 9000 50569 9056 50576
rect 9000 50520 9002 50569
rect 9002 50520 9054 50569
rect 9054 50520 9056 50569
rect 9124 50569 9180 50576
rect 9124 50520 9126 50569
rect 9126 50520 9178 50569
rect 9178 50520 9180 50569
rect 9248 50569 9304 50576
rect 9248 50520 9250 50569
rect 9250 50520 9302 50569
rect 9302 50520 9304 50569
rect 9372 50569 9428 50576
rect 9372 50520 9374 50569
rect 9374 50520 9426 50569
rect 9426 50520 9428 50569
rect 9496 50569 9552 50576
rect 9496 50520 9498 50569
rect 9498 50520 9550 50569
rect 9550 50520 9552 50569
rect 9620 50569 9676 50576
rect 9620 50520 9622 50569
rect 9622 50520 9674 50569
rect 9674 50520 9676 50569
rect 9744 50569 9800 50576
rect 9744 50520 9746 50569
rect 9746 50520 9798 50569
rect 9798 50520 9800 50569
rect 7884 50396 7940 50452
rect 8008 50396 8064 50452
rect 8132 50396 8188 50452
rect 8256 50396 8312 50452
rect 8380 50396 8436 50452
rect 8504 50396 8560 50452
rect 8628 50396 8684 50452
rect 8752 50396 8808 50452
rect 8876 50396 8932 50452
rect 9000 50396 9056 50452
rect 9124 50396 9180 50452
rect 9248 50396 9304 50452
rect 9372 50396 9428 50452
rect 9496 50396 9552 50452
rect 9620 50396 9676 50452
rect 9744 50396 9800 50452
rect 7884 50272 7940 50328
rect 8008 50272 8064 50328
rect 8132 50272 8188 50328
rect 8256 50272 8312 50328
rect 8380 50272 8436 50328
rect 8504 50272 8560 50328
rect 8628 50272 8684 50328
rect 8752 50272 8808 50328
rect 8876 50272 8932 50328
rect 9000 50272 9056 50328
rect 9124 50272 9180 50328
rect 9248 50272 9304 50328
rect 9372 50272 9428 50328
rect 9496 50272 9552 50328
rect 9620 50272 9676 50328
rect 9744 50272 9800 50328
rect 7884 50148 7940 50204
rect 8008 50148 8064 50204
rect 8132 50148 8188 50204
rect 8256 50148 8312 50204
rect 8380 50148 8436 50204
rect 8504 50148 8560 50204
rect 8628 50148 8684 50204
rect 8752 50148 8808 50204
rect 8876 50148 8932 50204
rect 9000 50148 9056 50204
rect 9124 50148 9180 50204
rect 9248 50148 9304 50204
rect 9372 50148 9428 50204
rect 9496 50148 9552 50204
rect 9620 50148 9676 50204
rect 9744 50148 9800 50204
rect 7884 50024 7940 50080
rect 8008 50024 8064 50080
rect 8132 50024 8188 50080
rect 8256 50024 8312 50080
rect 8380 50024 8436 50080
rect 8504 50024 8560 50080
rect 8628 50024 8684 50080
rect 8752 50024 8808 50080
rect 8876 50024 8932 50080
rect 9000 50024 9056 50080
rect 9124 50024 9180 50080
rect 9248 50024 9304 50080
rect 9372 50024 9428 50080
rect 9496 50024 9552 50080
rect 9620 50024 9676 50080
rect 9744 50024 9800 50080
rect 7884 49900 7940 49956
rect 8008 49900 8064 49956
rect 8132 49900 8188 49956
rect 8256 49900 8312 49956
rect 8380 49900 8436 49956
rect 8504 49900 8560 49956
rect 8628 49900 8684 49956
rect 8752 49900 8808 49956
rect 8876 49900 8932 49956
rect 9000 49900 9056 49956
rect 9124 49900 9180 49956
rect 9248 49900 9304 49956
rect 9372 49900 9428 49956
rect 9496 49900 9552 49956
rect 9620 49900 9676 49956
rect 9744 49900 9800 49956
rect 7884 49776 7940 49832
rect 8008 49776 8064 49832
rect 8132 49776 8188 49832
rect 8256 49776 8312 49832
rect 8380 49776 8436 49832
rect 8504 49776 8560 49832
rect 8628 49776 8684 49832
rect 8752 49776 8808 49832
rect 8876 49776 8932 49832
rect 9000 49776 9056 49832
rect 9124 49776 9180 49832
rect 9248 49776 9304 49832
rect 9372 49776 9428 49832
rect 9496 49776 9552 49832
rect 9620 49776 9676 49832
rect 9744 49776 9800 49832
rect 7884 49707 7886 49708
rect 7886 49707 7938 49708
rect 7938 49707 7940 49708
rect 7884 49652 7940 49707
rect 8008 49707 8010 49708
rect 8010 49707 8062 49708
rect 8062 49707 8064 49708
rect 8008 49652 8064 49707
rect 8132 49707 8134 49708
rect 8134 49707 8186 49708
rect 8186 49707 8188 49708
rect 8132 49652 8188 49707
rect 8256 49707 8258 49708
rect 8258 49707 8310 49708
rect 8310 49707 8312 49708
rect 8256 49652 8312 49707
rect 8380 49707 8382 49708
rect 8382 49707 8434 49708
rect 8434 49707 8436 49708
rect 8380 49652 8436 49707
rect 8504 49707 8506 49708
rect 8506 49707 8558 49708
rect 8558 49707 8560 49708
rect 8504 49652 8560 49707
rect 8628 49707 8630 49708
rect 8630 49707 8682 49708
rect 8682 49707 8684 49708
rect 8628 49652 8684 49707
rect 8752 49707 8754 49708
rect 8754 49707 8806 49708
rect 8806 49707 8808 49708
rect 8752 49652 8808 49707
rect 8876 49707 8878 49708
rect 8878 49707 8930 49708
rect 8930 49707 8932 49708
rect 8876 49652 8932 49707
rect 9000 49707 9002 49708
rect 9002 49707 9054 49708
rect 9054 49707 9056 49708
rect 9000 49652 9056 49707
rect 9124 49707 9126 49708
rect 9126 49707 9178 49708
rect 9178 49707 9180 49708
rect 9124 49652 9180 49707
rect 9248 49707 9250 49708
rect 9250 49707 9302 49708
rect 9302 49707 9304 49708
rect 9248 49652 9304 49707
rect 9372 49707 9374 49708
rect 9374 49707 9426 49708
rect 9426 49707 9428 49708
rect 9372 49652 9428 49707
rect 9496 49707 9498 49708
rect 9498 49707 9550 49708
rect 9550 49707 9552 49708
rect 9496 49652 9552 49707
rect 9620 49707 9622 49708
rect 9622 49707 9674 49708
rect 9674 49707 9676 49708
rect 9620 49652 9676 49707
rect 9744 49707 9746 49708
rect 9746 49707 9798 49708
rect 9798 49707 9800 49708
rect 9744 49652 9800 49707
rect 9937 52492 9993 52548
rect 10061 52492 10117 52548
rect 9937 52368 9993 52424
rect 10061 52368 10117 52424
rect 9937 52244 9993 52300
rect 10061 52244 10117 52300
rect 9937 52120 9993 52176
rect 10061 52120 10117 52176
rect 9937 52017 9993 52052
rect 9937 51996 9939 52017
rect 9939 51996 9991 52017
rect 9991 51996 9993 52017
rect 10061 52017 10117 52052
rect 10061 51996 10063 52017
rect 10063 51996 10115 52017
rect 10115 51996 10117 52017
rect 9937 51893 9993 51928
rect 9937 51872 9939 51893
rect 9939 51872 9991 51893
rect 9991 51872 9993 51893
rect 10061 51893 10117 51928
rect 10061 51872 10063 51893
rect 10063 51872 10115 51893
rect 10115 51872 10117 51893
rect 9937 51748 9993 51804
rect 10061 51748 10117 51804
rect 9937 51624 9993 51680
rect 10061 51624 10117 51680
rect 9937 51500 9993 51556
rect 10061 51500 10117 51556
rect 9937 51376 9993 51432
rect 10061 51376 10117 51432
rect 9937 51252 9993 51308
rect 10061 51252 10117 51308
rect 10254 50892 10310 50948
rect 10378 50892 10434 50948
rect 10502 50892 10558 50948
rect 10626 50892 10682 50948
rect 10750 50892 10806 50948
rect 10874 50892 10930 50948
rect 10998 50892 11054 50948
rect 11122 50892 11178 50948
rect 11246 50892 11302 50948
rect 11370 50892 11426 50948
rect 11494 50892 11550 50948
rect 11618 50892 11674 50948
rect 11742 50892 11798 50948
rect 11866 50892 11922 50948
rect 11990 50892 12046 50948
rect 12114 50892 12170 50948
rect 10254 50768 10310 50824
rect 10378 50768 10434 50824
rect 10502 50768 10558 50824
rect 10626 50768 10682 50824
rect 10750 50768 10806 50824
rect 10874 50768 10930 50824
rect 10998 50768 11054 50824
rect 11122 50768 11178 50824
rect 11246 50768 11302 50824
rect 11370 50768 11426 50824
rect 11494 50768 11550 50824
rect 11618 50768 11674 50824
rect 11742 50768 11798 50824
rect 11866 50768 11922 50824
rect 11990 50768 12046 50824
rect 12114 50768 12170 50824
rect 10254 50693 10310 50700
rect 10378 50693 10434 50700
rect 10502 50693 10558 50700
rect 10626 50693 10682 50700
rect 10750 50693 10806 50700
rect 10874 50693 10930 50700
rect 10998 50693 11054 50700
rect 11122 50693 11178 50700
rect 11246 50693 11302 50700
rect 11370 50693 11426 50700
rect 10254 50644 10303 50693
rect 10303 50644 10310 50693
rect 10378 50644 10427 50693
rect 10427 50644 10434 50693
rect 10502 50644 10551 50693
rect 10551 50644 10558 50693
rect 10626 50644 10675 50693
rect 10675 50644 10682 50693
rect 10750 50644 10799 50693
rect 10799 50644 10806 50693
rect 10874 50644 10923 50693
rect 10923 50644 10930 50693
rect 10998 50644 11047 50693
rect 11047 50644 11054 50693
rect 11122 50644 11171 50693
rect 11171 50644 11178 50693
rect 11246 50644 11295 50693
rect 11295 50644 11302 50693
rect 11370 50644 11419 50693
rect 11419 50644 11426 50693
rect 11494 50644 11550 50700
rect 11618 50644 11674 50700
rect 11742 50644 11798 50700
rect 11866 50644 11922 50700
rect 11990 50644 12046 50700
rect 12114 50644 12170 50700
rect 10254 50569 10310 50576
rect 10378 50569 10434 50576
rect 10502 50569 10558 50576
rect 10626 50569 10682 50576
rect 10750 50569 10806 50576
rect 10874 50569 10930 50576
rect 10998 50569 11054 50576
rect 11122 50569 11178 50576
rect 11246 50569 11302 50576
rect 11370 50569 11426 50576
rect 10254 50520 10303 50569
rect 10303 50520 10310 50569
rect 10378 50520 10427 50569
rect 10427 50520 10434 50569
rect 10502 50520 10551 50569
rect 10551 50520 10558 50569
rect 10626 50520 10675 50569
rect 10675 50520 10682 50569
rect 10750 50520 10799 50569
rect 10799 50520 10806 50569
rect 10874 50520 10923 50569
rect 10923 50520 10930 50569
rect 10998 50520 11047 50569
rect 11047 50520 11054 50569
rect 11122 50520 11171 50569
rect 11171 50520 11178 50569
rect 11246 50520 11295 50569
rect 11295 50520 11302 50569
rect 11370 50520 11419 50569
rect 11419 50520 11426 50569
rect 11494 50520 11550 50576
rect 11618 50520 11674 50576
rect 11742 50520 11798 50576
rect 11866 50520 11922 50576
rect 11990 50520 12046 50576
rect 12114 50520 12170 50576
rect 10254 50396 10310 50452
rect 10378 50396 10434 50452
rect 10502 50396 10558 50452
rect 10626 50396 10682 50452
rect 10750 50396 10806 50452
rect 10874 50396 10930 50452
rect 10998 50396 11054 50452
rect 11122 50396 11178 50452
rect 11246 50396 11302 50452
rect 11370 50396 11426 50452
rect 11494 50396 11550 50452
rect 11618 50396 11674 50452
rect 11742 50396 11798 50452
rect 11866 50396 11922 50452
rect 11990 50396 12046 50452
rect 12114 50396 12170 50452
rect 10254 50272 10310 50328
rect 10378 50272 10434 50328
rect 10502 50272 10558 50328
rect 10626 50272 10682 50328
rect 10750 50272 10806 50328
rect 10874 50272 10930 50328
rect 10998 50272 11054 50328
rect 11122 50272 11178 50328
rect 11246 50272 11302 50328
rect 11370 50272 11426 50328
rect 11494 50272 11550 50328
rect 11618 50272 11674 50328
rect 11742 50272 11798 50328
rect 11866 50272 11922 50328
rect 11990 50272 12046 50328
rect 12114 50272 12170 50328
rect 10254 50148 10310 50204
rect 10378 50148 10434 50204
rect 10502 50148 10558 50204
rect 10626 50148 10682 50204
rect 10750 50148 10806 50204
rect 10874 50148 10930 50204
rect 10998 50148 11054 50204
rect 11122 50148 11178 50204
rect 11246 50148 11302 50204
rect 11370 50148 11426 50204
rect 11494 50148 11550 50204
rect 11618 50148 11674 50204
rect 11742 50148 11798 50204
rect 11866 50148 11922 50204
rect 11990 50148 12046 50204
rect 12114 50148 12170 50204
rect 10254 50024 10310 50080
rect 10378 50024 10434 50080
rect 10502 50024 10558 50080
rect 10626 50024 10682 50080
rect 10750 50024 10806 50080
rect 10874 50024 10930 50080
rect 10998 50024 11054 50080
rect 11122 50024 11178 50080
rect 11246 50024 11302 50080
rect 11370 50024 11426 50080
rect 11494 50024 11550 50080
rect 11618 50024 11674 50080
rect 11742 50024 11798 50080
rect 11866 50024 11922 50080
rect 11990 50024 12046 50080
rect 12114 50024 12170 50080
rect 10254 49900 10310 49956
rect 10378 49900 10434 49956
rect 10502 49900 10558 49956
rect 10626 49900 10682 49956
rect 10750 49900 10806 49956
rect 10874 49900 10930 49956
rect 10998 49900 11054 49956
rect 11122 49900 11178 49956
rect 11246 49900 11302 49956
rect 11370 49900 11426 49956
rect 11494 49900 11550 49956
rect 11618 49900 11674 49956
rect 11742 49900 11798 49956
rect 11866 49900 11922 49956
rect 11990 49900 12046 49956
rect 12114 49900 12170 49956
rect 10254 49776 10310 49832
rect 10378 49776 10434 49832
rect 10502 49776 10558 49832
rect 10626 49776 10682 49832
rect 10750 49776 10806 49832
rect 10874 49776 10930 49832
rect 10998 49776 11054 49832
rect 11122 49776 11178 49832
rect 11246 49776 11302 49832
rect 11370 49776 11426 49832
rect 11494 49776 11550 49832
rect 11618 49776 11674 49832
rect 11742 49776 11798 49832
rect 11866 49776 11922 49832
rect 11990 49776 12046 49832
rect 12114 49776 12170 49832
rect 10254 49707 10303 49708
rect 10303 49707 10310 49708
rect 10378 49707 10427 49708
rect 10427 49707 10434 49708
rect 10502 49707 10551 49708
rect 10551 49707 10558 49708
rect 10626 49707 10675 49708
rect 10675 49707 10682 49708
rect 10750 49707 10799 49708
rect 10799 49707 10806 49708
rect 10874 49707 10923 49708
rect 10923 49707 10930 49708
rect 10998 49707 11047 49708
rect 11047 49707 11054 49708
rect 11122 49707 11171 49708
rect 11171 49707 11178 49708
rect 11246 49707 11295 49708
rect 11295 49707 11302 49708
rect 11370 49707 11419 49708
rect 11419 49707 11426 49708
rect 10254 49652 10310 49707
rect 10378 49652 10434 49707
rect 10502 49652 10558 49707
rect 10626 49652 10682 49707
rect 10750 49652 10806 49707
rect 10874 49652 10930 49707
rect 10998 49652 11054 49707
rect 11122 49652 11178 49707
rect 11246 49652 11302 49707
rect 11370 49652 11426 49707
rect 11494 49652 11550 49708
rect 11618 49652 11674 49708
rect 11742 49652 11798 49708
rect 11866 49652 11922 49708
rect 11990 49652 12046 49708
rect 12114 49652 12170 49708
rect 12307 52492 12363 52548
rect 12431 52492 12487 52548
rect 12307 52368 12363 52424
rect 12431 52368 12487 52424
rect 12307 52244 12363 52300
rect 12431 52244 12487 52300
rect 12307 52120 12363 52176
rect 12431 52120 12487 52176
rect 12307 51996 12363 52052
rect 12431 51996 12487 52052
rect 12307 51872 12363 51928
rect 12431 51872 12487 51928
rect 12307 51748 12363 51804
rect 12431 51748 12487 51804
rect 12307 51624 12363 51680
rect 12431 51624 12487 51680
rect 12307 51500 12363 51556
rect 12431 51500 12487 51556
rect 12307 51376 12363 51432
rect 12431 51376 12487 51432
rect 12307 51252 12363 51308
rect 12431 51252 12487 51308
rect 14902 52574 14958 52576
rect 14902 52522 14904 52574
rect 14904 52522 14956 52574
rect 14956 52522 14958 52574
rect 14902 52466 14958 52522
rect 14902 52414 14904 52466
rect 14904 52414 14956 52466
rect 14956 52414 14958 52466
rect 14902 52358 14958 52414
rect 14902 52306 14904 52358
rect 14904 52306 14956 52358
rect 14956 52306 14958 52358
rect 14902 52250 14958 52306
rect 14902 52198 14904 52250
rect 14904 52198 14956 52250
rect 14956 52198 14958 52250
rect 14902 52142 14958 52198
rect 14902 52090 14904 52142
rect 14904 52090 14956 52142
rect 14956 52090 14958 52142
rect 14902 52034 14958 52090
rect 14902 51982 14904 52034
rect 14904 51982 14956 52034
rect 14956 51982 14958 52034
rect 14902 51926 14958 51982
rect 14902 51874 14904 51926
rect 14904 51874 14956 51926
rect 14956 51874 14958 51926
rect 14902 51818 14958 51874
rect 14902 51766 14904 51818
rect 14904 51766 14956 51818
rect 14956 51766 14958 51818
rect 14902 51710 14958 51766
rect 14902 51658 14904 51710
rect 14904 51658 14956 51710
rect 14956 51658 14958 51710
rect 14902 51602 14958 51658
rect 14902 51550 14904 51602
rect 14904 51550 14956 51602
rect 14956 51550 14958 51602
rect 14902 51494 14958 51550
rect 14902 51442 14904 51494
rect 14904 51442 14956 51494
rect 14956 51442 14958 51494
rect 14902 51386 14958 51442
rect 14902 51334 14904 51386
rect 14904 51334 14956 51386
rect 14956 51334 14958 51386
rect 14902 51278 14958 51334
rect 14902 51226 14904 51278
rect 14904 51226 14956 51278
rect 14956 51226 14958 51278
rect 14902 51224 14958 51226
rect 12871 50892 12927 50948
rect 12995 50892 13051 50948
rect 13119 50892 13175 50948
rect 13243 50892 13299 50948
rect 13367 50892 13423 50948
rect 13491 50892 13547 50948
rect 13615 50892 13671 50948
rect 13739 50892 13795 50948
rect 13863 50892 13919 50948
rect 13987 50892 14043 50948
rect 14111 50892 14167 50948
rect 14235 50892 14291 50948
rect 14359 50892 14415 50948
rect 14483 50892 14539 50948
rect 14607 50892 14663 50948
rect 12871 50768 12927 50824
rect 12995 50768 13051 50824
rect 13119 50768 13175 50824
rect 13243 50768 13299 50824
rect 13367 50768 13423 50824
rect 13491 50768 13547 50824
rect 13615 50768 13671 50824
rect 13739 50768 13795 50824
rect 13863 50768 13919 50824
rect 13987 50768 14043 50824
rect 14111 50768 14167 50824
rect 14235 50768 14291 50824
rect 14359 50768 14415 50824
rect 14483 50768 14539 50824
rect 14607 50768 14663 50824
rect 12871 50644 12927 50700
rect 12995 50644 13051 50700
rect 13119 50644 13175 50700
rect 13243 50644 13299 50700
rect 13367 50644 13423 50700
rect 13491 50644 13547 50700
rect 13615 50644 13671 50700
rect 13739 50644 13795 50700
rect 13863 50644 13919 50700
rect 13987 50644 14043 50700
rect 14111 50644 14167 50700
rect 14235 50644 14291 50700
rect 14359 50644 14415 50700
rect 14483 50644 14539 50700
rect 14607 50644 14663 50700
rect 12871 50520 12927 50576
rect 12995 50520 13051 50576
rect 13119 50520 13175 50576
rect 13243 50520 13299 50576
rect 13367 50520 13423 50576
rect 13491 50520 13547 50576
rect 13615 50520 13671 50576
rect 13739 50520 13795 50576
rect 13863 50520 13919 50576
rect 13987 50520 14043 50576
rect 14111 50520 14167 50576
rect 14235 50520 14291 50576
rect 14359 50520 14415 50576
rect 14483 50520 14539 50576
rect 14607 50520 14663 50576
rect 12871 50396 12927 50452
rect 12995 50396 13051 50452
rect 13119 50396 13175 50452
rect 13243 50396 13299 50452
rect 13367 50396 13423 50452
rect 13491 50396 13547 50452
rect 13615 50396 13671 50452
rect 13739 50396 13795 50452
rect 13863 50396 13919 50452
rect 13987 50396 14043 50452
rect 14111 50396 14167 50452
rect 14235 50396 14291 50452
rect 14359 50396 14415 50452
rect 14483 50396 14539 50452
rect 14607 50396 14663 50452
rect 12871 50272 12927 50328
rect 12995 50272 13051 50328
rect 13119 50272 13175 50328
rect 13243 50272 13299 50328
rect 13367 50272 13423 50328
rect 13491 50272 13547 50328
rect 13615 50272 13671 50328
rect 13739 50272 13795 50328
rect 13863 50272 13919 50328
rect 13987 50272 14043 50328
rect 14111 50272 14167 50328
rect 14235 50272 14291 50328
rect 14359 50272 14415 50328
rect 14483 50272 14539 50328
rect 14607 50272 14663 50328
rect 12871 50148 12927 50204
rect 12995 50148 13051 50204
rect 13119 50148 13175 50204
rect 13243 50148 13299 50204
rect 13367 50148 13423 50204
rect 13491 50148 13547 50204
rect 13615 50148 13671 50204
rect 13739 50148 13795 50204
rect 13863 50148 13919 50204
rect 13987 50148 14043 50204
rect 14111 50148 14167 50204
rect 14235 50148 14291 50204
rect 14359 50148 14415 50204
rect 14483 50148 14539 50204
rect 14607 50148 14663 50204
rect 12871 50024 12927 50080
rect 12995 50024 13051 50080
rect 13119 50024 13175 50080
rect 13243 50024 13299 50080
rect 13367 50024 13423 50080
rect 13491 50024 13547 50080
rect 13615 50024 13671 50080
rect 13739 50024 13795 50080
rect 13863 50024 13919 50080
rect 13987 50024 14043 50080
rect 14111 50024 14167 50080
rect 14235 50024 14291 50080
rect 14359 50024 14415 50080
rect 14483 50024 14539 50080
rect 14607 50024 14663 50080
rect 12871 49900 12927 49956
rect 12995 49900 13051 49956
rect 13119 49900 13175 49956
rect 13243 49900 13299 49956
rect 13367 49900 13423 49956
rect 13491 49900 13547 49956
rect 13615 49900 13671 49956
rect 13739 49900 13795 49956
rect 13863 49900 13919 49956
rect 13987 49900 14043 49956
rect 14111 49900 14167 49956
rect 14235 49900 14291 49956
rect 14359 49900 14415 49956
rect 14483 49900 14539 49956
rect 14607 49900 14663 49956
rect 12871 49776 12927 49832
rect 12995 49776 13051 49832
rect 13119 49776 13175 49832
rect 13243 49776 13299 49832
rect 13367 49776 13423 49832
rect 13491 49776 13547 49832
rect 13615 49776 13671 49832
rect 13739 49776 13795 49832
rect 13863 49776 13919 49832
rect 13987 49776 14043 49832
rect 14111 49776 14167 49832
rect 14235 49776 14291 49832
rect 14359 49776 14415 49832
rect 14483 49776 14539 49832
rect 14607 49776 14663 49832
rect 12871 49652 12927 49708
rect 12995 49652 13051 49708
rect 13119 49652 13175 49708
rect 13243 49652 13299 49708
rect 13367 49652 13423 49708
rect 13491 49652 13547 49708
rect 13615 49652 13671 49708
rect 13739 49652 13795 49708
rect 13863 49652 13919 49708
rect 13987 49652 14043 49708
rect 14111 49652 14167 49708
rect 14235 49652 14291 49708
rect 14359 49652 14415 49708
rect 14483 49652 14539 49708
rect 14607 49652 14663 49708
rect 2808 39692 2864 39748
rect 2932 39692 2988 39748
rect 3056 39692 3112 39748
rect 3180 39692 3236 39748
rect 3304 39692 3360 39748
rect 3428 39692 3484 39748
rect 3552 39692 3608 39748
rect 3676 39692 3732 39748
rect 3800 39692 3856 39748
rect 3924 39692 3980 39748
rect 4048 39692 4104 39748
rect 4172 39692 4228 39748
rect 4296 39692 4352 39748
rect 4420 39692 4476 39748
rect 4544 39692 4600 39748
rect 4668 39692 4724 39748
rect 2808 39568 2864 39624
rect 2932 39568 2988 39624
rect 3056 39568 3112 39624
rect 3180 39568 3236 39624
rect 3304 39568 3360 39624
rect 3428 39568 3484 39624
rect 3552 39568 3608 39624
rect 3676 39568 3732 39624
rect 3800 39568 3856 39624
rect 3924 39568 3980 39624
rect 4048 39568 4104 39624
rect 4172 39568 4228 39624
rect 4296 39568 4352 39624
rect 4420 39568 4476 39624
rect 4544 39568 4600 39624
rect 4668 39568 4724 39624
rect 2808 39444 2864 39500
rect 2932 39444 2988 39500
rect 3056 39444 3112 39500
rect 3180 39444 3236 39500
rect 3304 39444 3360 39500
rect 3428 39444 3484 39500
rect 3552 39444 3608 39500
rect 3676 39444 3732 39500
rect 3800 39444 3856 39500
rect 3924 39444 3980 39500
rect 4048 39444 4104 39500
rect 4172 39444 4228 39500
rect 4296 39444 4352 39500
rect 4420 39444 4476 39500
rect 4544 39444 4600 39500
rect 4668 39444 4724 39500
rect 2808 39320 2864 39376
rect 2932 39320 2988 39376
rect 3056 39320 3112 39376
rect 3180 39320 3236 39376
rect 3304 39320 3360 39376
rect 3428 39320 3484 39376
rect 3552 39320 3608 39376
rect 3676 39320 3732 39376
rect 3800 39320 3856 39376
rect 3924 39320 3980 39376
rect 4048 39320 4104 39376
rect 4172 39320 4228 39376
rect 4296 39320 4352 39376
rect 4420 39320 4476 39376
rect 4544 39320 4600 39376
rect 4668 39320 4724 39376
rect 2808 39196 2864 39252
rect 2932 39196 2988 39252
rect 3056 39196 3112 39252
rect 3180 39196 3236 39252
rect 3304 39196 3360 39252
rect 3428 39196 3484 39252
rect 3552 39196 3608 39252
rect 3676 39196 3732 39252
rect 3800 39196 3856 39252
rect 3924 39196 3980 39252
rect 4048 39196 4104 39252
rect 4172 39196 4228 39252
rect 4296 39196 4352 39252
rect 4420 39196 4476 39252
rect 4544 39196 4600 39252
rect 4668 39196 4724 39252
rect 2808 39072 2864 39128
rect 2932 39072 2988 39128
rect 3056 39072 3112 39128
rect 3180 39072 3236 39128
rect 3304 39072 3360 39128
rect 3428 39072 3484 39128
rect 3552 39072 3608 39128
rect 3676 39072 3732 39128
rect 3800 39072 3856 39128
rect 3924 39072 3980 39128
rect 4048 39072 4104 39128
rect 4172 39072 4228 39128
rect 4296 39072 4352 39128
rect 4420 39072 4476 39128
rect 4544 39072 4600 39128
rect 4668 39072 4724 39128
rect 2808 38948 2864 39004
rect 2932 38948 2988 39004
rect 3056 38948 3112 39004
rect 3180 38948 3236 39004
rect 3304 38948 3360 39004
rect 3428 38948 3484 39004
rect 3552 38948 3608 39004
rect 3676 38948 3732 39004
rect 3800 38948 3856 39004
rect 3924 38948 3980 39004
rect 4048 38948 4104 39004
rect 4172 38948 4228 39004
rect 4296 38948 4352 39004
rect 4420 38948 4476 39004
rect 4544 38948 4600 39004
rect 4668 38948 4724 39004
rect 2808 38824 2864 38880
rect 2932 38824 2988 38880
rect 3056 38824 3112 38880
rect 3180 38824 3236 38880
rect 3304 38824 3360 38880
rect 3428 38824 3484 38880
rect 3552 38824 3608 38880
rect 3676 38824 3732 38880
rect 3800 38824 3856 38880
rect 3924 38824 3980 38880
rect 4048 38824 4104 38880
rect 4172 38824 4228 38880
rect 4296 38824 4352 38880
rect 4420 38824 4476 38880
rect 4544 38824 4600 38880
rect 4668 38824 4724 38880
rect 2808 38700 2864 38756
rect 2932 38700 2988 38756
rect 3056 38700 3112 38756
rect 3180 38700 3236 38756
rect 3304 38700 3360 38756
rect 3428 38700 3484 38756
rect 3552 38700 3608 38756
rect 3676 38700 3732 38756
rect 3800 38700 3856 38756
rect 3924 38700 3980 38756
rect 4048 38700 4104 38756
rect 4172 38700 4228 38756
rect 4296 38700 4352 38756
rect 4420 38700 4476 38756
rect 4544 38700 4600 38756
rect 4668 38700 4724 38756
rect 2808 38576 2864 38632
rect 2932 38576 2988 38632
rect 3056 38576 3112 38632
rect 3180 38576 3236 38632
rect 3304 38576 3360 38632
rect 3428 38576 3484 38632
rect 3552 38576 3608 38632
rect 3676 38576 3732 38632
rect 3800 38576 3856 38632
rect 3924 38576 3980 38632
rect 4048 38576 4104 38632
rect 4172 38576 4228 38632
rect 4296 38576 4352 38632
rect 4420 38576 4476 38632
rect 4544 38576 4600 38632
rect 4668 38576 4724 38632
rect 2808 38452 2864 38508
rect 2932 38452 2988 38508
rect 3056 38452 3112 38508
rect 3180 38452 3236 38508
rect 3304 38452 3360 38508
rect 3428 38452 3484 38508
rect 3552 38452 3608 38508
rect 3676 38452 3732 38508
rect 3800 38452 3856 38508
rect 3924 38452 3980 38508
rect 4048 38452 4104 38508
rect 4172 38452 4228 38508
rect 4296 38452 4352 38508
rect 4420 38452 4476 38508
rect 4544 38452 4600 38508
rect 4668 38452 4724 38508
rect 5178 39692 5234 39748
rect 5302 39692 5358 39748
rect 5426 39692 5482 39748
rect 5550 39692 5606 39748
rect 5674 39692 5730 39748
rect 5798 39692 5854 39748
rect 5922 39692 5978 39748
rect 6046 39692 6102 39748
rect 6170 39692 6226 39748
rect 6294 39692 6350 39748
rect 6418 39692 6474 39748
rect 6542 39692 6598 39748
rect 6666 39692 6722 39748
rect 6790 39692 6846 39748
rect 6914 39692 6970 39748
rect 7038 39692 7094 39748
rect 5178 39568 5234 39624
rect 5302 39568 5358 39624
rect 5426 39568 5482 39624
rect 5550 39568 5606 39624
rect 5674 39568 5730 39624
rect 5798 39568 5854 39624
rect 5922 39568 5978 39624
rect 6046 39568 6102 39624
rect 6170 39568 6226 39624
rect 6294 39568 6350 39624
rect 6418 39568 6474 39624
rect 6542 39568 6598 39624
rect 6666 39568 6722 39624
rect 6790 39568 6846 39624
rect 6914 39568 6970 39624
rect 7038 39568 7094 39624
rect 5178 39444 5234 39500
rect 5302 39444 5358 39500
rect 5426 39444 5482 39500
rect 5550 39444 5606 39500
rect 5674 39444 5730 39500
rect 5798 39444 5854 39500
rect 5922 39444 5978 39500
rect 6046 39444 6102 39500
rect 6170 39444 6226 39500
rect 6294 39444 6350 39500
rect 6418 39444 6474 39500
rect 6542 39444 6598 39500
rect 6666 39444 6722 39500
rect 6790 39444 6846 39500
rect 6914 39444 6970 39500
rect 7038 39444 7094 39500
rect 5178 39320 5234 39376
rect 5302 39320 5358 39376
rect 5426 39320 5482 39376
rect 5550 39320 5606 39376
rect 5674 39320 5730 39376
rect 5798 39320 5854 39376
rect 5922 39320 5978 39376
rect 6046 39320 6102 39376
rect 6170 39320 6226 39376
rect 6294 39320 6350 39376
rect 6418 39320 6474 39376
rect 6542 39320 6598 39376
rect 6666 39320 6722 39376
rect 6790 39320 6846 39376
rect 6914 39320 6970 39376
rect 7038 39320 7094 39376
rect 5178 39196 5234 39252
rect 5302 39196 5358 39252
rect 5426 39196 5482 39252
rect 5550 39196 5606 39252
rect 5674 39196 5730 39252
rect 5798 39196 5854 39252
rect 5922 39196 5978 39252
rect 6046 39196 6102 39252
rect 6170 39196 6226 39252
rect 6294 39196 6350 39252
rect 6418 39196 6474 39252
rect 6542 39196 6598 39252
rect 6666 39196 6722 39252
rect 6790 39196 6846 39252
rect 6914 39196 6970 39252
rect 7038 39196 7094 39252
rect 5178 39072 5234 39128
rect 5302 39072 5358 39128
rect 5426 39072 5482 39128
rect 5550 39072 5606 39128
rect 5674 39072 5730 39128
rect 5798 39072 5854 39128
rect 5922 39072 5978 39128
rect 6046 39072 6102 39128
rect 6170 39072 6226 39128
rect 6294 39072 6350 39128
rect 6418 39072 6474 39128
rect 6542 39072 6598 39128
rect 6666 39072 6722 39128
rect 6790 39072 6846 39128
rect 6914 39072 6970 39128
rect 7038 39072 7094 39128
rect 5178 38948 5234 39004
rect 5302 38948 5358 39004
rect 5426 38948 5482 39004
rect 5550 38948 5606 39004
rect 5674 38948 5730 39004
rect 5798 38948 5854 39004
rect 5922 38948 5978 39004
rect 6046 38948 6102 39004
rect 6170 38948 6226 39004
rect 6294 38948 6350 39004
rect 6418 38948 6474 39004
rect 6542 38948 6598 39004
rect 6666 38948 6722 39004
rect 6790 38948 6846 39004
rect 6914 38948 6970 39004
rect 7038 38948 7094 39004
rect 5178 38824 5234 38880
rect 5302 38824 5358 38880
rect 5426 38824 5482 38880
rect 5550 38824 5606 38880
rect 5674 38824 5730 38880
rect 5798 38824 5854 38880
rect 5922 38824 5978 38880
rect 6046 38824 6102 38880
rect 6170 38824 6226 38880
rect 6294 38824 6350 38880
rect 6418 38824 6474 38880
rect 6542 38824 6598 38880
rect 6666 38824 6722 38880
rect 6790 38824 6846 38880
rect 6914 38824 6970 38880
rect 7038 38824 7094 38880
rect 5178 38700 5234 38756
rect 5302 38700 5358 38756
rect 5426 38700 5482 38756
rect 5550 38700 5606 38756
rect 5674 38700 5730 38756
rect 5798 38700 5854 38756
rect 5922 38700 5978 38756
rect 6046 38700 6102 38756
rect 6170 38700 6226 38756
rect 6294 38700 6350 38756
rect 6418 38700 6474 38756
rect 6542 38700 6598 38756
rect 6666 38700 6722 38756
rect 6790 38700 6846 38756
rect 6914 38700 6970 38756
rect 7038 38700 7094 38756
rect 5178 38576 5234 38632
rect 5302 38576 5358 38632
rect 5426 38576 5482 38632
rect 5550 38576 5606 38632
rect 5674 38576 5730 38632
rect 5798 38576 5854 38632
rect 5922 38576 5978 38632
rect 6046 38576 6102 38632
rect 6170 38576 6226 38632
rect 6294 38576 6350 38632
rect 6418 38576 6474 38632
rect 6542 38576 6598 38632
rect 6666 38576 6722 38632
rect 6790 38576 6846 38632
rect 6914 38576 6970 38632
rect 7038 38576 7094 38632
rect 5178 38452 5234 38508
rect 5302 38452 5358 38508
rect 5426 38452 5482 38508
rect 5550 38452 5606 38508
rect 5674 38452 5730 38508
rect 5798 38452 5854 38508
rect 5922 38452 5978 38508
rect 6046 38452 6102 38508
rect 6170 38452 6226 38508
rect 6294 38452 6350 38508
rect 6418 38452 6474 38508
rect 6542 38452 6598 38508
rect 6666 38452 6722 38508
rect 6790 38452 6846 38508
rect 6914 38452 6970 38508
rect 7038 38452 7094 38508
rect 7884 39692 7940 39748
rect 8008 39692 8064 39748
rect 8132 39692 8188 39748
rect 8256 39692 8312 39748
rect 8380 39692 8436 39748
rect 8504 39692 8560 39748
rect 8628 39692 8684 39748
rect 8752 39692 8808 39748
rect 8876 39692 8932 39748
rect 9000 39692 9056 39748
rect 9124 39692 9180 39748
rect 9248 39692 9304 39748
rect 9372 39692 9428 39748
rect 9496 39692 9552 39748
rect 9620 39692 9676 39748
rect 9744 39692 9800 39748
rect 7884 39568 7940 39624
rect 8008 39568 8064 39624
rect 8132 39568 8188 39624
rect 8256 39568 8312 39624
rect 8380 39568 8436 39624
rect 8504 39568 8560 39624
rect 8628 39568 8684 39624
rect 8752 39568 8808 39624
rect 8876 39568 8932 39624
rect 9000 39568 9056 39624
rect 9124 39568 9180 39624
rect 9248 39568 9304 39624
rect 9372 39568 9428 39624
rect 9496 39568 9552 39624
rect 9620 39568 9676 39624
rect 9744 39568 9800 39624
rect 7884 39444 7940 39500
rect 8008 39444 8064 39500
rect 8132 39444 8188 39500
rect 8256 39444 8312 39500
rect 8380 39444 8436 39500
rect 8504 39444 8560 39500
rect 8628 39444 8684 39500
rect 8752 39444 8808 39500
rect 8876 39444 8932 39500
rect 9000 39444 9056 39500
rect 9124 39444 9180 39500
rect 9248 39444 9304 39500
rect 9372 39444 9428 39500
rect 9496 39444 9552 39500
rect 9620 39444 9676 39500
rect 9744 39444 9800 39500
rect 7884 39320 7940 39376
rect 8008 39320 8064 39376
rect 8132 39320 8188 39376
rect 8256 39320 8312 39376
rect 8380 39320 8436 39376
rect 8504 39320 8560 39376
rect 8628 39320 8684 39376
rect 8752 39320 8808 39376
rect 8876 39320 8932 39376
rect 9000 39320 9056 39376
rect 9124 39320 9180 39376
rect 9248 39320 9304 39376
rect 9372 39320 9428 39376
rect 9496 39320 9552 39376
rect 9620 39320 9676 39376
rect 9744 39320 9800 39376
rect 7884 39196 7940 39252
rect 8008 39196 8064 39252
rect 8132 39196 8188 39252
rect 8256 39196 8312 39252
rect 8380 39196 8436 39252
rect 8504 39196 8560 39252
rect 8628 39196 8684 39252
rect 8752 39196 8808 39252
rect 8876 39196 8932 39252
rect 9000 39196 9056 39252
rect 9124 39196 9180 39252
rect 9248 39196 9304 39252
rect 9372 39196 9428 39252
rect 9496 39196 9552 39252
rect 9620 39196 9676 39252
rect 9744 39196 9800 39252
rect 7884 39072 7940 39128
rect 8008 39072 8064 39128
rect 8132 39072 8188 39128
rect 8256 39072 8312 39128
rect 8380 39072 8436 39128
rect 8504 39072 8560 39128
rect 8628 39072 8684 39128
rect 8752 39072 8808 39128
rect 8876 39072 8932 39128
rect 9000 39072 9056 39128
rect 9124 39072 9180 39128
rect 9248 39072 9304 39128
rect 9372 39072 9428 39128
rect 9496 39072 9552 39128
rect 9620 39072 9676 39128
rect 9744 39072 9800 39128
rect 7884 38948 7940 39004
rect 8008 38948 8064 39004
rect 8132 38948 8188 39004
rect 8256 38948 8312 39004
rect 8380 38948 8436 39004
rect 8504 38948 8560 39004
rect 8628 38948 8684 39004
rect 8752 38948 8808 39004
rect 8876 38948 8932 39004
rect 9000 38948 9056 39004
rect 9124 38948 9180 39004
rect 9248 38948 9304 39004
rect 9372 38948 9428 39004
rect 9496 38948 9552 39004
rect 9620 38948 9676 39004
rect 9744 38948 9800 39004
rect 7884 38824 7940 38880
rect 8008 38824 8064 38880
rect 8132 38824 8188 38880
rect 8256 38824 8312 38880
rect 8380 38824 8436 38880
rect 8504 38824 8560 38880
rect 8628 38824 8684 38880
rect 8752 38824 8808 38880
rect 8876 38824 8932 38880
rect 9000 38824 9056 38880
rect 9124 38824 9180 38880
rect 9248 38824 9304 38880
rect 9372 38824 9428 38880
rect 9496 38824 9552 38880
rect 9620 38824 9676 38880
rect 9744 38824 9800 38880
rect 7884 38700 7940 38756
rect 8008 38700 8064 38756
rect 8132 38700 8188 38756
rect 8256 38700 8312 38756
rect 8380 38700 8436 38756
rect 8504 38700 8560 38756
rect 8628 38700 8684 38756
rect 8752 38700 8808 38756
rect 8876 38700 8932 38756
rect 9000 38700 9056 38756
rect 9124 38700 9180 38756
rect 9248 38700 9304 38756
rect 9372 38700 9428 38756
rect 9496 38700 9552 38756
rect 9620 38700 9676 38756
rect 9744 38700 9800 38756
rect 7884 38576 7940 38632
rect 8008 38576 8064 38632
rect 8132 38576 8188 38632
rect 8256 38576 8312 38632
rect 8380 38576 8436 38632
rect 8504 38576 8560 38632
rect 8628 38576 8684 38632
rect 8752 38576 8808 38632
rect 8876 38576 8932 38632
rect 9000 38576 9056 38632
rect 9124 38576 9180 38632
rect 9248 38576 9304 38632
rect 9372 38576 9428 38632
rect 9496 38576 9552 38632
rect 9620 38576 9676 38632
rect 9744 38576 9800 38632
rect 7884 38452 7940 38508
rect 8008 38452 8064 38508
rect 8132 38452 8188 38508
rect 8256 38452 8312 38508
rect 8380 38452 8436 38508
rect 8504 38452 8560 38508
rect 8628 38452 8684 38508
rect 8752 38452 8808 38508
rect 8876 38452 8932 38508
rect 9000 38452 9056 38508
rect 9124 38452 9180 38508
rect 9248 38452 9304 38508
rect 9372 38452 9428 38508
rect 9496 38452 9552 38508
rect 9620 38452 9676 38508
rect 9744 38452 9800 38508
rect 10254 39692 10310 39748
rect 10378 39692 10434 39748
rect 10502 39692 10558 39748
rect 10626 39692 10682 39748
rect 10750 39692 10806 39748
rect 10874 39692 10930 39748
rect 10998 39692 11054 39748
rect 11122 39692 11178 39748
rect 11246 39692 11302 39748
rect 11370 39692 11426 39748
rect 11494 39692 11550 39748
rect 11618 39692 11674 39748
rect 11742 39692 11798 39748
rect 11866 39692 11922 39748
rect 11990 39692 12046 39748
rect 12114 39692 12170 39748
rect 10254 39568 10310 39624
rect 10378 39568 10434 39624
rect 10502 39568 10558 39624
rect 10626 39568 10682 39624
rect 10750 39568 10806 39624
rect 10874 39568 10930 39624
rect 10998 39568 11054 39624
rect 11122 39568 11178 39624
rect 11246 39568 11302 39624
rect 11370 39568 11426 39624
rect 11494 39568 11550 39624
rect 11618 39568 11674 39624
rect 11742 39568 11798 39624
rect 11866 39568 11922 39624
rect 11990 39568 12046 39624
rect 12114 39568 12170 39624
rect 10254 39444 10310 39500
rect 10378 39444 10434 39500
rect 10502 39444 10558 39500
rect 10626 39444 10682 39500
rect 10750 39444 10806 39500
rect 10874 39444 10930 39500
rect 10998 39444 11054 39500
rect 11122 39444 11178 39500
rect 11246 39444 11302 39500
rect 11370 39444 11426 39500
rect 11494 39444 11550 39500
rect 11618 39444 11674 39500
rect 11742 39444 11798 39500
rect 11866 39444 11922 39500
rect 11990 39444 12046 39500
rect 12114 39444 12170 39500
rect 10254 39320 10310 39376
rect 10378 39320 10434 39376
rect 10502 39320 10558 39376
rect 10626 39320 10682 39376
rect 10750 39320 10806 39376
rect 10874 39320 10930 39376
rect 10998 39320 11054 39376
rect 11122 39320 11178 39376
rect 11246 39320 11302 39376
rect 11370 39320 11426 39376
rect 11494 39320 11550 39376
rect 11618 39320 11674 39376
rect 11742 39320 11798 39376
rect 11866 39320 11922 39376
rect 11990 39320 12046 39376
rect 12114 39320 12170 39376
rect 10254 39196 10310 39252
rect 10378 39196 10434 39252
rect 10502 39196 10558 39252
rect 10626 39196 10682 39252
rect 10750 39196 10806 39252
rect 10874 39196 10930 39252
rect 10998 39196 11054 39252
rect 11122 39196 11178 39252
rect 11246 39196 11302 39252
rect 11370 39196 11426 39252
rect 11494 39196 11550 39252
rect 11618 39196 11674 39252
rect 11742 39196 11798 39252
rect 11866 39196 11922 39252
rect 11990 39196 12046 39252
rect 12114 39196 12170 39252
rect 10254 39072 10310 39128
rect 10378 39072 10434 39128
rect 10502 39072 10558 39128
rect 10626 39072 10682 39128
rect 10750 39072 10806 39128
rect 10874 39072 10930 39128
rect 10998 39072 11054 39128
rect 11122 39072 11178 39128
rect 11246 39072 11302 39128
rect 11370 39072 11426 39128
rect 11494 39072 11550 39128
rect 11618 39072 11674 39128
rect 11742 39072 11798 39128
rect 11866 39072 11922 39128
rect 11990 39072 12046 39128
rect 12114 39072 12170 39128
rect 10254 38948 10310 39004
rect 10378 38948 10434 39004
rect 10502 38948 10558 39004
rect 10626 38948 10682 39004
rect 10750 38948 10806 39004
rect 10874 38948 10930 39004
rect 10998 38948 11054 39004
rect 11122 38948 11178 39004
rect 11246 38948 11302 39004
rect 11370 38948 11426 39004
rect 11494 38948 11550 39004
rect 11618 38948 11674 39004
rect 11742 38948 11798 39004
rect 11866 38948 11922 39004
rect 11990 38948 12046 39004
rect 12114 38948 12170 39004
rect 10254 38824 10310 38880
rect 10378 38824 10434 38880
rect 10502 38824 10558 38880
rect 10626 38824 10682 38880
rect 10750 38824 10806 38880
rect 10874 38824 10930 38880
rect 10998 38824 11054 38880
rect 11122 38824 11178 38880
rect 11246 38824 11302 38880
rect 11370 38824 11426 38880
rect 11494 38824 11550 38880
rect 11618 38824 11674 38880
rect 11742 38824 11798 38880
rect 11866 38824 11922 38880
rect 11990 38824 12046 38880
rect 12114 38824 12170 38880
rect 10254 38700 10310 38756
rect 10378 38700 10434 38756
rect 10502 38700 10558 38756
rect 10626 38700 10682 38756
rect 10750 38700 10806 38756
rect 10874 38700 10930 38756
rect 10998 38700 11054 38756
rect 11122 38700 11178 38756
rect 11246 38700 11302 38756
rect 11370 38700 11426 38756
rect 11494 38700 11550 38756
rect 11618 38700 11674 38756
rect 11742 38700 11798 38756
rect 11866 38700 11922 38756
rect 11990 38700 12046 38756
rect 12114 38700 12170 38756
rect 10254 38576 10310 38632
rect 10378 38576 10434 38632
rect 10502 38576 10558 38632
rect 10626 38576 10682 38632
rect 10750 38576 10806 38632
rect 10874 38576 10930 38632
rect 10998 38576 11054 38632
rect 11122 38576 11178 38632
rect 11246 38576 11302 38632
rect 11370 38576 11426 38632
rect 11494 38576 11550 38632
rect 11618 38576 11674 38632
rect 11742 38576 11798 38632
rect 11866 38576 11922 38632
rect 11990 38576 12046 38632
rect 12114 38576 12170 38632
rect 10254 38452 10310 38508
rect 10378 38452 10434 38508
rect 10502 38452 10558 38508
rect 10626 38452 10682 38508
rect 10750 38452 10806 38508
rect 10874 38452 10930 38508
rect 10998 38452 11054 38508
rect 11122 38452 11178 38508
rect 11246 38452 11302 38508
rect 11370 38452 11426 38508
rect 11494 38452 11550 38508
rect 11618 38452 11674 38508
rect 11742 38452 11798 38508
rect 11866 38452 11922 38508
rect 11990 38452 12046 38508
rect 12114 38452 12170 38508
rect 12871 39692 12927 39748
rect 12995 39692 13051 39748
rect 13119 39692 13175 39748
rect 13243 39692 13299 39748
rect 13367 39692 13423 39748
rect 13491 39692 13547 39748
rect 13615 39692 13671 39748
rect 13739 39692 13795 39748
rect 13863 39692 13919 39748
rect 13987 39692 14043 39748
rect 14111 39692 14167 39748
rect 14235 39692 14291 39748
rect 14359 39692 14415 39748
rect 14483 39692 14539 39748
rect 14607 39692 14663 39748
rect 12871 39568 12927 39624
rect 12995 39568 13051 39624
rect 13119 39568 13175 39624
rect 13243 39568 13299 39624
rect 13367 39568 13423 39624
rect 13491 39568 13547 39624
rect 13615 39568 13671 39624
rect 13739 39568 13795 39624
rect 13863 39568 13919 39624
rect 13987 39568 14043 39624
rect 14111 39568 14167 39624
rect 14235 39568 14291 39624
rect 14359 39568 14415 39624
rect 14483 39568 14539 39624
rect 14607 39568 14663 39624
rect 12871 39444 12927 39500
rect 12995 39444 13051 39500
rect 13119 39444 13175 39500
rect 13243 39444 13299 39500
rect 13367 39444 13423 39500
rect 13491 39444 13547 39500
rect 13615 39444 13671 39500
rect 13739 39444 13795 39500
rect 13863 39444 13919 39500
rect 13987 39444 14043 39500
rect 14111 39444 14167 39500
rect 14235 39444 14291 39500
rect 14359 39444 14415 39500
rect 14483 39444 14539 39500
rect 14607 39444 14663 39500
rect 12871 39320 12927 39376
rect 12995 39320 13051 39376
rect 13119 39320 13175 39376
rect 13243 39320 13299 39376
rect 13367 39320 13423 39376
rect 13491 39320 13547 39376
rect 13615 39320 13671 39376
rect 13739 39320 13795 39376
rect 13863 39320 13919 39376
rect 13987 39320 14043 39376
rect 14111 39320 14167 39376
rect 14235 39320 14291 39376
rect 14359 39320 14415 39376
rect 14483 39320 14539 39376
rect 14607 39320 14663 39376
rect 12871 39196 12927 39252
rect 12995 39196 13051 39252
rect 13119 39196 13175 39252
rect 13243 39196 13299 39252
rect 13367 39196 13423 39252
rect 13491 39196 13547 39252
rect 13615 39196 13671 39252
rect 13739 39196 13795 39252
rect 13863 39196 13919 39252
rect 13987 39196 14043 39252
rect 14111 39196 14167 39252
rect 14235 39196 14291 39252
rect 14359 39196 14415 39252
rect 14483 39196 14539 39252
rect 14607 39196 14663 39252
rect 12871 39072 12927 39128
rect 12995 39072 13051 39128
rect 13119 39072 13175 39128
rect 13243 39072 13299 39128
rect 13367 39072 13423 39128
rect 13491 39072 13547 39128
rect 13615 39072 13671 39128
rect 13739 39072 13795 39128
rect 13863 39072 13919 39128
rect 13987 39072 14043 39128
rect 14111 39072 14167 39128
rect 14235 39072 14291 39128
rect 14359 39072 14415 39128
rect 14483 39072 14539 39128
rect 14607 39072 14663 39128
rect 12871 38948 12927 39004
rect 12995 38948 13051 39004
rect 13119 38948 13175 39004
rect 13243 38948 13299 39004
rect 13367 38948 13423 39004
rect 13491 38948 13547 39004
rect 13615 38948 13671 39004
rect 13739 38948 13795 39004
rect 13863 38948 13919 39004
rect 13987 38948 14043 39004
rect 14111 38948 14167 39004
rect 14235 38948 14291 39004
rect 14359 38948 14415 39004
rect 14483 38948 14539 39004
rect 14607 38948 14663 39004
rect 12871 38824 12927 38880
rect 12995 38824 13051 38880
rect 13119 38824 13175 38880
rect 13243 38824 13299 38880
rect 13367 38824 13423 38880
rect 13491 38824 13547 38880
rect 13615 38824 13671 38880
rect 13739 38824 13795 38880
rect 13863 38824 13919 38880
rect 13987 38824 14043 38880
rect 14111 38824 14167 38880
rect 14235 38824 14291 38880
rect 14359 38824 14415 38880
rect 14483 38824 14539 38880
rect 14607 38824 14663 38880
rect 12871 38700 12927 38756
rect 12995 38700 13051 38756
rect 13119 38700 13175 38756
rect 13243 38700 13299 38756
rect 13367 38700 13423 38756
rect 13491 38700 13547 38756
rect 13615 38700 13671 38756
rect 13739 38700 13795 38756
rect 13863 38700 13919 38756
rect 13987 38700 14043 38756
rect 14111 38700 14167 38756
rect 14235 38700 14291 38756
rect 14359 38700 14415 38756
rect 14483 38700 14539 38756
rect 14607 38700 14663 38756
rect 12871 38576 12927 38632
rect 12995 38576 13051 38632
rect 13119 38576 13175 38632
rect 13243 38576 13299 38632
rect 13367 38576 13423 38632
rect 13491 38576 13547 38632
rect 13615 38576 13671 38632
rect 13739 38576 13795 38632
rect 13863 38576 13919 38632
rect 13987 38576 14043 38632
rect 14111 38576 14167 38632
rect 14235 38576 14291 38632
rect 14359 38576 14415 38632
rect 14483 38576 14539 38632
rect 14607 38576 14663 38632
rect 12871 38452 12927 38508
rect 12995 38452 13051 38508
rect 13119 38452 13175 38508
rect 13243 38452 13299 38508
rect 13367 38452 13423 38508
rect 13491 38452 13547 38508
rect 13615 38452 13671 38508
rect 13739 38452 13795 38508
rect 13863 38452 13919 38508
rect 13987 38452 14043 38508
rect 14111 38452 14167 38508
rect 14235 38452 14291 38508
rect 14359 38452 14415 38508
rect 14483 38452 14539 38508
rect 14607 38452 14663 38508
rect 2289 38079 2345 38135
rect 2491 38098 2547 38154
rect 2615 38098 2671 38154
rect 4861 38098 4917 38154
rect 4985 38098 5041 38154
rect 7275 38098 7331 38154
rect 7399 38098 7455 38154
rect 7523 38098 7579 38154
rect 7647 38098 7703 38154
rect 9937 38098 9993 38154
rect 10061 38098 10117 38154
rect 12307 38098 12363 38154
rect 12431 38098 12487 38154
rect 2289 37947 2345 38003
rect 2491 37974 2547 38030
rect 2615 37974 2671 38030
rect 4861 37974 4917 38030
rect 4985 37974 5041 38030
rect 7275 37974 7331 38030
rect 7399 37974 7455 38030
rect 7523 37974 7579 38030
rect 7647 37974 7703 38030
rect 9937 37974 9993 38030
rect 10061 37974 10117 38030
rect 12307 37974 12363 38030
rect 12431 37974 12487 38030
rect 2289 37815 2345 37871
rect 2491 37850 2547 37906
rect 2615 37850 2671 37906
rect 4861 37850 4917 37906
rect 4985 37850 5041 37906
rect 7275 37850 7331 37906
rect 7399 37850 7455 37906
rect 7523 37850 7579 37906
rect 7647 37850 7703 37906
rect 9937 37850 9993 37906
rect 10061 37850 10117 37906
rect 12307 37850 12363 37906
rect 12431 37850 12487 37906
rect 2289 37683 2345 37739
rect 2491 37726 2547 37782
rect 2615 37726 2671 37782
rect 4861 37726 4917 37782
rect 4985 37726 5041 37782
rect 7275 37726 7331 37782
rect 7399 37726 7455 37782
rect 7523 37726 7579 37782
rect 7647 37726 7703 37782
rect 9937 37726 9993 37782
rect 10061 37726 10117 37782
rect 12307 37726 12363 37782
rect 12431 37726 12487 37782
rect 2289 37551 2345 37607
rect 2491 37602 2547 37658
rect 2615 37602 2671 37658
rect 4861 37602 4917 37658
rect 4985 37602 5041 37658
rect 7275 37602 7331 37658
rect 7399 37602 7455 37658
rect 7523 37602 7579 37658
rect 7647 37602 7703 37658
rect 9937 37602 9993 37658
rect 10061 37602 10117 37658
rect 12307 37602 12363 37658
rect 12431 37602 12487 37658
rect 2491 37478 2547 37534
rect 2615 37478 2671 37534
rect 4861 37478 4917 37534
rect 4985 37478 5041 37534
rect 7275 37478 7331 37534
rect 7399 37478 7455 37534
rect 7523 37478 7579 37534
rect 7647 37478 7703 37534
rect 9937 37478 9993 37534
rect 10061 37478 10117 37534
rect 12307 37478 12363 37534
rect 12431 37478 12487 37534
rect 2289 37419 2345 37475
rect 2491 37354 2547 37410
rect 2615 37354 2671 37410
rect 4861 37354 4917 37410
rect 4985 37354 5041 37410
rect 7275 37354 7331 37410
rect 7399 37354 7455 37410
rect 7523 37354 7579 37410
rect 7647 37354 7703 37410
rect 9937 37354 9993 37410
rect 10061 37354 10117 37410
rect 12307 37354 12363 37410
rect 12431 37354 12487 37410
rect 2289 37287 2345 37343
rect 2491 37230 2547 37286
rect 2615 37230 2671 37286
rect 4861 37230 4917 37286
rect 4985 37230 5041 37286
rect 7275 37230 7331 37286
rect 7399 37230 7455 37286
rect 7523 37230 7579 37286
rect 7647 37230 7703 37286
rect 9937 37230 9993 37286
rect 10061 37230 10117 37286
rect 12307 37230 12363 37286
rect 12431 37230 12487 37286
rect 2289 37155 2345 37211
rect 2491 37106 2547 37162
rect 2615 37106 2671 37162
rect 4861 37106 4917 37162
rect 4985 37106 5041 37162
rect 7275 37106 7331 37162
rect 7399 37106 7455 37162
rect 7523 37106 7579 37162
rect 7647 37106 7703 37162
rect 9937 37106 9993 37162
rect 10061 37106 10117 37162
rect 12307 37106 12363 37162
rect 12431 37106 12487 37162
rect 2289 37023 2345 37079
rect 2491 36982 2547 37038
rect 2615 36982 2671 37038
rect 4861 36982 4917 37038
rect 4985 36982 5041 37038
rect 7275 36982 7331 37038
rect 7399 36982 7455 37038
rect 7523 36982 7579 37038
rect 7647 36982 7703 37038
rect 9937 36982 9993 37038
rect 10061 36982 10117 37038
rect 12307 36982 12363 37038
rect 12431 36982 12487 37038
rect 2289 36891 2345 36947
rect 2491 36858 2547 36914
rect 2615 36858 2671 36914
rect 4861 36858 4917 36914
rect 4985 36858 5041 36914
rect 7275 36858 7331 36914
rect 7399 36858 7455 36914
rect 7523 36858 7579 36914
rect 7647 36858 7703 36914
rect 9937 36858 9993 36914
rect 10061 36858 10117 36914
rect 12307 36858 12363 36914
rect 12431 36858 12487 36914
rect 14902 38174 14958 38176
rect 14902 38122 14904 38174
rect 14904 38122 14956 38174
rect 14956 38122 14958 38174
rect 14902 38066 14958 38122
rect 14902 38014 14904 38066
rect 14904 38014 14956 38066
rect 14956 38014 14958 38066
rect 14902 37958 14958 38014
rect 14902 37906 14904 37958
rect 14904 37906 14956 37958
rect 14956 37906 14958 37958
rect 14902 37850 14958 37906
rect 14902 37798 14904 37850
rect 14904 37798 14956 37850
rect 14956 37798 14958 37850
rect 14902 37742 14958 37798
rect 14902 37690 14904 37742
rect 14904 37690 14956 37742
rect 14956 37690 14958 37742
rect 14902 37634 14958 37690
rect 14902 37582 14904 37634
rect 14904 37582 14956 37634
rect 14956 37582 14958 37634
rect 14902 37526 14958 37582
rect 14902 37474 14904 37526
rect 14904 37474 14956 37526
rect 14956 37474 14958 37526
rect 14902 37418 14958 37474
rect 14902 37366 14904 37418
rect 14904 37366 14956 37418
rect 14956 37366 14958 37418
rect 14902 37310 14958 37366
rect 14902 37258 14904 37310
rect 14904 37258 14956 37310
rect 14956 37258 14958 37310
rect 14902 37202 14958 37258
rect 14902 37150 14904 37202
rect 14904 37150 14956 37202
rect 14956 37150 14958 37202
rect 14902 37094 14958 37150
rect 14902 37042 14904 37094
rect 14904 37042 14956 37094
rect 14956 37042 14958 37094
rect 14902 36986 14958 37042
rect 14902 36934 14904 36986
rect 14904 36934 14956 36986
rect 14956 36934 14958 36986
rect 14902 36878 14958 36934
rect 14902 36826 14904 36878
rect 14904 36826 14956 36878
rect 14956 36826 14958 36878
rect 14902 36824 14958 36826
<< metal3 >>
rect 2481 56043 2681 57235
rect 4851 56043 5051 57235
rect 7265 56043 7713 57235
rect 9927 56043 10127 57235
rect 12297 56043 12497 57235
rect 305 54442 2117 55758
rect 2798 54442 4734 55758
rect 5168 54442 7104 55758
rect 7874 54442 9810 55758
rect 10244 54442 12180 55758
rect 12861 54442 14673 55758
rect 2481 52842 2681 54158
rect 4851 52842 5051 54158
rect 7265 52842 7713 54158
rect 9927 52842 10127 54158
rect 12297 52842 12497 54158
rect -11 52576 14989 52600
rect -11 51224 20 52576
rect 76 52548 14902 52576
rect 76 52521 2491 52548
rect 76 52465 2289 52521
rect 2345 52492 2491 52521
rect 2547 52492 2615 52548
rect 2671 52492 4861 52548
rect 4917 52492 4985 52548
rect 5041 52492 7275 52548
rect 7331 52492 7399 52548
rect 7455 52492 7523 52548
rect 7579 52492 7647 52548
rect 7703 52492 9937 52548
rect 9993 52492 10061 52548
rect 10117 52492 12307 52548
rect 12363 52492 12431 52548
rect 12487 52492 14902 52548
rect 2345 52465 14902 52492
rect 76 52424 14902 52465
rect 76 52389 2491 52424
rect 76 52333 2289 52389
rect 2345 52368 2491 52389
rect 2547 52368 2615 52424
rect 2671 52368 4861 52424
rect 4917 52368 4985 52424
rect 5041 52368 7275 52424
rect 7331 52368 7399 52424
rect 7455 52368 7523 52424
rect 7579 52368 7647 52424
rect 7703 52368 9937 52424
rect 9993 52368 10061 52424
rect 10117 52368 12307 52424
rect 12363 52368 12431 52424
rect 12487 52368 14902 52424
rect 2345 52333 14902 52368
rect 76 52300 14902 52333
rect 76 52257 2491 52300
rect 76 52201 2289 52257
rect 2345 52244 2491 52257
rect 2547 52244 2615 52300
rect 2671 52244 4861 52300
rect 4917 52244 4985 52300
rect 5041 52244 7275 52300
rect 7331 52244 7399 52300
rect 7455 52244 7523 52300
rect 7579 52244 7647 52300
rect 7703 52244 9937 52300
rect 9993 52244 10061 52300
rect 10117 52244 12307 52300
rect 12363 52244 12431 52300
rect 12487 52244 14902 52300
rect 2345 52201 14902 52244
rect 76 52176 14902 52201
rect 76 52125 2491 52176
rect 76 52069 2289 52125
rect 2345 52120 2491 52125
rect 2547 52120 2615 52176
rect 2671 52120 4861 52176
rect 4917 52120 4985 52176
rect 5041 52120 7275 52176
rect 7331 52120 7399 52176
rect 7455 52120 7523 52176
rect 7579 52120 7647 52176
rect 7703 52120 9937 52176
rect 9993 52120 10061 52176
rect 10117 52120 12307 52176
rect 12363 52120 12431 52176
rect 12487 52120 14902 52176
rect 2345 52069 14902 52120
rect 76 52052 14902 52069
rect 76 51996 2491 52052
rect 2547 51996 2615 52052
rect 2671 51996 4861 52052
rect 4917 51996 4985 52052
rect 5041 51996 7275 52052
rect 7331 51996 7399 52052
rect 7455 51996 7523 52052
rect 7579 51996 7647 52052
rect 7703 51996 9937 52052
rect 9993 51996 10061 52052
rect 10117 51996 12307 52052
rect 12363 51996 12431 52052
rect 12487 51996 14902 52052
rect 76 51993 14902 51996
rect 76 51937 2289 51993
rect 2345 51937 14902 51993
rect 76 51928 14902 51937
rect 76 51872 2491 51928
rect 2547 51872 2615 51928
rect 2671 51872 4861 51928
rect 4917 51872 4985 51928
rect 5041 51872 7275 51928
rect 7331 51872 7399 51928
rect 7455 51872 7523 51928
rect 7579 51872 7647 51928
rect 7703 51872 9937 51928
rect 9993 51872 10061 51928
rect 10117 51872 12307 51928
rect 12363 51872 12431 51928
rect 12487 51872 14902 51928
rect 76 51861 14902 51872
rect 76 51805 2289 51861
rect 2345 51805 14902 51861
rect 76 51804 14902 51805
rect 76 51748 2491 51804
rect 2547 51748 2615 51804
rect 2671 51748 4861 51804
rect 4917 51748 4985 51804
rect 5041 51748 7275 51804
rect 7331 51748 7399 51804
rect 7455 51748 7523 51804
rect 7579 51748 7647 51804
rect 7703 51748 9937 51804
rect 9993 51748 10061 51804
rect 10117 51748 12307 51804
rect 12363 51748 12431 51804
rect 12487 51748 14902 51804
rect 76 51729 14902 51748
rect 76 51673 2289 51729
rect 2345 51680 14902 51729
rect 2345 51673 2491 51680
rect 76 51624 2491 51673
rect 2547 51624 2615 51680
rect 2671 51624 4861 51680
rect 4917 51624 4985 51680
rect 5041 51624 7275 51680
rect 7331 51624 7399 51680
rect 7455 51624 7523 51680
rect 7579 51624 7647 51680
rect 7703 51624 9937 51680
rect 9993 51624 10061 51680
rect 10117 51624 12307 51680
rect 12363 51624 12431 51680
rect 12487 51624 14902 51680
rect 76 51597 14902 51624
rect 76 51541 2289 51597
rect 2345 51556 14902 51597
rect 2345 51541 2491 51556
rect 76 51500 2491 51541
rect 2547 51500 2615 51556
rect 2671 51500 4861 51556
rect 4917 51500 4985 51556
rect 5041 51500 7275 51556
rect 7331 51500 7399 51556
rect 7455 51500 7523 51556
rect 7579 51500 7647 51556
rect 7703 51500 9937 51556
rect 9993 51500 10061 51556
rect 10117 51500 12307 51556
rect 12363 51500 12431 51556
rect 12487 51500 14902 51556
rect 76 51465 14902 51500
rect 76 51409 2289 51465
rect 2345 51432 14902 51465
rect 2345 51409 2491 51432
rect 76 51376 2491 51409
rect 2547 51376 2615 51432
rect 2671 51376 4861 51432
rect 4917 51376 4985 51432
rect 5041 51376 7275 51432
rect 7331 51376 7399 51432
rect 7455 51376 7523 51432
rect 7579 51376 7647 51432
rect 7703 51376 9937 51432
rect 9993 51376 10061 51432
rect 10117 51376 12307 51432
rect 12363 51376 12431 51432
rect 12487 51376 14902 51432
rect 76 51333 14902 51376
rect 76 51277 2289 51333
rect 2345 51308 14902 51333
rect 2345 51277 2491 51308
rect 76 51252 2491 51277
rect 2547 51252 2615 51308
rect 2671 51252 4861 51308
rect 4917 51252 4985 51308
rect 5041 51252 7275 51308
rect 7331 51252 7399 51308
rect 7455 51252 7523 51308
rect 7579 51252 7647 51308
rect 7703 51252 9937 51308
rect 9993 51252 10061 51308
rect 10117 51252 12307 51308
rect 12363 51252 12431 51308
rect 12487 51252 14902 51308
rect 76 51224 14902 51252
rect 14958 51224 14989 52576
rect -11 51200 14989 51224
rect 139 50948 14839 50980
rect 139 50892 315 50948
rect 371 50892 439 50948
rect 495 50892 563 50948
rect 619 50892 687 50948
rect 743 50892 811 50948
rect 867 50892 935 50948
rect 991 50892 1059 50948
rect 1115 50892 1183 50948
rect 1239 50892 1307 50948
rect 1363 50892 1431 50948
rect 1487 50892 1555 50948
rect 1611 50892 1679 50948
rect 1735 50892 1803 50948
rect 1859 50892 1927 50948
rect 1983 50892 2051 50948
rect 2107 50892 2808 50948
rect 2864 50892 2932 50948
rect 2988 50892 3056 50948
rect 3112 50892 3180 50948
rect 3236 50892 3304 50948
rect 3360 50892 3428 50948
rect 3484 50892 3552 50948
rect 3608 50892 3676 50948
rect 3732 50892 3800 50948
rect 3856 50892 3924 50948
rect 3980 50892 4048 50948
rect 4104 50892 4172 50948
rect 4228 50892 4296 50948
rect 4352 50892 4420 50948
rect 4476 50892 4544 50948
rect 4600 50892 4668 50948
rect 4724 50892 5178 50948
rect 5234 50892 5302 50948
rect 5358 50892 5426 50948
rect 5482 50892 5550 50948
rect 5606 50892 5674 50948
rect 5730 50892 5798 50948
rect 5854 50892 5922 50948
rect 5978 50892 6046 50948
rect 6102 50892 6170 50948
rect 6226 50892 6294 50948
rect 6350 50892 6418 50948
rect 6474 50892 6542 50948
rect 6598 50892 6666 50948
rect 6722 50892 6790 50948
rect 6846 50892 6914 50948
rect 6970 50892 7038 50948
rect 7094 50892 7884 50948
rect 7940 50892 8008 50948
rect 8064 50892 8132 50948
rect 8188 50892 8256 50948
rect 8312 50892 8380 50948
rect 8436 50892 8504 50948
rect 8560 50892 8628 50948
rect 8684 50892 8752 50948
rect 8808 50892 8876 50948
rect 8932 50892 9000 50948
rect 9056 50892 9124 50948
rect 9180 50892 9248 50948
rect 9304 50892 9372 50948
rect 9428 50892 9496 50948
rect 9552 50892 9620 50948
rect 9676 50892 9744 50948
rect 9800 50892 10254 50948
rect 10310 50892 10378 50948
rect 10434 50892 10502 50948
rect 10558 50892 10626 50948
rect 10682 50892 10750 50948
rect 10806 50892 10874 50948
rect 10930 50892 10998 50948
rect 11054 50892 11122 50948
rect 11178 50892 11246 50948
rect 11302 50892 11370 50948
rect 11426 50892 11494 50948
rect 11550 50892 11618 50948
rect 11674 50892 11742 50948
rect 11798 50892 11866 50948
rect 11922 50892 11990 50948
rect 12046 50892 12114 50948
rect 12170 50892 12871 50948
rect 12927 50892 12995 50948
rect 13051 50892 13119 50948
rect 13175 50892 13243 50948
rect 13299 50892 13367 50948
rect 13423 50892 13491 50948
rect 13547 50892 13615 50948
rect 13671 50892 13739 50948
rect 13795 50892 13863 50948
rect 13919 50892 13987 50948
rect 14043 50892 14111 50948
rect 14167 50892 14235 50948
rect 14291 50892 14359 50948
rect 14415 50892 14483 50948
rect 14539 50892 14607 50948
rect 14663 50892 14839 50948
rect 139 50824 14839 50892
rect 139 50768 315 50824
rect 371 50768 439 50824
rect 495 50768 563 50824
rect 619 50768 687 50824
rect 743 50768 811 50824
rect 867 50768 935 50824
rect 991 50768 1059 50824
rect 1115 50768 1183 50824
rect 1239 50768 1307 50824
rect 1363 50768 1431 50824
rect 1487 50768 1555 50824
rect 1611 50768 1679 50824
rect 1735 50768 1803 50824
rect 1859 50768 1927 50824
rect 1983 50768 2051 50824
rect 2107 50768 2808 50824
rect 2864 50768 2932 50824
rect 2988 50768 3056 50824
rect 3112 50768 3180 50824
rect 3236 50768 3304 50824
rect 3360 50768 3428 50824
rect 3484 50768 3552 50824
rect 3608 50768 3676 50824
rect 3732 50768 3800 50824
rect 3856 50768 3924 50824
rect 3980 50768 4048 50824
rect 4104 50768 4172 50824
rect 4228 50768 4296 50824
rect 4352 50768 4420 50824
rect 4476 50768 4544 50824
rect 4600 50768 4668 50824
rect 4724 50768 5178 50824
rect 5234 50768 5302 50824
rect 5358 50768 5426 50824
rect 5482 50768 5550 50824
rect 5606 50768 5674 50824
rect 5730 50768 5798 50824
rect 5854 50768 5922 50824
rect 5978 50768 6046 50824
rect 6102 50768 6170 50824
rect 6226 50768 6294 50824
rect 6350 50768 6418 50824
rect 6474 50768 6542 50824
rect 6598 50768 6666 50824
rect 6722 50768 6790 50824
rect 6846 50768 6914 50824
rect 6970 50768 7038 50824
rect 7094 50768 7884 50824
rect 7940 50768 8008 50824
rect 8064 50768 8132 50824
rect 8188 50768 8256 50824
rect 8312 50768 8380 50824
rect 8436 50768 8504 50824
rect 8560 50768 8628 50824
rect 8684 50768 8752 50824
rect 8808 50768 8876 50824
rect 8932 50768 9000 50824
rect 9056 50768 9124 50824
rect 9180 50768 9248 50824
rect 9304 50768 9372 50824
rect 9428 50768 9496 50824
rect 9552 50768 9620 50824
rect 9676 50768 9744 50824
rect 9800 50768 10254 50824
rect 10310 50768 10378 50824
rect 10434 50768 10502 50824
rect 10558 50768 10626 50824
rect 10682 50768 10750 50824
rect 10806 50768 10874 50824
rect 10930 50768 10998 50824
rect 11054 50768 11122 50824
rect 11178 50768 11246 50824
rect 11302 50768 11370 50824
rect 11426 50768 11494 50824
rect 11550 50768 11618 50824
rect 11674 50768 11742 50824
rect 11798 50768 11866 50824
rect 11922 50768 11990 50824
rect 12046 50768 12114 50824
rect 12170 50768 12871 50824
rect 12927 50768 12995 50824
rect 13051 50768 13119 50824
rect 13175 50768 13243 50824
rect 13299 50768 13367 50824
rect 13423 50768 13491 50824
rect 13547 50768 13615 50824
rect 13671 50768 13739 50824
rect 13795 50768 13863 50824
rect 13919 50768 13987 50824
rect 14043 50768 14111 50824
rect 14167 50768 14235 50824
rect 14291 50768 14359 50824
rect 14415 50768 14483 50824
rect 14539 50768 14607 50824
rect 14663 50768 14839 50824
rect 139 50700 14839 50768
rect 139 50644 315 50700
rect 371 50644 439 50700
rect 495 50644 563 50700
rect 619 50644 687 50700
rect 743 50644 811 50700
rect 867 50644 935 50700
rect 991 50644 1059 50700
rect 1115 50644 1183 50700
rect 1239 50644 1307 50700
rect 1363 50644 1431 50700
rect 1487 50644 1555 50700
rect 1611 50644 1679 50700
rect 1735 50644 1803 50700
rect 1859 50644 1927 50700
rect 1983 50644 2051 50700
rect 2107 50644 2808 50700
rect 2864 50644 2932 50700
rect 2988 50644 3056 50700
rect 3112 50644 3180 50700
rect 3236 50644 3304 50700
rect 3360 50644 3428 50700
rect 3484 50644 3552 50700
rect 3608 50644 3676 50700
rect 3732 50644 3800 50700
rect 3856 50644 3924 50700
rect 3980 50644 4048 50700
rect 4104 50644 4172 50700
rect 4228 50644 4296 50700
rect 4352 50644 4420 50700
rect 4476 50644 4544 50700
rect 4600 50644 4668 50700
rect 4724 50644 5178 50700
rect 5234 50644 5302 50700
rect 5358 50644 5426 50700
rect 5482 50644 5550 50700
rect 5606 50644 5674 50700
rect 5730 50644 5798 50700
rect 5854 50644 5922 50700
rect 5978 50644 6046 50700
rect 6102 50644 6170 50700
rect 6226 50644 6294 50700
rect 6350 50644 6418 50700
rect 6474 50644 6542 50700
rect 6598 50644 6666 50700
rect 6722 50644 6790 50700
rect 6846 50644 6914 50700
rect 6970 50644 7038 50700
rect 7094 50644 7884 50700
rect 7940 50644 8008 50700
rect 8064 50644 8132 50700
rect 8188 50644 8256 50700
rect 8312 50644 8380 50700
rect 8436 50644 8504 50700
rect 8560 50644 8628 50700
rect 8684 50644 8752 50700
rect 8808 50644 8876 50700
rect 8932 50644 9000 50700
rect 9056 50644 9124 50700
rect 9180 50644 9248 50700
rect 9304 50644 9372 50700
rect 9428 50644 9496 50700
rect 9552 50644 9620 50700
rect 9676 50644 9744 50700
rect 9800 50644 10254 50700
rect 10310 50644 10378 50700
rect 10434 50644 10502 50700
rect 10558 50644 10626 50700
rect 10682 50644 10750 50700
rect 10806 50644 10874 50700
rect 10930 50644 10998 50700
rect 11054 50644 11122 50700
rect 11178 50644 11246 50700
rect 11302 50644 11370 50700
rect 11426 50644 11494 50700
rect 11550 50644 11618 50700
rect 11674 50644 11742 50700
rect 11798 50644 11866 50700
rect 11922 50644 11990 50700
rect 12046 50644 12114 50700
rect 12170 50644 12871 50700
rect 12927 50644 12995 50700
rect 13051 50644 13119 50700
rect 13175 50644 13243 50700
rect 13299 50644 13367 50700
rect 13423 50644 13491 50700
rect 13547 50644 13615 50700
rect 13671 50644 13739 50700
rect 13795 50644 13863 50700
rect 13919 50644 13987 50700
rect 14043 50644 14111 50700
rect 14167 50644 14235 50700
rect 14291 50644 14359 50700
rect 14415 50644 14483 50700
rect 14539 50644 14607 50700
rect 14663 50644 14839 50700
rect 139 50576 14839 50644
rect 139 50520 315 50576
rect 371 50520 439 50576
rect 495 50520 563 50576
rect 619 50520 687 50576
rect 743 50520 811 50576
rect 867 50520 935 50576
rect 991 50520 1059 50576
rect 1115 50520 1183 50576
rect 1239 50520 1307 50576
rect 1363 50520 1431 50576
rect 1487 50520 1555 50576
rect 1611 50520 1679 50576
rect 1735 50520 1803 50576
rect 1859 50520 1927 50576
rect 1983 50520 2051 50576
rect 2107 50520 2808 50576
rect 2864 50520 2932 50576
rect 2988 50520 3056 50576
rect 3112 50520 3180 50576
rect 3236 50520 3304 50576
rect 3360 50520 3428 50576
rect 3484 50520 3552 50576
rect 3608 50520 3676 50576
rect 3732 50520 3800 50576
rect 3856 50520 3924 50576
rect 3980 50520 4048 50576
rect 4104 50520 4172 50576
rect 4228 50520 4296 50576
rect 4352 50520 4420 50576
rect 4476 50520 4544 50576
rect 4600 50520 4668 50576
rect 4724 50520 5178 50576
rect 5234 50520 5302 50576
rect 5358 50520 5426 50576
rect 5482 50520 5550 50576
rect 5606 50520 5674 50576
rect 5730 50520 5798 50576
rect 5854 50520 5922 50576
rect 5978 50520 6046 50576
rect 6102 50520 6170 50576
rect 6226 50520 6294 50576
rect 6350 50520 6418 50576
rect 6474 50520 6542 50576
rect 6598 50520 6666 50576
rect 6722 50520 6790 50576
rect 6846 50520 6914 50576
rect 6970 50520 7038 50576
rect 7094 50520 7884 50576
rect 7940 50520 8008 50576
rect 8064 50520 8132 50576
rect 8188 50520 8256 50576
rect 8312 50520 8380 50576
rect 8436 50520 8504 50576
rect 8560 50520 8628 50576
rect 8684 50520 8752 50576
rect 8808 50520 8876 50576
rect 8932 50520 9000 50576
rect 9056 50520 9124 50576
rect 9180 50520 9248 50576
rect 9304 50520 9372 50576
rect 9428 50520 9496 50576
rect 9552 50520 9620 50576
rect 9676 50520 9744 50576
rect 9800 50520 10254 50576
rect 10310 50520 10378 50576
rect 10434 50520 10502 50576
rect 10558 50520 10626 50576
rect 10682 50520 10750 50576
rect 10806 50520 10874 50576
rect 10930 50520 10998 50576
rect 11054 50520 11122 50576
rect 11178 50520 11246 50576
rect 11302 50520 11370 50576
rect 11426 50520 11494 50576
rect 11550 50520 11618 50576
rect 11674 50520 11742 50576
rect 11798 50520 11866 50576
rect 11922 50520 11990 50576
rect 12046 50520 12114 50576
rect 12170 50520 12871 50576
rect 12927 50520 12995 50576
rect 13051 50520 13119 50576
rect 13175 50520 13243 50576
rect 13299 50520 13367 50576
rect 13423 50520 13491 50576
rect 13547 50520 13615 50576
rect 13671 50520 13739 50576
rect 13795 50520 13863 50576
rect 13919 50520 13987 50576
rect 14043 50520 14111 50576
rect 14167 50520 14235 50576
rect 14291 50520 14359 50576
rect 14415 50520 14483 50576
rect 14539 50520 14607 50576
rect 14663 50520 14839 50576
rect 139 50452 14839 50520
rect 139 50396 315 50452
rect 371 50396 439 50452
rect 495 50396 563 50452
rect 619 50396 687 50452
rect 743 50396 811 50452
rect 867 50396 935 50452
rect 991 50396 1059 50452
rect 1115 50396 1183 50452
rect 1239 50396 1307 50452
rect 1363 50396 1431 50452
rect 1487 50396 1555 50452
rect 1611 50396 1679 50452
rect 1735 50396 1803 50452
rect 1859 50396 1927 50452
rect 1983 50396 2051 50452
rect 2107 50396 2808 50452
rect 2864 50396 2932 50452
rect 2988 50396 3056 50452
rect 3112 50396 3180 50452
rect 3236 50396 3304 50452
rect 3360 50396 3428 50452
rect 3484 50396 3552 50452
rect 3608 50396 3676 50452
rect 3732 50396 3800 50452
rect 3856 50396 3924 50452
rect 3980 50396 4048 50452
rect 4104 50396 4172 50452
rect 4228 50396 4296 50452
rect 4352 50396 4420 50452
rect 4476 50396 4544 50452
rect 4600 50396 4668 50452
rect 4724 50396 5178 50452
rect 5234 50396 5302 50452
rect 5358 50396 5426 50452
rect 5482 50396 5550 50452
rect 5606 50396 5674 50452
rect 5730 50396 5798 50452
rect 5854 50396 5922 50452
rect 5978 50396 6046 50452
rect 6102 50396 6170 50452
rect 6226 50396 6294 50452
rect 6350 50396 6418 50452
rect 6474 50396 6542 50452
rect 6598 50396 6666 50452
rect 6722 50396 6790 50452
rect 6846 50396 6914 50452
rect 6970 50396 7038 50452
rect 7094 50396 7884 50452
rect 7940 50396 8008 50452
rect 8064 50396 8132 50452
rect 8188 50396 8256 50452
rect 8312 50396 8380 50452
rect 8436 50396 8504 50452
rect 8560 50396 8628 50452
rect 8684 50396 8752 50452
rect 8808 50396 8876 50452
rect 8932 50396 9000 50452
rect 9056 50396 9124 50452
rect 9180 50396 9248 50452
rect 9304 50396 9372 50452
rect 9428 50396 9496 50452
rect 9552 50396 9620 50452
rect 9676 50396 9744 50452
rect 9800 50396 10254 50452
rect 10310 50396 10378 50452
rect 10434 50396 10502 50452
rect 10558 50396 10626 50452
rect 10682 50396 10750 50452
rect 10806 50396 10874 50452
rect 10930 50396 10998 50452
rect 11054 50396 11122 50452
rect 11178 50396 11246 50452
rect 11302 50396 11370 50452
rect 11426 50396 11494 50452
rect 11550 50396 11618 50452
rect 11674 50396 11742 50452
rect 11798 50396 11866 50452
rect 11922 50396 11990 50452
rect 12046 50396 12114 50452
rect 12170 50396 12871 50452
rect 12927 50396 12995 50452
rect 13051 50396 13119 50452
rect 13175 50396 13243 50452
rect 13299 50396 13367 50452
rect 13423 50396 13491 50452
rect 13547 50396 13615 50452
rect 13671 50396 13739 50452
rect 13795 50396 13863 50452
rect 13919 50396 13987 50452
rect 14043 50396 14111 50452
rect 14167 50396 14235 50452
rect 14291 50396 14359 50452
rect 14415 50396 14483 50452
rect 14539 50396 14607 50452
rect 14663 50396 14839 50452
rect 139 50328 14839 50396
rect 139 50272 315 50328
rect 371 50272 439 50328
rect 495 50272 563 50328
rect 619 50272 687 50328
rect 743 50272 811 50328
rect 867 50272 935 50328
rect 991 50272 1059 50328
rect 1115 50272 1183 50328
rect 1239 50272 1307 50328
rect 1363 50272 1431 50328
rect 1487 50272 1555 50328
rect 1611 50272 1679 50328
rect 1735 50272 1803 50328
rect 1859 50272 1927 50328
rect 1983 50272 2051 50328
rect 2107 50272 2808 50328
rect 2864 50272 2932 50328
rect 2988 50272 3056 50328
rect 3112 50272 3180 50328
rect 3236 50272 3304 50328
rect 3360 50272 3428 50328
rect 3484 50272 3552 50328
rect 3608 50272 3676 50328
rect 3732 50272 3800 50328
rect 3856 50272 3924 50328
rect 3980 50272 4048 50328
rect 4104 50272 4172 50328
rect 4228 50272 4296 50328
rect 4352 50272 4420 50328
rect 4476 50272 4544 50328
rect 4600 50272 4668 50328
rect 4724 50272 5178 50328
rect 5234 50272 5302 50328
rect 5358 50272 5426 50328
rect 5482 50272 5550 50328
rect 5606 50272 5674 50328
rect 5730 50272 5798 50328
rect 5854 50272 5922 50328
rect 5978 50272 6046 50328
rect 6102 50272 6170 50328
rect 6226 50272 6294 50328
rect 6350 50272 6418 50328
rect 6474 50272 6542 50328
rect 6598 50272 6666 50328
rect 6722 50272 6790 50328
rect 6846 50272 6914 50328
rect 6970 50272 7038 50328
rect 7094 50272 7884 50328
rect 7940 50272 8008 50328
rect 8064 50272 8132 50328
rect 8188 50272 8256 50328
rect 8312 50272 8380 50328
rect 8436 50272 8504 50328
rect 8560 50272 8628 50328
rect 8684 50272 8752 50328
rect 8808 50272 8876 50328
rect 8932 50272 9000 50328
rect 9056 50272 9124 50328
rect 9180 50272 9248 50328
rect 9304 50272 9372 50328
rect 9428 50272 9496 50328
rect 9552 50272 9620 50328
rect 9676 50272 9744 50328
rect 9800 50272 10254 50328
rect 10310 50272 10378 50328
rect 10434 50272 10502 50328
rect 10558 50272 10626 50328
rect 10682 50272 10750 50328
rect 10806 50272 10874 50328
rect 10930 50272 10998 50328
rect 11054 50272 11122 50328
rect 11178 50272 11246 50328
rect 11302 50272 11370 50328
rect 11426 50272 11494 50328
rect 11550 50272 11618 50328
rect 11674 50272 11742 50328
rect 11798 50272 11866 50328
rect 11922 50272 11990 50328
rect 12046 50272 12114 50328
rect 12170 50272 12871 50328
rect 12927 50272 12995 50328
rect 13051 50272 13119 50328
rect 13175 50272 13243 50328
rect 13299 50272 13367 50328
rect 13423 50272 13491 50328
rect 13547 50272 13615 50328
rect 13671 50272 13739 50328
rect 13795 50272 13863 50328
rect 13919 50272 13987 50328
rect 14043 50272 14111 50328
rect 14167 50272 14235 50328
rect 14291 50272 14359 50328
rect 14415 50272 14483 50328
rect 14539 50272 14607 50328
rect 14663 50272 14839 50328
rect 139 50204 14839 50272
rect 139 50148 315 50204
rect 371 50148 439 50204
rect 495 50148 563 50204
rect 619 50148 687 50204
rect 743 50148 811 50204
rect 867 50148 935 50204
rect 991 50148 1059 50204
rect 1115 50148 1183 50204
rect 1239 50148 1307 50204
rect 1363 50148 1431 50204
rect 1487 50148 1555 50204
rect 1611 50148 1679 50204
rect 1735 50148 1803 50204
rect 1859 50148 1927 50204
rect 1983 50148 2051 50204
rect 2107 50148 2808 50204
rect 2864 50148 2932 50204
rect 2988 50148 3056 50204
rect 3112 50148 3180 50204
rect 3236 50148 3304 50204
rect 3360 50148 3428 50204
rect 3484 50148 3552 50204
rect 3608 50148 3676 50204
rect 3732 50148 3800 50204
rect 3856 50148 3924 50204
rect 3980 50148 4048 50204
rect 4104 50148 4172 50204
rect 4228 50148 4296 50204
rect 4352 50148 4420 50204
rect 4476 50148 4544 50204
rect 4600 50148 4668 50204
rect 4724 50148 5178 50204
rect 5234 50148 5302 50204
rect 5358 50148 5426 50204
rect 5482 50148 5550 50204
rect 5606 50148 5674 50204
rect 5730 50148 5798 50204
rect 5854 50148 5922 50204
rect 5978 50148 6046 50204
rect 6102 50148 6170 50204
rect 6226 50148 6294 50204
rect 6350 50148 6418 50204
rect 6474 50148 6542 50204
rect 6598 50148 6666 50204
rect 6722 50148 6790 50204
rect 6846 50148 6914 50204
rect 6970 50148 7038 50204
rect 7094 50148 7884 50204
rect 7940 50148 8008 50204
rect 8064 50148 8132 50204
rect 8188 50148 8256 50204
rect 8312 50148 8380 50204
rect 8436 50148 8504 50204
rect 8560 50148 8628 50204
rect 8684 50148 8752 50204
rect 8808 50148 8876 50204
rect 8932 50148 9000 50204
rect 9056 50148 9124 50204
rect 9180 50148 9248 50204
rect 9304 50148 9372 50204
rect 9428 50148 9496 50204
rect 9552 50148 9620 50204
rect 9676 50148 9744 50204
rect 9800 50148 10254 50204
rect 10310 50148 10378 50204
rect 10434 50148 10502 50204
rect 10558 50148 10626 50204
rect 10682 50148 10750 50204
rect 10806 50148 10874 50204
rect 10930 50148 10998 50204
rect 11054 50148 11122 50204
rect 11178 50148 11246 50204
rect 11302 50148 11370 50204
rect 11426 50148 11494 50204
rect 11550 50148 11618 50204
rect 11674 50148 11742 50204
rect 11798 50148 11866 50204
rect 11922 50148 11990 50204
rect 12046 50148 12114 50204
rect 12170 50148 12871 50204
rect 12927 50148 12995 50204
rect 13051 50148 13119 50204
rect 13175 50148 13243 50204
rect 13299 50148 13367 50204
rect 13423 50148 13491 50204
rect 13547 50148 13615 50204
rect 13671 50148 13739 50204
rect 13795 50148 13863 50204
rect 13919 50148 13987 50204
rect 14043 50148 14111 50204
rect 14167 50148 14235 50204
rect 14291 50148 14359 50204
rect 14415 50148 14483 50204
rect 14539 50148 14607 50204
rect 14663 50148 14839 50204
rect 139 50080 14839 50148
rect 139 50024 315 50080
rect 371 50024 439 50080
rect 495 50024 563 50080
rect 619 50024 687 50080
rect 743 50024 811 50080
rect 867 50024 935 50080
rect 991 50024 1059 50080
rect 1115 50024 1183 50080
rect 1239 50024 1307 50080
rect 1363 50024 1431 50080
rect 1487 50024 1555 50080
rect 1611 50024 1679 50080
rect 1735 50024 1803 50080
rect 1859 50024 1927 50080
rect 1983 50024 2051 50080
rect 2107 50024 2808 50080
rect 2864 50024 2932 50080
rect 2988 50024 3056 50080
rect 3112 50024 3180 50080
rect 3236 50024 3304 50080
rect 3360 50024 3428 50080
rect 3484 50024 3552 50080
rect 3608 50024 3676 50080
rect 3732 50024 3800 50080
rect 3856 50024 3924 50080
rect 3980 50024 4048 50080
rect 4104 50024 4172 50080
rect 4228 50024 4296 50080
rect 4352 50024 4420 50080
rect 4476 50024 4544 50080
rect 4600 50024 4668 50080
rect 4724 50024 5178 50080
rect 5234 50024 5302 50080
rect 5358 50024 5426 50080
rect 5482 50024 5550 50080
rect 5606 50024 5674 50080
rect 5730 50024 5798 50080
rect 5854 50024 5922 50080
rect 5978 50024 6046 50080
rect 6102 50024 6170 50080
rect 6226 50024 6294 50080
rect 6350 50024 6418 50080
rect 6474 50024 6542 50080
rect 6598 50024 6666 50080
rect 6722 50024 6790 50080
rect 6846 50024 6914 50080
rect 6970 50024 7038 50080
rect 7094 50024 7884 50080
rect 7940 50024 8008 50080
rect 8064 50024 8132 50080
rect 8188 50024 8256 50080
rect 8312 50024 8380 50080
rect 8436 50024 8504 50080
rect 8560 50024 8628 50080
rect 8684 50024 8752 50080
rect 8808 50024 8876 50080
rect 8932 50024 9000 50080
rect 9056 50024 9124 50080
rect 9180 50024 9248 50080
rect 9304 50024 9372 50080
rect 9428 50024 9496 50080
rect 9552 50024 9620 50080
rect 9676 50024 9744 50080
rect 9800 50024 10254 50080
rect 10310 50024 10378 50080
rect 10434 50024 10502 50080
rect 10558 50024 10626 50080
rect 10682 50024 10750 50080
rect 10806 50024 10874 50080
rect 10930 50024 10998 50080
rect 11054 50024 11122 50080
rect 11178 50024 11246 50080
rect 11302 50024 11370 50080
rect 11426 50024 11494 50080
rect 11550 50024 11618 50080
rect 11674 50024 11742 50080
rect 11798 50024 11866 50080
rect 11922 50024 11990 50080
rect 12046 50024 12114 50080
rect 12170 50024 12871 50080
rect 12927 50024 12995 50080
rect 13051 50024 13119 50080
rect 13175 50024 13243 50080
rect 13299 50024 13367 50080
rect 13423 50024 13491 50080
rect 13547 50024 13615 50080
rect 13671 50024 13739 50080
rect 13795 50024 13863 50080
rect 13919 50024 13987 50080
rect 14043 50024 14111 50080
rect 14167 50024 14235 50080
rect 14291 50024 14359 50080
rect 14415 50024 14483 50080
rect 14539 50024 14607 50080
rect 14663 50024 14839 50080
rect 139 49956 14839 50024
rect 139 49900 315 49956
rect 371 49900 439 49956
rect 495 49900 563 49956
rect 619 49900 687 49956
rect 743 49900 811 49956
rect 867 49900 935 49956
rect 991 49900 1059 49956
rect 1115 49900 1183 49956
rect 1239 49900 1307 49956
rect 1363 49900 1431 49956
rect 1487 49900 1555 49956
rect 1611 49900 1679 49956
rect 1735 49900 1803 49956
rect 1859 49900 1927 49956
rect 1983 49900 2051 49956
rect 2107 49900 2808 49956
rect 2864 49900 2932 49956
rect 2988 49900 3056 49956
rect 3112 49900 3180 49956
rect 3236 49900 3304 49956
rect 3360 49900 3428 49956
rect 3484 49900 3552 49956
rect 3608 49900 3676 49956
rect 3732 49900 3800 49956
rect 3856 49900 3924 49956
rect 3980 49900 4048 49956
rect 4104 49900 4172 49956
rect 4228 49900 4296 49956
rect 4352 49900 4420 49956
rect 4476 49900 4544 49956
rect 4600 49900 4668 49956
rect 4724 49900 5178 49956
rect 5234 49900 5302 49956
rect 5358 49900 5426 49956
rect 5482 49900 5550 49956
rect 5606 49900 5674 49956
rect 5730 49900 5798 49956
rect 5854 49900 5922 49956
rect 5978 49900 6046 49956
rect 6102 49900 6170 49956
rect 6226 49900 6294 49956
rect 6350 49900 6418 49956
rect 6474 49900 6542 49956
rect 6598 49900 6666 49956
rect 6722 49900 6790 49956
rect 6846 49900 6914 49956
rect 6970 49900 7038 49956
rect 7094 49900 7884 49956
rect 7940 49900 8008 49956
rect 8064 49900 8132 49956
rect 8188 49900 8256 49956
rect 8312 49900 8380 49956
rect 8436 49900 8504 49956
rect 8560 49900 8628 49956
rect 8684 49900 8752 49956
rect 8808 49900 8876 49956
rect 8932 49900 9000 49956
rect 9056 49900 9124 49956
rect 9180 49900 9248 49956
rect 9304 49900 9372 49956
rect 9428 49900 9496 49956
rect 9552 49900 9620 49956
rect 9676 49900 9744 49956
rect 9800 49900 10254 49956
rect 10310 49900 10378 49956
rect 10434 49900 10502 49956
rect 10558 49900 10626 49956
rect 10682 49900 10750 49956
rect 10806 49900 10874 49956
rect 10930 49900 10998 49956
rect 11054 49900 11122 49956
rect 11178 49900 11246 49956
rect 11302 49900 11370 49956
rect 11426 49900 11494 49956
rect 11550 49900 11618 49956
rect 11674 49900 11742 49956
rect 11798 49900 11866 49956
rect 11922 49900 11990 49956
rect 12046 49900 12114 49956
rect 12170 49900 12871 49956
rect 12927 49900 12995 49956
rect 13051 49900 13119 49956
rect 13175 49900 13243 49956
rect 13299 49900 13367 49956
rect 13423 49900 13491 49956
rect 13547 49900 13615 49956
rect 13671 49900 13739 49956
rect 13795 49900 13863 49956
rect 13919 49900 13987 49956
rect 14043 49900 14111 49956
rect 14167 49900 14235 49956
rect 14291 49900 14359 49956
rect 14415 49900 14483 49956
rect 14539 49900 14607 49956
rect 14663 49900 14839 49956
rect 139 49832 14839 49900
rect 139 49776 315 49832
rect 371 49776 439 49832
rect 495 49776 563 49832
rect 619 49776 687 49832
rect 743 49776 811 49832
rect 867 49776 935 49832
rect 991 49776 1059 49832
rect 1115 49776 1183 49832
rect 1239 49776 1307 49832
rect 1363 49776 1431 49832
rect 1487 49776 1555 49832
rect 1611 49776 1679 49832
rect 1735 49776 1803 49832
rect 1859 49776 1927 49832
rect 1983 49776 2051 49832
rect 2107 49776 2808 49832
rect 2864 49776 2932 49832
rect 2988 49776 3056 49832
rect 3112 49776 3180 49832
rect 3236 49776 3304 49832
rect 3360 49776 3428 49832
rect 3484 49776 3552 49832
rect 3608 49776 3676 49832
rect 3732 49776 3800 49832
rect 3856 49776 3924 49832
rect 3980 49776 4048 49832
rect 4104 49776 4172 49832
rect 4228 49776 4296 49832
rect 4352 49776 4420 49832
rect 4476 49776 4544 49832
rect 4600 49776 4668 49832
rect 4724 49776 5178 49832
rect 5234 49776 5302 49832
rect 5358 49776 5426 49832
rect 5482 49776 5550 49832
rect 5606 49776 5674 49832
rect 5730 49776 5798 49832
rect 5854 49776 5922 49832
rect 5978 49776 6046 49832
rect 6102 49776 6170 49832
rect 6226 49776 6294 49832
rect 6350 49776 6418 49832
rect 6474 49776 6542 49832
rect 6598 49776 6666 49832
rect 6722 49776 6790 49832
rect 6846 49776 6914 49832
rect 6970 49776 7038 49832
rect 7094 49776 7884 49832
rect 7940 49776 8008 49832
rect 8064 49776 8132 49832
rect 8188 49776 8256 49832
rect 8312 49776 8380 49832
rect 8436 49776 8504 49832
rect 8560 49776 8628 49832
rect 8684 49776 8752 49832
rect 8808 49776 8876 49832
rect 8932 49776 9000 49832
rect 9056 49776 9124 49832
rect 9180 49776 9248 49832
rect 9304 49776 9372 49832
rect 9428 49776 9496 49832
rect 9552 49776 9620 49832
rect 9676 49776 9744 49832
rect 9800 49776 10254 49832
rect 10310 49776 10378 49832
rect 10434 49776 10502 49832
rect 10558 49776 10626 49832
rect 10682 49776 10750 49832
rect 10806 49776 10874 49832
rect 10930 49776 10998 49832
rect 11054 49776 11122 49832
rect 11178 49776 11246 49832
rect 11302 49776 11370 49832
rect 11426 49776 11494 49832
rect 11550 49776 11618 49832
rect 11674 49776 11742 49832
rect 11798 49776 11866 49832
rect 11922 49776 11990 49832
rect 12046 49776 12114 49832
rect 12170 49776 12871 49832
rect 12927 49776 12995 49832
rect 13051 49776 13119 49832
rect 13175 49776 13243 49832
rect 13299 49776 13367 49832
rect 13423 49776 13491 49832
rect 13547 49776 13615 49832
rect 13671 49776 13739 49832
rect 13795 49776 13863 49832
rect 13919 49776 13987 49832
rect 14043 49776 14111 49832
rect 14167 49776 14235 49832
rect 14291 49776 14359 49832
rect 14415 49776 14483 49832
rect 14539 49776 14607 49832
rect 14663 49776 14839 49832
rect 139 49708 14839 49776
rect 139 49652 315 49708
rect 371 49652 439 49708
rect 495 49652 563 49708
rect 619 49652 687 49708
rect 743 49652 811 49708
rect 867 49652 935 49708
rect 991 49652 1059 49708
rect 1115 49652 1183 49708
rect 1239 49652 1307 49708
rect 1363 49652 1431 49708
rect 1487 49652 1555 49708
rect 1611 49652 1679 49708
rect 1735 49652 1803 49708
rect 1859 49652 1927 49708
rect 1983 49652 2051 49708
rect 2107 49652 2808 49708
rect 2864 49652 2932 49708
rect 2988 49652 3056 49708
rect 3112 49652 3180 49708
rect 3236 49652 3304 49708
rect 3360 49652 3428 49708
rect 3484 49652 3552 49708
rect 3608 49652 3676 49708
rect 3732 49652 3800 49708
rect 3856 49652 3924 49708
rect 3980 49652 4048 49708
rect 4104 49652 4172 49708
rect 4228 49652 4296 49708
rect 4352 49652 4420 49708
rect 4476 49652 4544 49708
rect 4600 49652 4668 49708
rect 4724 49652 5178 49708
rect 5234 49652 5302 49708
rect 5358 49652 5426 49708
rect 5482 49652 5550 49708
rect 5606 49652 5674 49708
rect 5730 49652 5798 49708
rect 5854 49652 5922 49708
rect 5978 49652 6046 49708
rect 6102 49652 6170 49708
rect 6226 49652 6294 49708
rect 6350 49652 6418 49708
rect 6474 49652 6542 49708
rect 6598 49652 6666 49708
rect 6722 49652 6790 49708
rect 6846 49652 6914 49708
rect 6970 49652 7038 49708
rect 7094 49652 7884 49708
rect 7940 49652 8008 49708
rect 8064 49652 8132 49708
rect 8188 49652 8256 49708
rect 8312 49652 8380 49708
rect 8436 49652 8504 49708
rect 8560 49652 8628 49708
rect 8684 49652 8752 49708
rect 8808 49652 8876 49708
rect 8932 49652 9000 49708
rect 9056 49652 9124 49708
rect 9180 49652 9248 49708
rect 9304 49652 9372 49708
rect 9428 49652 9496 49708
rect 9552 49652 9620 49708
rect 9676 49652 9744 49708
rect 9800 49652 10254 49708
rect 10310 49652 10378 49708
rect 10434 49652 10502 49708
rect 10558 49652 10626 49708
rect 10682 49652 10750 49708
rect 10806 49652 10874 49708
rect 10930 49652 10998 49708
rect 11054 49652 11122 49708
rect 11178 49652 11246 49708
rect 11302 49652 11370 49708
rect 11426 49652 11494 49708
rect 11550 49652 11618 49708
rect 11674 49652 11742 49708
rect 11798 49652 11866 49708
rect 11922 49652 11990 49708
rect 12046 49652 12114 49708
rect 12170 49652 12871 49708
rect 12927 49652 12995 49708
rect 13051 49652 13119 49708
rect 13175 49652 13243 49708
rect 13299 49652 13367 49708
rect 13423 49652 13491 49708
rect 13547 49652 13615 49708
rect 13671 49652 13739 49708
rect 13795 49652 13863 49708
rect 13919 49652 13987 49708
rect 14043 49652 14111 49708
rect 14167 49652 14235 49708
rect 14291 49652 14359 49708
rect 14415 49652 14483 49708
rect 14539 49652 14607 49708
rect 14663 49652 14839 49708
rect 139 49630 14839 49652
rect 2481 48042 2681 49358
rect 4851 48042 5051 49358
rect 7265 48042 7713 49358
rect 9927 48042 10127 49358
rect 12297 48042 12497 49358
rect 139 46430 14839 47780
rect 2481 44842 2681 46158
rect 4851 44842 5051 46158
rect 7265 44842 7713 46158
rect 9927 44842 10127 46158
rect 12297 44842 12497 46158
rect 305 43242 2117 44558
rect 2798 43242 4734 44558
rect 5168 43242 7104 44558
rect 7874 43242 9810 44558
rect 10244 43242 12180 44558
rect 12861 43242 14673 44558
rect 305 41642 2117 42958
rect 2798 41642 4734 42958
rect 5168 41642 7104 42958
rect 7874 41642 9810 42958
rect 10244 41642 12180 42958
rect 12861 41642 14673 42958
rect 309 41358 14669 41360
rect 305 40050 14673 41358
rect 305 40042 2117 40050
rect 2798 40042 4734 40050
rect 5168 40042 7104 40050
rect 7874 40042 9810 40050
rect 10244 40042 12180 40050
rect 12861 40042 14673 40050
rect 139 39748 14839 39780
rect 139 39692 315 39748
rect 371 39692 439 39748
rect 495 39692 563 39748
rect 619 39692 687 39748
rect 743 39692 811 39748
rect 867 39692 935 39748
rect 991 39692 1059 39748
rect 1115 39692 1183 39748
rect 1239 39692 1307 39748
rect 1363 39692 1431 39748
rect 1487 39692 1555 39748
rect 1611 39692 1679 39748
rect 1735 39692 1803 39748
rect 1859 39692 1927 39748
rect 1983 39692 2051 39748
rect 2107 39692 2808 39748
rect 2864 39692 2932 39748
rect 2988 39692 3056 39748
rect 3112 39692 3180 39748
rect 3236 39692 3304 39748
rect 3360 39692 3428 39748
rect 3484 39692 3552 39748
rect 3608 39692 3676 39748
rect 3732 39692 3800 39748
rect 3856 39692 3924 39748
rect 3980 39692 4048 39748
rect 4104 39692 4172 39748
rect 4228 39692 4296 39748
rect 4352 39692 4420 39748
rect 4476 39692 4544 39748
rect 4600 39692 4668 39748
rect 4724 39692 5178 39748
rect 5234 39692 5302 39748
rect 5358 39692 5426 39748
rect 5482 39692 5550 39748
rect 5606 39692 5674 39748
rect 5730 39692 5798 39748
rect 5854 39692 5922 39748
rect 5978 39692 6046 39748
rect 6102 39692 6170 39748
rect 6226 39692 6294 39748
rect 6350 39692 6418 39748
rect 6474 39692 6542 39748
rect 6598 39692 6666 39748
rect 6722 39692 6790 39748
rect 6846 39692 6914 39748
rect 6970 39692 7038 39748
rect 7094 39692 7884 39748
rect 7940 39692 8008 39748
rect 8064 39692 8132 39748
rect 8188 39692 8256 39748
rect 8312 39692 8380 39748
rect 8436 39692 8504 39748
rect 8560 39692 8628 39748
rect 8684 39692 8752 39748
rect 8808 39692 8876 39748
rect 8932 39692 9000 39748
rect 9056 39692 9124 39748
rect 9180 39692 9248 39748
rect 9304 39692 9372 39748
rect 9428 39692 9496 39748
rect 9552 39692 9620 39748
rect 9676 39692 9744 39748
rect 9800 39692 10254 39748
rect 10310 39692 10378 39748
rect 10434 39692 10502 39748
rect 10558 39692 10626 39748
rect 10682 39692 10750 39748
rect 10806 39692 10874 39748
rect 10930 39692 10998 39748
rect 11054 39692 11122 39748
rect 11178 39692 11246 39748
rect 11302 39692 11370 39748
rect 11426 39692 11494 39748
rect 11550 39692 11618 39748
rect 11674 39692 11742 39748
rect 11798 39692 11866 39748
rect 11922 39692 11990 39748
rect 12046 39692 12114 39748
rect 12170 39692 12871 39748
rect 12927 39692 12995 39748
rect 13051 39692 13119 39748
rect 13175 39692 13243 39748
rect 13299 39692 13367 39748
rect 13423 39692 13491 39748
rect 13547 39692 13615 39748
rect 13671 39692 13739 39748
rect 13795 39692 13863 39748
rect 13919 39692 13987 39748
rect 14043 39692 14111 39748
rect 14167 39692 14235 39748
rect 14291 39692 14359 39748
rect 14415 39692 14483 39748
rect 14539 39692 14607 39748
rect 14663 39692 14839 39748
rect 139 39624 14839 39692
rect 139 39568 315 39624
rect 371 39568 439 39624
rect 495 39568 563 39624
rect 619 39568 687 39624
rect 743 39568 811 39624
rect 867 39568 935 39624
rect 991 39568 1059 39624
rect 1115 39568 1183 39624
rect 1239 39568 1307 39624
rect 1363 39568 1431 39624
rect 1487 39568 1555 39624
rect 1611 39568 1679 39624
rect 1735 39568 1803 39624
rect 1859 39568 1927 39624
rect 1983 39568 2051 39624
rect 2107 39568 2808 39624
rect 2864 39568 2932 39624
rect 2988 39568 3056 39624
rect 3112 39568 3180 39624
rect 3236 39568 3304 39624
rect 3360 39568 3428 39624
rect 3484 39568 3552 39624
rect 3608 39568 3676 39624
rect 3732 39568 3800 39624
rect 3856 39568 3924 39624
rect 3980 39568 4048 39624
rect 4104 39568 4172 39624
rect 4228 39568 4296 39624
rect 4352 39568 4420 39624
rect 4476 39568 4544 39624
rect 4600 39568 4668 39624
rect 4724 39568 5178 39624
rect 5234 39568 5302 39624
rect 5358 39568 5426 39624
rect 5482 39568 5550 39624
rect 5606 39568 5674 39624
rect 5730 39568 5798 39624
rect 5854 39568 5922 39624
rect 5978 39568 6046 39624
rect 6102 39568 6170 39624
rect 6226 39568 6294 39624
rect 6350 39568 6418 39624
rect 6474 39568 6542 39624
rect 6598 39568 6666 39624
rect 6722 39568 6790 39624
rect 6846 39568 6914 39624
rect 6970 39568 7038 39624
rect 7094 39568 7884 39624
rect 7940 39568 8008 39624
rect 8064 39568 8132 39624
rect 8188 39568 8256 39624
rect 8312 39568 8380 39624
rect 8436 39568 8504 39624
rect 8560 39568 8628 39624
rect 8684 39568 8752 39624
rect 8808 39568 8876 39624
rect 8932 39568 9000 39624
rect 9056 39568 9124 39624
rect 9180 39568 9248 39624
rect 9304 39568 9372 39624
rect 9428 39568 9496 39624
rect 9552 39568 9620 39624
rect 9676 39568 9744 39624
rect 9800 39568 10254 39624
rect 10310 39568 10378 39624
rect 10434 39568 10502 39624
rect 10558 39568 10626 39624
rect 10682 39568 10750 39624
rect 10806 39568 10874 39624
rect 10930 39568 10998 39624
rect 11054 39568 11122 39624
rect 11178 39568 11246 39624
rect 11302 39568 11370 39624
rect 11426 39568 11494 39624
rect 11550 39568 11618 39624
rect 11674 39568 11742 39624
rect 11798 39568 11866 39624
rect 11922 39568 11990 39624
rect 12046 39568 12114 39624
rect 12170 39568 12871 39624
rect 12927 39568 12995 39624
rect 13051 39568 13119 39624
rect 13175 39568 13243 39624
rect 13299 39568 13367 39624
rect 13423 39568 13491 39624
rect 13547 39568 13615 39624
rect 13671 39568 13739 39624
rect 13795 39568 13863 39624
rect 13919 39568 13987 39624
rect 14043 39568 14111 39624
rect 14167 39568 14235 39624
rect 14291 39568 14359 39624
rect 14415 39568 14483 39624
rect 14539 39568 14607 39624
rect 14663 39568 14839 39624
rect 139 39500 14839 39568
rect 139 39444 315 39500
rect 371 39444 439 39500
rect 495 39444 563 39500
rect 619 39444 687 39500
rect 743 39444 811 39500
rect 867 39444 935 39500
rect 991 39444 1059 39500
rect 1115 39444 1183 39500
rect 1239 39444 1307 39500
rect 1363 39444 1431 39500
rect 1487 39444 1555 39500
rect 1611 39444 1679 39500
rect 1735 39444 1803 39500
rect 1859 39444 1927 39500
rect 1983 39444 2051 39500
rect 2107 39444 2808 39500
rect 2864 39444 2932 39500
rect 2988 39444 3056 39500
rect 3112 39444 3180 39500
rect 3236 39444 3304 39500
rect 3360 39444 3428 39500
rect 3484 39444 3552 39500
rect 3608 39444 3676 39500
rect 3732 39444 3800 39500
rect 3856 39444 3924 39500
rect 3980 39444 4048 39500
rect 4104 39444 4172 39500
rect 4228 39444 4296 39500
rect 4352 39444 4420 39500
rect 4476 39444 4544 39500
rect 4600 39444 4668 39500
rect 4724 39444 5178 39500
rect 5234 39444 5302 39500
rect 5358 39444 5426 39500
rect 5482 39444 5550 39500
rect 5606 39444 5674 39500
rect 5730 39444 5798 39500
rect 5854 39444 5922 39500
rect 5978 39444 6046 39500
rect 6102 39444 6170 39500
rect 6226 39444 6294 39500
rect 6350 39444 6418 39500
rect 6474 39444 6542 39500
rect 6598 39444 6666 39500
rect 6722 39444 6790 39500
rect 6846 39444 6914 39500
rect 6970 39444 7038 39500
rect 7094 39444 7884 39500
rect 7940 39444 8008 39500
rect 8064 39444 8132 39500
rect 8188 39444 8256 39500
rect 8312 39444 8380 39500
rect 8436 39444 8504 39500
rect 8560 39444 8628 39500
rect 8684 39444 8752 39500
rect 8808 39444 8876 39500
rect 8932 39444 9000 39500
rect 9056 39444 9124 39500
rect 9180 39444 9248 39500
rect 9304 39444 9372 39500
rect 9428 39444 9496 39500
rect 9552 39444 9620 39500
rect 9676 39444 9744 39500
rect 9800 39444 10254 39500
rect 10310 39444 10378 39500
rect 10434 39444 10502 39500
rect 10558 39444 10626 39500
rect 10682 39444 10750 39500
rect 10806 39444 10874 39500
rect 10930 39444 10998 39500
rect 11054 39444 11122 39500
rect 11178 39444 11246 39500
rect 11302 39444 11370 39500
rect 11426 39444 11494 39500
rect 11550 39444 11618 39500
rect 11674 39444 11742 39500
rect 11798 39444 11866 39500
rect 11922 39444 11990 39500
rect 12046 39444 12114 39500
rect 12170 39444 12871 39500
rect 12927 39444 12995 39500
rect 13051 39444 13119 39500
rect 13175 39444 13243 39500
rect 13299 39444 13367 39500
rect 13423 39444 13491 39500
rect 13547 39444 13615 39500
rect 13671 39444 13739 39500
rect 13795 39444 13863 39500
rect 13919 39444 13987 39500
rect 14043 39444 14111 39500
rect 14167 39444 14235 39500
rect 14291 39444 14359 39500
rect 14415 39444 14483 39500
rect 14539 39444 14607 39500
rect 14663 39444 14839 39500
rect 139 39376 14839 39444
rect 139 39320 315 39376
rect 371 39320 439 39376
rect 495 39320 563 39376
rect 619 39320 687 39376
rect 743 39320 811 39376
rect 867 39320 935 39376
rect 991 39320 1059 39376
rect 1115 39320 1183 39376
rect 1239 39320 1307 39376
rect 1363 39320 1431 39376
rect 1487 39320 1555 39376
rect 1611 39320 1679 39376
rect 1735 39320 1803 39376
rect 1859 39320 1927 39376
rect 1983 39320 2051 39376
rect 2107 39320 2808 39376
rect 2864 39320 2932 39376
rect 2988 39320 3056 39376
rect 3112 39320 3180 39376
rect 3236 39320 3304 39376
rect 3360 39320 3428 39376
rect 3484 39320 3552 39376
rect 3608 39320 3676 39376
rect 3732 39320 3800 39376
rect 3856 39320 3924 39376
rect 3980 39320 4048 39376
rect 4104 39320 4172 39376
rect 4228 39320 4296 39376
rect 4352 39320 4420 39376
rect 4476 39320 4544 39376
rect 4600 39320 4668 39376
rect 4724 39320 5178 39376
rect 5234 39320 5302 39376
rect 5358 39320 5426 39376
rect 5482 39320 5550 39376
rect 5606 39320 5674 39376
rect 5730 39320 5798 39376
rect 5854 39320 5922 39376
rect 5978 39320 6046 39376
rect 6102 39320 6170 39376
rect 6226 39320 6294 39376
rect 6350 39320 6418 39376
rect 6474 39320 6542 39376
rect 6598 39320 6666 39376
rect 6722 39320 6790 39376
rect 6846 39320 6914 39376
rect 6970 39320 7038 39376
rect 7094 39320 7884 39376
rect 7940 39320 8008 39376
rect 8064 39320 8132 39376
rect 8188 39320 8256 39376
rect 8312 39320 8380 39376
rect 8436 39320 8504 39376
rect 8560 39320 8628 39376
rect 8684 39320 8752 39376
rect 8808 39320 8876 39376
rect 8932 39320 9000 39376
rect 9056 39320 9124 39376
rect 9180 39320 9248 39376
rect 9304 39320 9372 39376
rect 9428 39320 9496 39376
rect 9552 39320 9620 39376
rect 9676 39320 9744 39376
rect 9800 39320 10254 39376
rect 10310 39320 10378 39376
rect 10434 39320 10502 39376
rect 10558 39320 10626 39376
rect 10682 39320 10750 39376
rect 10806 39320 10874 39376
rect 10930 39320 10998 39376
rect 11054 39320 11122 39376
rect 11178 39320 11246 39376
rect 11302 39320 11370 39376
rect 11426 39320 11494 39376
rect 11550 39320 11618 39376
rect 11674 39320 11742 39376
rect 11798 39320 11866 39376
rect 11922 39320 11990 39376
rect 12046 39320 12114 39376
rect 12170 39320 12871 39376
rect 12927 39320 12995 39376
rect 13051 39320 13119 39376
rect 13175 39320 13243 39376
rect 13299 39320 13367 39376
rect 13423 39320 13491 39376
rect 13547 39320 13615 39376
rect 13671 39320 13739 39376
rect 13795 39320 13863 39376
rect 13919 39320 13987 39376
rect 14043 39320 14111 39376
rect 14167 39320 14235 39376
rect 14291 39320 14359 39376
rect 14415 39320 14483 39376
rect 14539 39320 14607 39376
rect 14663 39320 14839 39376
rect 139 39252 14839 39320
rect 139 39196 315 39252
rect 371 39196 439 39252
rect 495 39196 563 39252
rect 619 39196 687 39252
rect 743 39196 811 39252
rect 867 39196 935 39252
rect 991 39196 1059 39252
rect 1115 39196 1183 39252
rect 1239 39196 1307 39252
rect 1363 39196 1431 39252
rect 1487 39196 1555 39252
rect 1611 39196 1679 39252
rect 1735 39196 1803 39252
rect 1859 39196 1927 39252
rect 1983 39196 2051 39252
rect 2107 39196 2808 39252
rect 2864 39196 2932 39252
rect 2988 39196 3056 39252
rect 3112 39196 3180 39252
rect 3236 39196 3304 39252
rect 3360 39196 3428 39252
rect 3484 39196 3552 39252
rect 3608 39196 3676 39252
rect 3732 39196 3800 39252
rect 3856 39196 3924 39252
rect 3980 39196 4048 39252
rect 4104 39196 4172 39252
rect 4228 39196 4296 39252
rect 4352 39196 4420 39252
rect 4476 39196 4544 39252
rect 4600 39196 4668 39252
rect 4724 39196 5178 39252
rect 5234 39196 5302 39252
rect 5358 39196 5426 39252
rect 5482 39196 5550 39252
rect 5606 39196 5674 39252
rect 5730 39196 5798 39252
rect 5854 39196 5922 39252
rect 5978 39196 6046 39252
rect 6102 39196 6170 39252
rect 6226 39196 6294 39252
rect 6350 39196 6418 39252
rect 6474 39196 6542 39252
rect 6598 39196 6666 39252
rect 6722 39196 6790 39252
rect 6846 39196 6914 39252
rect 6970 39196 7038 39252
rect 7094 39196 7884 39252
rect 7940 39196 8008 39252
rect 8064 39196 8132 39252
rect 8188 39196 8256 39252
rect 8312 39196 8380 39252
rect 8436 39196 8504 39252
rect 8560 39196 8628 39252
rect 8684 39196 8752 39252
rect 8808 39196 8876 39252
rect 8932 39196 9000 39252
rect 9056 39196 9124 39252
rect 9180 39196 9248 39252
rect 9304 39196 9372 39252
rect 9428 39196 9496 39252
rect 9552 39196 9620 39252
rect 9676 39196 9744 39252
rect 9800 39196 10254 39252
rect 10310 39196 10378 39252
rect 10434 39196 10502 39252
rect 10558 39196 10626 39252
rect 10682 39196 10750 39252
rect 10806 39196 10874 39252
rect 10930 39196 10998 39252
rect 11054 39196 11122 39252
rect 11178 39196 11246 39252
rect 11302 39196 11370 39252
rect 11426 39196 11494 39252
rect 11550 39196 11618 39252
rect 11674 39196 11742 39252
rect 11798 39196 11866 39252
rect 11922 39196 11990 39252
rect 12046 39196 12114 39252
rect 12170 39196 12871 39252
rect 12927 39196 12995 39252
rect 13051 39196 13119 39252
rect 13175 39196 13243 39252
rect 13299 39196 13367 39252
rect 13423 39196 13491 39252
rect 13547 39196 13615 39252
rect 13671 39196 13739 39252
rect 13795 39196 13863 39252
rect 13919 39196 13987 39252
rect 14043 39196 14111 39252
rect 14167 39196 14235 39252
rect 14291 39196 14359 39252
rect 14415 39196 14483 39252
rect 14539 39196 14607 39252
rect 14663 39196 14839 39252
rect 139 39128 14839 39196
rect 139 39072 315 39128
rect 371 39072 439 39128
rect 495 39072 563 39128
rect 619 39072 687 39128
rect 743 39072 811 39128
rect 867 39072 935 39128
rect 991 39072 1059 39128
rect 1115 39072 1183 39128
rect 1239 39072 1307 39128
rect 1363 39072 1431 39128
rect 1487 39072 1555 39128
rect 1611 39072 1679 39128
rect 1735 39072 1803 39128
rect 1859 39072 1927 39128
rect 1983 39072 2051 39128
rect 2107 39072 2808 39128
rect 2864 39072 2932 39128
rect 2988 39072 3056 39128
rect 3112 39072 3180 39128
rect 3236 39072 3304 39128
rect 3360 39072 3428 39128
rect 3484 39072 3552 39128
rect 3608 39072 3676 39128
rect 3732 39072 3800 39128
rect 3856 39072 3924 39128
rect 3980 39072 4048 39128
rect 4104 39072 4172 39128
rect 4228 39072 4296 39128
rect 4352 39072 4420 39128
rect 4476 39072 4544 39128
rect 4600 39072 4668 39128
rect 4724 39072 5178 39128
rect 5234 39072 5302 39128
rect 5358 39072 5426 39128
rect 5482 39072 5550 39128
rect 5606 39072 5674 39128
rect 5730 39072 5798 39128
rect 5854 39072 5922 39128
rect 5978 39072 6046 39128
rect 6102 39072 6170 39128
rect 6226 39072 6294 39128
rect 6350 39072 6418 39128
rect 6474 39072 6542 39128
rect 6598 39072 6666 39128
rect 6722 39072 6790 39128
rect 6846 39072 6914 39128
rect 6970 39072 7038 39128
rect 7094 39072 7884 39128
rect 7940 39072 8008 39128
rect 8064 39072 8132 39128
rect 8188 39072 8256 39128
rect 8312 39072 8380 39128
rect 8436 39072 8504 39128
rect 8560 39072 8628 39128
rect 8684 39072 8752 39128
rect 8808 39072 8876 39128
rect 8932 39072 9000 39128
rect 9056 39072 9124 39128
rect 9180 39072 9248 39128
rect 9304 39072 9372 39128
rect 9428 39072 9496 39128
rect 9552 39072 9620 39128
rect 9676 39072 9744 39128
rect 9800 39072 10254 39128
rect 10310 39072 10378 39128
rect 10434 39072 10502 39128
rect 10558 39072 10626 39128
rect 10682 39072 10750 39128
rect 10806 39072 10874 39128
rect 10930 39072 10998 39128
rect 11054 39072 11122 39128
rect 11178 39072 11246 39128
rect 11302 39072 11370 39128
rect 11426 39072 11494 39128
rect 11550 39072 11618 39128
rect 11674 39072 11742 39128
rect 11798 39072 11866 39128
rect 11922 39072 11990 39128
rect 12046 39072 12114 39128
rect 12170 39072 12871 39128
rect 12927 39072 12995 39128
rect 13051 39072 13119 39128
rect 13175 39072 13243 39128
rect 13299 39072 13367 39128
rect 13423 39072 13491 39128
rect 13547 39072 13615 39128
rect 13671 39072 13739 39128
rect 13795 39072 13863 39128
rect 13919 39072 13987 39128
rect 14043 39072 14111 39128
rect 14167 39072 14235 39128
rect 14291 39072 14359 39128
rect 14415 39072 14483 39128
rect 14539 39072 14607 39128
rect 14663 39072 14839 39128
rect 139 39004 14839 39072
rect 139 38948 315 39004
rect 371 38948 439 39004
rect 495 38948 563 39004
rect 619 38948 687 39004
rect 743 38948 811 39004
rect 867 38948 935 39004
rect 991 38948 1059 39004
rect 1115 38948 1183 39004
rect 1239 38948 1307 39004
rect 1363 38948 1431 39004
rect 1487 38948 1555 39004
rect 1611 38948 1679 39004
rect 1735 38948 1803 39004
rect 1859 38948 1927 39004
rect 1983 38948 2051 39004
rect 2107 38948 2808 39004
rect 2864 38948 2932 39004
rect 2988 38948 3056 39004
rect 3112 38948 3180 39004
rect 3236 38948 3304 39004
rect 3360 38948 3428 39004
rect 3484 38948 3552 39004
rect 3608 38948 3676 39004
rect 3732 38948 3800 39004
rect 3856 38948 3924 39004
rect 3980 38948 4048 39004
rect 4104 38948 4172 39004
rect 4228 38948 4296 39004
rect 4352 38948 4420 39004
rect 4476 38948 4544 39004
rect 4600 38948 4668 39004
rect 4724 38948 5178 39004
rect 5234 38948 5302 39004
rect 5358 38948 5426 39004
rect 5482 38948 5550 39004
rect 5606 38948 5674 39004
rect 5730 38948 5798 39004
rect 5854 38948 5922 39004
rect 5978 38948 6046 39004
rect 6102 38948 6170 39004
rect 6226 38948 6294 39004
rect 6350 38948 6418 39004
rect 6474 38948 6542 39004
rect 6598 38948 6666 39004
rect 6722 38948 6790 39004
rect 6846 38948 6914 39004
rect 6970 38948 7038 39004
rect 7094 38948 7884 39004
rect 7940 38948 8008 39004
rect 8064 38948 8132 39004
rect 8188 38948 8256 39004
rect 8312 38948 8380 39004
rect 8436 38948 8504 39004
rect 8560 38948 8628 39004
rect 8684 38948 8752 39004
rect 8808 38948 8876 39004
rect 8932 38948 9000 39004
rect 9056 38948 9124 39004
rect 9180 38948 9248 39004
rect 9304 38948 9372 39004
rect 9428 38948 9496 39004
rect 9552 38948 9620 39004
rect 9676 38948 9744 39004
rect 9800 38948 10254 39004
rect 10310 38948 10378 39004
rect 10434 38948 10502 39004
rect 10558 38948 10626 39004
rect 10682 38948 10750 39004
rect 10806 38948 10874 39004
rect 10930 38948 10998 39004
rect 11054 38948 11122 39004
rect 11178 38948 11246 39004
rect 11302 38948 11370 39004
rect 11426 38948 11494 39004
rect 11550 38948 11618 39004
rect 11674 38948 11742 39004
rect 11798 38948 11866 39004
rect 11922 38948 11990 39004
rect 12046 38948 12114 39004
rect 12170 38948 12871 39004
rect 12927 38948 12995 39004
rect 13051 38948 13119 39004
rect 13175 38948 13243 39004
rect 13299 38948 13367 39004
rect 13423 38948 13491 39004
rect 13547 38948 13615 39004
rect 13671 38948 13739 39004
rect 13795 38948 13863 39004
rect 13919 38948 13987 39004
rect 14043 38948 14111 39004
rect 14167 38948 14235 39004
rect 14291 38948 14359 39004
rect 14415 38948 14483 39004
rect 14539 38948 14607 39004
rect 14663 38948 14839 39004
rect 139 38880 14839 38948
rect 139 38824 315 38880
rect 371 38824 439 38880
rect 495 38824 563 38880
rect 619 38824 687 38880
rect 743 38824 811 38880
rect 867 38824 935 38880
rect 991 38824 1059 38880
rect 1115 38824 1183 38880
rect 1239 38824 1307 38880
rect 1363 38824 1431 38880
rect 1487 38824 1555 38880
rect 1611 38824 1679 38880
rect 1735 38824 1803 38880
rect 1859 38824 1927 38880
rect 1983 38824 2051 38880
rect 2107 38824 2808 38880
rect 2864 38824 2932 38880
rect 2988 38824 3056 38880
rect 3112 38824 3180 38880
rect 3236 38824 3304 38880
rect 3360 38824 3428 38880
rect 3484 38824 3552 38880
rect 3608 38824 3676 38880
rect 3732 38824 3800 38880
rect 3856 38824 3924 38880
rect 3980 38824 4048 38880
rect 4104 38824 4172 38880
rect 4228 38824 4296 38880
rect 4352 38824 4420 38880
rect 4476 38824 4544 38880
rect 4600 38824 4668 38880
rect 4724 38824 5178 38880
rect 5234 38824 5302 38880
rect 5358 38824 5426 38880
rect 5482 38824 5550 38880
rect 5606 38824 5674 38880
rect 5730 38824 5798 38880
rect 5854 38824 5922 38880
rect 5978 38824 6046 38880
rect 6102 38824 6170 38880
rect 6226 38824 6294 38880
rect 6350 38824 6418 38880
rect 6474 38824 6542 38880
rect 6598 38824 6666 38880
rect 6722 38824 6790 38880
rect 6846 38824 6914 38880
rect 6970 38824 7038 38880
rect 7094 38824 7884 38880
rect 7940 38824 8008 38880
rect 8064 38824 8132 38880
rect 8188 38824 8256 38880
rect 8312 38824 8380 38880
rect 8436 38824 8504 38880
rect 8560 38824 8628 38880
rect 8684 38824 8752 38880
rect 8808 38824 8876 38880
rect 8932 38824 9000 38880
rect 9056 38824 9124 38880
rect 9180 38824 9248 38880
rect 9304 38824 9372 38880
rect 9428 38824 9496 38880
rect 9552 38824 9620 38880
rect 9676 38824 9744 38880
rect 9800 38824 10254 38880
rect 10310 38824 10378 38880
rect 10434 38824 10502 38880
rect 10558 38824 10626 38880
rect 10682 38824 10750 38880
rect 10806 38824 10874 38880
rect 10930 38824 10998 38880
rect 11054 38824 11122 38880
rect 11178 38824 11246 38880
rect 11302 38824 11370 38880
rect 11426 38824 11494 38880
rect 11550 38824 11618 38880
rect 11674 38824 11742 38880
rect 11798 38824 11866 38880
rect 11922 38824 11990 38880
rect 12046 38824 12114 38880
rect 12170 38824 12871 38880
rect 12927 38824 12995 38880
rect 13051 38824 13119 38880
rect 13175 38824 13243 38880
rect 13299 38824 13367 38880
rect 13423 38824 13491 38880
rect 13547 38824 13615 38880
rect 13671 38824 13739 38880
rect 13795 38824 13863 38880
rect 13919 38824 13987 38880
rect 14043 38824 14111 38880
rect 14167 38824 14235 38880
rect 14291 38824 14359 38880
rect 14415 38824 14483 38880
rect 14539 38824 14607 38880
rect 14663 38824 14839 38880
rect 139 38756 14839 38824
rect 139 38700 315 38756
rect 371 38700 439 38756
rect 495 38700 563 38756
rect 619 38700 687 38756
rect 743 38700 811 38756
rect 867 38700 935 38756
rect 991 38700 1059 38756
rect 1115 38700 1183 38756
rect 1239 38700 1307 38756
rect 1363 38700 1431 38756
rect 1487 38700 1555 38756
rect 1611 38700 1679 38756
rect 1735 38700 1803 38756
rect 1859 38700 1927 38756
rect 1983 38700 2051 38756
rect 2107 38700 2808 38756
rect 2864 38700 2932 38756
rect 2988 38700 3056 38756
rect 3112 38700 3180 38756
rect 3236 38700 3304 38756
rect 3360 38700 3428 38756
rect 3484 38700 3552 38756
rect 3608 38700 3676 38756
rect 3732 38700 3800 38756
rect 3856 38700 3924 38756
rect 3980 38700 4048 38756
rect 4104 38700 4172 38756
rect 4228 38700 4296 38756
rect 4352 38700 4420 38756
rect 4476 38700 4544 38756
rect 4600 38700 4668 38756
rect 4724 38700 5178 38756
rect 5234 38700 5302 38756
rect 5358 38700 5426 38756
rect 5482 38700 5550 38756
rect 5606 38700 5674 38756
rect 5730 38700 5798 38756
rect 5854 38700 5922 38756
rect 5978 38700 6046 38756
rect 6102 38700 6170 38756
rect 6226 38700 6294 38756
rect 6350 38700 6418 38756
rect 6474 38700 6542 38756
rect 6598 38700 6666 38756
rect 6722 38700 6790 38756
rect 6846 38700 6914 38756
rect 6970 38700 7038 38756
rect 7094 38700 7884 38756
rect 7940 38700 8008 38756
rect 8064 38700 8132 38756
rect 8188 38700 8256 38756
rect 8312 38700 8380 38756
rect 8436 38700 8504 38756
rect 8560 38700 8628 38756
rect 8684 38700 8752 38756
rect 8808 38700 8876 38756
rect 8932 38700 9000 38756
rect 9056 38700 9124 38756
rect 9180 38700 9248 38756
rect 9304 38700 9372 38756
rect 9428 38700 9496 38756
rect 9552 38700 9620 38756
rect 9676 38700 9744 38756
rect 9800 38700 10254 38756
rect 10310 38700 10378 38756
rect 10434 38700 10502 38756
rect 10558 38700 10626 38756
rect 10682 38700 10750 38756
rect 10806 38700 10874 38756
rect 10930 38700 10998 38756
rect 11054 38700 11122 38756
rect 11178 38700 11246 38756
rect 11302 38700 11370 38756
rect 11426 38700 11494 38756
rect 11550 38700 11618 38756
rect 11674 38700 11742 38756
rect 11798 38700 11866 38756
rect 11922 38700 11990 38756
rect 12046 38700 12114 38756
rect 12170 38700 12871 38756
rect 12927 38700 12995 38756
rect 13051 38700 13119 38756
rect 13175 38700 13243 38756
rect 13299 38700 13367 38756
rect 13423 38700 13491 38756
rect 13547 38700 13615 38756
rect 13671 38700 13739 38756
rect 13795 38700 13863 38756
rect 13919 38700 13987 38756
rect 14043 38700 14111 38756
rect 14167 38700 14235 38756
rect 14291 38700 14359 38756
rect 14415 38700 14483 38756
rect 14539 38700 14607 38756
rect 14663 38700 14839 38756
rect 139 38632 14839 38700
rect 139 38576 315 38632
rect 371 38576 439 38632
rect 495 38576 563 38632
rect 619 38576 687 38632
rect 743 38576 811 38632
rect 867 38576 935 38632
rect 991 38576 1059 38632
rect 1115 38576 1183 38632
rect 1239 38576 1307 38632
rect 1363 38576 1431 38632
rect 1487 38576 1555 38632
rect 1611 38576 1679 38632
rect 1735 38576 1803 38632
rect 1859 38576 1927 38632
rect 1983 38576 2051 38632
rect 2107 38576 2808 38632
rect 2864 38576 2932 38632
rect 2988 38576 3056 38632
rect 3112 38576 3180 38632
rect 3236 38576 3304 38632
rect 3360 38576 3428 38632
rect 3484 38576 3552 38632
rect 3608 38576 3676 38632
rect 3732 38576 3800 38632
rect 3856 38576 3924 38632
rect 3980 38576 4048 38632
rect 4104 38576 4172 38632
rect 4228 38576 4296 38632
rect 4352 38576 4420 38632
rect 4476 38576 4544 38632
rect 4600 38576 4668 38632
rect 4724 38576 5178 38632
rect 5234 38576 5302 38632
rect 5358 38576 5426 38632
rect 5482 38576 5550 38632
rect 5606 38576 5674 38632
rect 5730 38576 5798 38632
rect 5854 38576 5922 38632
rect 5978 38576 6046 38632
rect 6102 38576 6170 38632
rect 6226 38576 6294 38632
rect 6350 38576 6418 38632
rect 6474 38576 6542 38632
rect 6598 38576 6666 38632
rect 6722 38576 6790 38632
rect 6846 38576 6914 38632
rect 6970 38576 7038 38632
rect 7094 38576 7884 38632
rect 7940 38576 8008 38632
rect 8064 38576 8132 38632
rect 8188 38576 8256 38632
rect 8312 38576 8380 38632
rect 8436 38576 8504 38632
rect 8560 38576 8628 38632
rect 8684 38576 8752 38632
rect 8808 38576 8876 38632
rect 8932 38576 9000 38632
rect 9056 38576 9124 38632
rect 9180 38576 9248 38632
rect 9304 38576 9372 38632
rect 9428 38576 9496 38632
rect 9552 38576 9620 38632
rect 9676 38576 9744 38632
rect 9800 38576 10254 38632
rect 10310 38576 10378 38632
rect 10434 38576 10502 38632
rect 10558 38576 10626 38632
rect 10682 38576 10750 38632
rect 10806 38576 10874 38632
rect 10930 38576 10998 38632
rect 11054 38576 11122 38632
rect 11178 38576 11246 38632
rect 11302 38576 11370 38632
rect 11426 38576 11494 38632
rect 11550 38576 11618 38632
rect 11674 38576 11742 38632
rect 11798 38576 11866 38632
rect 11922 38576 11990 38632
rect 12046 38576 12114 38632
rect 12170 38576 12871 38632
rect 12927 38576 12995 38632
rect 13051 38576 13119 38632
rect 13175 38576 13243 38632
rect 13299 38576 13367 38632
rect 13423 38576 13491 38632
rect 13547 38576 13615 38632
rect 13671 38576 13739 38632
rect 13795 38576 13863 38632
rect 13919 38576 13987 38632
rect 14043 38576 14111 38632
rect 14167 38576 14235 38632
rect 14291 38576 14359 38632
rect 14415 38576 14483 38632
rect 14539 38576 14607 38632
rect 14663 38576 14839 38632
rect 139 38508 14839 38576
rect 139 38452 315 38508
rect 371 38452 439 38508
rect 495 38452 563 38508
rect 619 38452 687 38508
rect 743 38452 811 38508
rect 867 38452 935 38508
rect 991 38452 1059 38508
rect 1115 38452 1183 38508
rect 1239 38452 1307 38508
rect 1363 38452 1431 38508
rect 1487 38452 1555 38508
rect 1611 38452 1679 38508
rect 1735 38452 1803 38508
rect 1859 38452 1927 38508
rect 1983 38452 2051 38508
rect 2107 38452 2808 38508
rect 2864 38452 2932 38508
rect 2988 38452 3056 38508
rect 3112 38452 3180 38508
rect 3236 38452 3304 38508
rect 3360 38452 3428 38508
rect 3484 38452 3552 38508
rect 3608 38452 3676 38508
rect 3732 38452 3800 38508
rect 3856 38452 3924 38508
rect 3980 38452 4048 38508
rect 4104 38452 4172 38508
rect 4228 38452 4296 38508
rect 4352 38452 4420 38508
rect 4476 38452 4544 38508
rect 4600 38452 4668 38508
rect 4724 38452 5178 38508
rect 5234 38452 5302 38508
rect 5358 38452 5426 38508
rect 5482 38452 5550 38508
rect 5606 38452 5674 38508
rect 5730 38452 5798 38508
rect 5854 38452 5922 38508
rect 5978 38452 6046 38508
rect 6102 38452 6170 38508
rect 6226 38452 6294 38508
rect 6350 38452 6418 38508
rect 6474 38452 6542 38508
rect 6598 38452 6666 38508
rect 6722 38452 6790 38508
rect 6846 38452 6914 38508
rect 6970 38452 7038 38508
rect 7094 38452 7884 38508
rect 7940 38452 8008 38508
rect 8064 38452 8132 38508
rect 8188 38452 8256 38508
rect 8312 38452 8380 38508
rect 8436 38452 8504 38508
rect 8560 38452 8628 38508
rect 8684 38452 8752 38508
rect 8808 38452 8876 38508
rect 8932 38452 9000 38508
rect 9056 38452 9124 38508
rect 9180 38452 9248 38508
rect 9304 38452 9372 38508
rect 9428 38452 9496 38508
rect 9552 38452 9620 38508
rect 9676 38452 9744 38508
rect 9800 38452 10254 38508
rect 10310 38452 10378 38508
rect 10434 38452 10502 38508
rect 10558 38452 10626 38508
rect 10682 38452 10750 38508
rect 10806 38452 10874 38508
rect 10930 38452 10998 38508
rect 11054 38452 11122 38508
rect 11178 38452 11246 38508
rect 11302 38452 11370 38508
rect 11426 38452 11494 38508
rect 11550 38452 11618 38508
rect 11674 38452 11742 38508
rect 11798 38452 11866 38508
rect 11922 38452 11990 38508
rect 12046 38452 12114 38508
rect 12170 38452 12871 38508
rect 12927 38452 12995 38508
rect 13051 38452 13119 38508
rect 13175 38452 13243 38508
rect 13299 38452 13367 38508
rect 13423 38452 13491 38508
rect 13547 38452 13615 38508
rect 13671 38452 13739 38508
rect 13795 38452 13863 38508
rect 13919 38452 13987 38508
rect 14043 38452 14111 38508
rect 14167 38452 14235 38508
rect 14291 38452 14359 38508
rect 14415 38452 14483 38508
rect 14539 38452 14607 38508
rect 14663 38452 14839 38508
rect 139 38430 14839 38452
rect 10 38176 86 38186
rect 10 36824 20 38176
rect 76 38160 86 38176
rect 14892 38176 14968 38186
rect 14892 38160 14902 38176
rect 76 38154 14902 38160
rect 76 38135 2491 38154
rect 76 38079 2289 38135
rect 2345 38098 2491 38135
rect 2547 38098 2615 38154
rect 2671 38098 4861 38154
rect 4917 38098 4985 38154
rect 5041 38098 7275 38154
rect 7331 38098 7399 38154
rect 7455 38098 7523 38154
rect 7579 38098 7647 38154
rect 7703 38098 9937 38154
rect 9993 38098 10061 38154
rect 10117 38098 12307 38154
rect 12363 38098 12431 38154
rect 12487 38098 14902 38154
rect 2345 38079 14902 38098
rect 76 38030 14902 38079
rect 76 38003 2491 38030
rect 76 37947 2289 38003
rect 2345 37974 2491 38003
rect 2547 37974 2615 38030
rect 2671 37974 4861 38030
rect 4917 37974 4985 38030
rect 5041 37974 7275 38030
rect 7331 37974 7399 38030
rect 7455 37974 7523 38030
rect 7579 37974 7647 38030
rect 7703 37974 9937 38030
rect 9993 37974 10061 38030
rect 10117 37974 12307 38030
rect 12363 37974 12431 38030
rect 12487 37974 14902 38030
rect 2345 37947 14902 37974
rect 76 37906 14902 37947
rect 76 37871 2491 37906
rect 76 37815 2289 37871
rect 2345 37850 2491 37871
rect 2547 37850 2615 37906
rect 2671 37850 4861 37906
rect 4917 37850 4985 37906
rect 5041 37850 7275 37906
rect 7331 37850 7399 37906
rect 7455 37850 7523 37906
rect 7579 37850 7647 37906
rect 7703 37850 9937 37906
rect 9993 37850 10061 37906
rect 10117 37850 12307 37906
rect 12363 37850 12431 37906
rect 12487 37850 14902 37906
rect 2345 37815 14902 37850
rect 76 37782 14902 37815
rect 76 37739 2491 37782
rect 76 37683 2289 37739
rect 2345 37726 2491 37739
rect 2547 37726 2615 37782
rect 2671 37726 4861 37782
rect 4917 37726 4985 37782
rect 5041 37726 7275 37782
rect 7331 37726 7399 37782
rect 7455 37726 7523 37782
rect 7579 37726 7647 37782
rect 7703 37726 9937 37782
rect 9993 37726 10061 37782
rect 10117 37726 12307 37782
rect 12363 37726 12431 37782
rect 12487 37726 14902 37782
rect 2345 37683 14902 37726
rect 76 37658 14902 37683
rect 76 37607 2491 37658
rect 76 37551 2289 37607
rect 2345 37602 2491 37607
rect 2547 37602 2615 37658
rect 2671 37602 4861 37658
rect 4917 37602 4985 37658
rect 5041 37602 7275 37658
rect 7331 37602 7399 37658
rect 7455 37602 7523 37658
rect 7579 37602 7647 37658
rect 7703 37602 9937 37658
rect 9993 37602 10061 37658
rect 10117 37602 12307 37658
rect 12363 37602 12431 37658
rect 12487 37602 14902 37658
rect 2345 37551 14902 37602
rect 76 37534 14902 37551
rect 76 37478 2491 37534
rect 2547 37478 2615 37534
rect 2671 37478 4861 37534
rect 4917 37478 4985 37534
rect 5041 37478 7275 37534
rect 7331 37478 7399 37534
rect 7455 37478 7523 37534
rect 7579 37478 7647 37534
rect 7703 37478 9937 37534
rect 9993 37478 10061 37534
rect 10117 37478 12307 37534
rect 12363 37478 12431 37534
rect 12487 37478 14902 37534
rect 76 37475 14902 37478
rect 76 37419 2289 37475
rect 2345 37419 14902 37475
rect 76 37410 14902 37419
rect 76 37354 2491 37410
rect 2547 37354 2615 37410
rect 2671 37354 4861 37410
rect 4917 37354 4985 37410
rect 5041 37354 7275 37410
rect 7331 37354 7399 37410
rect 7455 37354 7523 37410
rect 7579 37354 7647 37410
rect 7703 37354 9937 37410
rect 9993 37354 10061 37410
rect 10117 37354 12307 37410
rect 12363 37354 12431 37410
rect 12487 37354 14902 37410
rect 76 37343 14902 37354
rect 76 37287 2289 37343
rect 2345 37287 14902 37343
rect 76 37286 14902 37287
rect 76 37230 2491 37286
rect 2547 37230 2615 37286
rect 2671 37230 4861 37286
rect 4917 37230 4985 37286
rect 5041 37230 7275 37286
rect 7331 37230 7399 37286
rect 7455 37230 7523 37286
rect 7579 37230 7647 37286
rect 7703 37230 9937 37286
rect 9993 37230 10061 37286
rect 10117 37230 12307 37286
rect 12363 37230 12431 37286
rect 12487 37230 14902 37286
rect 76 37211 14902 37230
rect 76 37155 2289 37211
rect 2345 37162 14902 37211
rect 2345 37155 2491 37162
rect 76 37106 2491 37155
rect 2547 37106 2615 37162
rect 2671 37106 4861 37162
rect 4917 37106 4985 37162
rect 5041 37106 7275 37162
rect 7331 37106 7399 37162
rect 7455 37106 7523 37162
rect 7579 37106 7647 37162
rect 7703 37106 9937 37162
rect 9993 37106 10061 37162
rect 10117 37106 12307 37162
rect 12363 37106 12431 37162
rect 12487 37106 14902 37162
rect 76 37079 14902 37106
rect 76 37023 2289 37079
rect 2345 37038 14902 37079
rect 2345 37023 2491 37038
rect 76 36982 2491 37023
rect 2547 36982 2615 37038
rect 2671 36982 4861 37038
rect 4917 36982 4985 37038
rect 5041 36982 7275 37038
rect 7331 36982 7399 37038
rect 7455 36982 7523 37038
rect 7579 36982 7647 37038
rect 7703 36982 9937 37038
rect 9993 36982 10061 37038
rect 10117 36982 12307 37038
rect 12363 36982 12431 37038
rect 12487 36982 14902 37038
rect 76 36947 14902 36982
rect 76 36891 2289 36947
rect 2345 36914 14902 36947
rect 2345 36891 2491 36914
rect 76 36858 2491 36891
rect 2547 36858 2615 36914
rect 2671 36858 4861 36914
rect 4917 36858 4985 36914
rect 5041 36858 7275 36914
rect 7331 36858 7399 36914
rect 7455 36858 7523 36914
rect 7579 36858 7647 36914
rect 7703 36858 9937 36914
rect 9993 36858 10061 36914
rect 10117 36858 12307 36914
rect 12363 36858 12431 36914
rect 12487 36858 14902 36914
rect 76 36850 14902 36858
rect 76 36824 86 36850
rect 10 36814 86 36824
rect 14892 36824 14902 36850
rect 14958 36824 14968 38176
rect 14892 36814 14968 36824
rect 2481 33636 2681 36564
rect 4851 33636 5051 36564
rect 7265 33636 7713 36564
rect 9927 33636 10127 36564
rect 12297 33636 12497 36564
rect 305 30436 2117 33364
rect 2798 30436 4734 33364
rect 5168 30436 7104 33364
rect 7874 30436 9810 33364
rect 10244 30436 12180 33364
rect 12861 30436 14673 33364
rect 305 28842 2117 30158
rect 2798 28842 4734 30158
rect 5168 28842 7104 30158
rect 7874 28842 9810 30158
rect 10244 28842 12180 30158
rect 12861 28842 14673 30158
rect 2481 27242 2681 28558
rect 4851 27242 5051 28558
rect 7265 27242 7713 28558
rect 9927 27242 10127 28558
rect 12297 27242 12497 28558
rect 305 24036 2117 26964
rect 2798 24036 4734 26964
rect 5168 24036 7104 26964
rect 7874 24036 9810 26964
rect 10244 24036 12180 26964
rect 12861 24036 14673 26964
rect 305 20836 2117 23764
rect 2798 20836 4734 23764
rect 5168 20836 7104 23764
rect 7874 20836 9810 23764
rect 10244 20836 12180 23764
rect 12861 20836 14673 23764
rect 305 17636 2117 20564
rect 2798 17636 4734 20564
rect 5168 17636 7104 20564
rect 7874 17636 9810 20564
rect 10244 17636 12180 20564
rect 12861 17636 14673 20564
rect 305 14436 2117 17364
rect 2798 14436 4734 17364
rect 5168 14436 7104 17364
rect 7874 14436 9810 17364
rect 10244 14436 12180 17364
rect 12861 14436 14673 17364
rect 2481 12842 2681 14158
rect 4851 12842 5051 14158
rect 7265 12842 7713 14158
rect 9927 12842 10127 14158
rect 12297 12842 12497 14158
rect 305 11242 2117 12558
rect 2798 11242 4734 12558
rect 5168 11242 7104 12558
rect 7874 11242 9810 12558
rect 10244 11242 12180 12558
rect 12861 11242 14673 12558
rect 2481 8036 2681 10964
rect 4851 8036 5051 10964
rect 7265 8036 7713 10964
rect 9927 8036 10127 10964
rect 12297 8036 12497 10964
rect 2481 4836 2681 7764
rect 4851 4836 5051 7764
rect 7265 4836 7713 7764
rect 9927 4836 10127 7764
rect 12297 4836 12497 7764
rect 2481 1636 2681 4564
rect 4851 1636 5051 4564
rect 7265 1636 7713 4564
rect 9927 1636 10127 4564
rect 12297 1636 12497 4564
use comp018green_esd_clamp_v5p0_DVDD  comp018green_esd_clamp_v5p0_DVDD_0
timestamp 1758727423
transform 1 0 1008 0 1 1147
box -747 -51 13709 46134
<< labels >>
rlabel metal3 s 705 6432 705 6432 4 DVSS
port 1 nsew
rlabel metal3 s 752 3261 752 3261 4 DVSS
port 1 nsew
rlabel metal3 s 774 9418 774 9418 4 DVSS
port 1 nsew
rlabel metal3 s 774 13611 774 13611 4 DVSS
port 1 nsew
rlabel metal3 s 774 11795 774 11795 4 DVDD
port 2 nsew
rlabel metal3 s 774 22234 774 22234 4 DVDD
port 2 nsew
rlabel metal3 s 774 19120 774 19120 4 DVDD
port 2 nsew
rlabel metal3 s 774 15905 774 15905 4 DVDD
port 2 nsew
rlabel metal3 s 774 27853 774 27853 4 DVSS
port 1 nsew
rlabel metal3 s 774 29488 774 29488 4 DVDD
port 2 nsew
rlabel metal3 s 774 25470 774 25470 4 DVDD
port 2 nsew
rlabel metal3 s 774 35106 774 35106 4 DVSS
port 1 nsew
rlabel metal3 s 774 31879 774 31879 4 DVDD
port 2 nsew
rlabel metal3 s 774 45369 774 45369 4 DVSS
port 1 nsew
rlabel metal3 s 774 43934 774 43934 4 DVDD
port 2 nsew
rlabel metal3 s 774 42169 774 42169 4 DVDD
port 2 nsew
rlabel metal3 s 774 40734 774 40734 4 DVDD
port 2 nsew
rlabel metal3 s 774 48569 774 48569 4 DVSS
port 1 nsew
rlabel metal3 s 774 53534 774 53534 4 DVSS
port 1 nsew
rlabel metal3 s 774 56560 774 56560 4 DVSS
port 1 nsew
rlabel metal3 s 774 54969 774 54969 4 DVDD
port 2 nsew
rlabel metal3 s 774 47134 774 47134 4 DVDD
port 2 nsew
rlabel metal3 s 774 50334 774 50334 4 VDD
port 3 nsew
rlabel metal3 s 774 39134 774 39134 4 VDD
port 3 nsew
rlabel metal3 s 774 37534 774 37534 4 VSS
port 4 nsew
<< end >>
