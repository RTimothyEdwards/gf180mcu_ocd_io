magic
tech gf180mcuD
magscale 1 10
timestamp 1758818392
<< metal2 >>
rect 272 69800 2172 70000
rect 2752 69800 4802 70000
rect 5122 69800 7172 70000
rect 7828 69800 9878 70000
rect 10198 69800 12248 70000
rect 12828 69800 14728 70000
<< metal5 >>
rect 0 68400 1000 69678
rect 14000 68400 15000 69678
rect 0 66800 1000 68200
rect 14000 66800 15000 68200
rect 0 65200 1000 66600
rect 14000 65200 15000 66600
rect 0 63600 1000 65000
rect 14000 63600 15000 65000
rect 0 62000 1000 63400
rect 14000 62000 15000 63400
rect 0 60400 1000 61800
rect 14000 60400 15000 61800
rect 0 58800 1000 60200
rect 14000 58800 15000 60200
rect 0 57200 1000 58600
rect 14000 57200 15000 58600
rect 0 55600 1000 57000
rect 14000 55600 15000 57000
rect 0 54000 1000 55400
rect 14000 54000 15000 55400
rect 0 52400 1000 53800
rect 14000 52400 15000 53800
rect 0 50800 1000 52200
rect 14000 50800 15000 52200
rect 0 49200 1000 50600
rect 14000 49200 15000 50600
rect 0 46000 1000 49000
rect 14000 46000 15000 49000
rect 0 42800 1000 45800
rect 14000 42800 15000 45800
rect 0 41200 1000 42600
rect 14000 41200 15000 42600
rect 0 39600 1000 41000
rect 14000 39600 15000 41000
rect 0 36400 1000 39400
rect 14000 36400 15000 39400
rect 0 33200 1000 36200
rect 14000 33200 15000 36200
rect 0 30000 1000 33000
rect 14000 30000 15000 33000
rect 0 26800 1000 29800
rect 14000 26800 15000 29800
rect 0 25200 1000 26600
rect 14000 25200 15000 26600
rect 0 23600 1000 25000
rect 14000 23600 15000 25000
rect 0 20400 1000 23400
rect 14000 20400 15000 23400
rect 0 17200 1000 20200
rect 14000 17200 15000 20200
rect 0 14000 1000 17000
rect 14000 14000 15000 17000
rect 1500 400 13500 12400
use 5LM_METAL_RAIL_PAD_60  5LM_METAL_RAIL_PAD_60_0
timestamp 1586916644
transform 1 0 0 0 1 0
box -32 0 15032 69968
use GF_NI_DVDD_BASE  GF_NI_DVDD_BASE_0
timestamp 1758741431
transform 1 0 11 0 1 12400
box -11 0 14989 57600
<< labels >>
flabel metal5 s 0 17200 1000 20200 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 0 14000 1000 17000 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 0 46000 1000 49000 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 0 39600 1000 41000 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 0 25200 1000 26600 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 0 20400 1000 23400 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 0 57200 1000 58600 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 0 60400 1000 61800 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 0 65200 1000 66600 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 0 68400 1000 69678 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 0 49200 1000 50600 0 FreeSans 1600 0 0 0 VSS
port 3 nsew ground bidirectional
flabel metal5 s 0 63600 1000 65000 0 FreeSans 1600 0 0 0 VSS
port 3 nsew ground bidirectional
flabel metal5 s 0 66800 1000 68200 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 0 58800 1000 60200 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 0 55600 1000 57000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 0 54000 1000 55400 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 0 52400 1000 53800 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 0 41200 1000 42600 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 0 42800 1000 45800 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 0 36400 1000 39400 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 0 33200 1000 36200 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 0 30000 1000 33000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 0 26800 1000 29800 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 0 23600 1000 25000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 1500 400 13500 12400 0 FreeSans 8000 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal2 s 272 69800 2172 70000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal2 s 2752 69800 4802 70000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal2 s 5122 69800 7172 70000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal2 s 7828 69800 9878 70000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal2 s 10198 69800 12248 70000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal2 s 12828 69800 14728 70000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 0 62000 1000 63400 0 FreeSans 1600 0 0 0 VDD
port 6 nsew power bidirectional
flabel metal5 s 0 50800 1000 52200 0 FreeSans 1600 0 0 0 VDD
port 6 nsew power bidirectional
flabel metal5 s 14000 17200 15000 20200 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 14000 14000 15000 17000 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 14000 46000 15000 49000 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 14000 39600 15000 41000 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 14000 25200 15000 26600 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 14000 20400 15000 23400 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 14000 57200 15000 58600 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 14000 60400 15000 61800 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 14000 65200 15000 66600 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 14000 68400 15000 69678 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal5 s 14000 49200 15000 50600 0 FreeSans 1600 0 0 0 VSS
port 3 nsew ground bidirectional
flabel metal5 s 14000 63600 15000 65000 0 FreeSans 1600 0 0 0 VSS
port 3 nsew ground bidirectional
flabel metal5 s 14000 66800 15000 68200 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 14000 58800 15000 60200 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 14000 55600 15000 57000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 14000 54000 15000 55400 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 14000 52400 15000 53800 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 14000 41200 15000 42600 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 14000 42800 15000 45800 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 14000 36400 15000 39400 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 14000 33200 15000 36200 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 14000 30000 15000 33000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 14000 26800 15000 29800 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 14000 23600 15000 25000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal5 s 14000 62000 15000 63400 0 FreeSans 1600 0 0 0 VDD
port 6 nsew power bidirectional
flabel metal5 s 14000 50800 15000 52200 0 FreeSans 1600 0 0 0 VDD
port 6 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 70000
string LEFclass PAD POWER
string LEFsymmetry X Y R90
string LEFsite GF_IO_Site
<< end >>
