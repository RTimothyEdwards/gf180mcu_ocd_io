magic
tech gf180mcuD
magscale 1 10
timestamp 1758722869
<< checkpaint >>
rect -2756 54700 -1466 56453
<< nwell >>
rect -2756 54700 -1466 56453
<< nsubdiff >>
rect -2673 56348 -1549 56370
rect -2673 56302 -2651 56348
rect -2135 56302 -1805 56348
rect -1571 56302 -1549 56348
rect -2673 56280 -1549 56302
rect -2673 56194 -2583 56280
rect -2673 54926 -2651 56194
rect -2605 54926 -2583 56194
rect -1639 56194 -1549 56280
rect -1639 55960 -1617 56194
rect -1571 55960 -1549 56194
rect -1639 55724 -1549 55960
rect -1639 55208 -1617 55724
rect -1571 55208 -1549 55724
rect -2673 54840 -2583 54926
rect -1639 54972 -1549 55208
rect -1639 54926 -1617 54972
rect -1571 54926 -1549 54972
rect -1639 54840 -1549 54926
rect -2673 54818 -1549 54840
rect -2673 54772 -2651 54818
rect -1571 54772 -1549 54818
rect -2673 54750 -1549 54772
<< nsubdiffcont >>
rect -2651 56302 -2135 56348
rect -1805 56302 -1571 56348
rect -2651 54926 -2605 56194
rect -1617 55960 -1571 56194
rect -1617 55208 -1571 55724
rect -1617 54926 -1571 54972
rect -2651 54772 -1571 54818
<< polysilicon >>
rect -2331 56032 -2171 56045
rect -2331 55986 -2274 56032
rect -2228 55986 -2171 56032
rect -2331 55943 -2171 55986
rect -2331 55120 -2171 55163
rect -2331 55074 -2274 55120
rect -2228 55074 -2171 55120
rect -2331 55061 -2171 55074
rect -2051 56032 -1891 56045
rect -2051 55986 -1994 56032
rect -1948 55986 -1891 56032
rect -2051 55943 -1891 55986
rect -2051 55120 -1891 55163
rect -2051 55074 -1994 55120
rect -1948 55074 -1891 55120
rect -2051 55061 -1891 55074
<< polycontact >>
rect -2274 55986 -2228 56032
rect -2274 55074 -2228 55120
rect -1994 55986 -1948 56032
rect -1994 55074 -1948 55120
<< ppolyres >>
rect -2331 55163 -2171 55943
rect -2051 55163 -1891 55943
<< metal1 >>
rect -2662 56348 -2111 56359
rect -2662 56302 -2651 56348
rect -2135 56302 -2111 56348
rect -2662 56291 -2111 56302
rect -2662 56194 -2594 56291
rect -2662 54926 -2651 56194
rect -2605 55131 -2594 56194
rect -2329 56032 -2173 56043
rect -2329 55986 -2274 56032
rect -2228 55986 -2173 56032
rect -2329 55975 -2173 55986
rect -2049 56032 -1893 56430
rect -1837 56348 -1560 56359
rect -1837 56302 -1805 56348
rect -1571 56302 -1560 56348
rect -1837 56291 -1560 56302
rect -2049 55986 -1994 56032
rect -1948 55986 -1893 56032
rect -2049 55975 -1893 55986
rect -1628 56194 -1560 56291
rect -2249 55885 -2173 55975
rect -1628 55960 -1617 56194
rect -1571 55960 -1560 56194
rect -1628 55945 -1560 55960
rect -2249 55809 -1480 55885
rect -1628 55724 -1560 55749
rect -1628 55208 -1617 55724
rect -1571 55208 -1560 55724
rect -1628 55180 -1560 55208
rect -2605 55120 -2173 55131
rect -2605 55074 -2274 55120
rect -2228 55074 -2173 55120
rect -2605 55063 -2173 55074
rect -2049 55120 -1480 55131
rect -2049 55074 -1994 55120
rect -1948 55074 -1480 55120
rect -2049 55063 -1480 55074
rect -2605 54926 -2594 55063
rect -2662 54829 -2594 54926
rect -1628 54972 -1560 55005
rect -1628 54926 -1617 54972
rect -1571 54926 -1560 54972
rect -1628 54829 -1560 54926
rect -2730 54818 -1480 54829
rect -2730 54772 -2651 54818
rect -1571 54772 -1480 54818
rect -2730 54700 -1480 54772
<< end >>
