magic
tech gf180mcuD
magscale 1 10
timestamp 1758724778
<< nwell >>
rect 0 -878 12382 14423
<< psubdiff >>
rect -975 15239 13355 15294
rect -975 15234 1290 15239
rect -975 14588 -953 15234
rect 793 14593 1290 15234
rect 2236 15238 13355 15239
rect 2236 15235 6604 15238
rect 2236 15233 4828 15235
rect 2236 14593 3060 15233
rect 793 14588 3060 14593
rect -975 14587 3060 14588
rect 4006 14589 4828 15233
rect 5774 14592 6604 15235
rect 7550 15227 13355 15238
rect 7550 14592 8368 15227
rect 5774 14589 8368 14592
rect 4006 14587 8368 14589
rect -975 14581 8368 14587
rect 9314 15214 11487 15227
rect 9314 14581 10141 15214
rect -975 14568 10141 14581
rect 11087 14581 11487 15214
rect 13333 14581 13355 15227
rect 11087 14568 13355 14581
rect -975 14516 13355 14568
rect -975 14501 12455 14516
rect -975 14481 -53 14501
rect -975 -865 -953 14481
rect -907 -865 -849 14481
rect -803 -865 -745 14481
rect -699 -865 -641 14481
rect -595 -865 -537 14481
rect -491 -865 -433 14481
rect -387 -865 -329 14481
rect -283 -865 -225 14481
rect -179 -865 -121 14481
rect -75 -865 -53 14481
rect -975 -910 -53 -865
rect 12433 -830 12455 14501
rect 12501 -830 12559 14516
rect 12605 -830 12663 14516
rect 12709 -830 12767 14516
rect 12813 -830 12871 14516
rect 12917 -830 12975 14516
rect 13021 -830 13079 14516
rect 13125 -830 13183 14516
rect 13229 -830 13287 14516
rect 13333 -830 13355 14516
rect 12433 -910 13355 -830
rect -975 -932 13355 -910
rect -975 -978 -913 -932
rect 13333 -978 13355 -932
rect -975 -1036 13355 -978
rect -975 -1082 -913 -1036
rect 13333 -1082 13355 -1036
rect -975 -1140 13355 -1082
rect -975 -1186 -913 -1140
rect 13333 -1186 13355 -1140
rect -975 -1244 13355 -1186
rect -975 -1290 -913 -1244
rect 13333 -1290 13355 -1244
rect -975 -1312 13355 -1290
<< nsubdiff >>
rect 96 14279 12299 14340
rect 96 13933 118 14279
rect 864 13933 11531 14279
rect 12277 13933 12299 14279
rect 96 13818 12299 13933
rect 96 272 183 13818
rect 429 12926 11953 13818
rect 429 272 451 12926
rect 96 54 451 272
rect 11931 272 11953 12926
rect 12199 272 12299 13818
rect 11931 250 12299 272
rect 11959 54 12299 250
rect 96 32 12299 54
rect 96 -714 118 32
rect 12264 -714 12299 32
rect 96 -736 12299 -714
<< psubdiffcont >>
rect -953 14588 793 15234
rect 1290 14593 2236 15239
rect 3060 14587 4006 15233
rect 4828 14589 5774 15235
rect 6604 14592 7550 15238
rect 8368 14581 9314 15227
rect 10141 14568 11087 15214
rect 11487 14581 13333 15227
rect -953 -865 -907 14481
rect -849 -865 -803 14481
rect -745 -865 -699 14481
rect -641 -865 -595 14481
rect -537 -865 -491 14481
rect -433 -865 -387 14481
rect -329 -865 -283 14481
rect -225 -865 -179 14481
rect -121 -865 -75 14481
rect 12455 -830 12501 14516
rect 12559 -830 12605 14516
rect 12663 -830 12709 14516
rect 12767 -830 12813 14516
rect 12871 -830 12917 14516
rect 12975 -830 13021 14516
rect 13079 -830 13125 14516
rect 13183 -830 13229 14516
rect 13287 -830 13333 14516
rect -913 -978 13333 -932
rect -913 -1082 13333 -1036
rect -913 -1186 13333 -1140
rect -913 -1290 13333 -1244
<< nsubdiffcont >>
rect 118 13933 864 14279
rect 11531 13933 12277 14279
rect 183 272 429 13818
rect 11953 272 12199 13818
rect 118 -714 12264 32
<< polysilicon >>
rect 974 12667 1185 12686
rect 974 12621 1009 12667
rect 1149 12621 1185 12667
rect 974 12602 1185 12621
rect 2360 12667 2571 12686
rect 2360 12621 2395 12667
rect 2535 12621 2571 12667
rect 2360 12602 2571 12621
rect 2746 12667 2957 12686
rect 2746 12621 2781 12667
rect 2921 12621 2957 12667
rect 2746 12602 2957 12621
rect 4120 12667 4331 12686
rect 4120 12621 4155 12667
rect 4295 12621 4331 12667
rect 4120 12602 4331 12621
rect 4511 12667 4722 12686
rect 4511 12621 4541 12667
rect 4681 12621 4722 12667
rect 4511 12602 4722 12621
rect 5892 12667 6103 12686
rect 5892 12621 5927 12667
rect 6067 12621 6103 12667
rect 5892 12602 6103 12621
rect 6280 12667 6491 12686
rect 6280 12621 6315 12667
rect 6455 12621 6491 12667
rect 6280 12602 6491 12621
rect 7662 12667 7873 12686
rect 7662 12621 7701 12667
rect 7841 12621 7873 12667
rect 7662 12602 7873 12621
rect 8049 12667 8260 12686
rect 8049 12621 8087 12667
rect 8227 12621 8260 12667
rect 8049 12602 8260 12621
rect 9428 12667 9639 12686
rect 9428 12621 9461 12667
rect 9601 12621 9639 12667
rect 9428 12602 9639 12621
rect 9815 12667 10026 12686
rect 9815 12621 9847 12667
rect 9987 12621 10026 12667
rect 9815 12602 10026 12621
rect 11201 12667 11412 12686
rect 11201 12621 11233 12667
rect 11373 12621 11412 12667
rect 11201 12602 11412 12621
rect 974 387 1185 406
rect 974 341 1009 387
rect 1149 341 1185 387
rect 974 322 1185 341
rect 2360 387 2571 406
rect 2360 341 2395 387
rect 2535 341 2571 387
rect 2360 322 2571 341
rect 2746 387 2957 406
rect 2746 341 2781 387
rect 2921 341 2957 387
rect 2746 322 2957 341
rect 4120 387 4331 406
rect 4120 341 4155 387
rect 4295 341 4331 387
rect 4120 322 4331 341
rect 4511 387 4722 406
rect 4511 341 4546 387
rect 4686 341 4722 387
rect 4511 322 4722 341
rect 5892 387 6103 406
rect 5892 341 5927 387
rect 6067 341 6103 387
rect 5892 322 6103 341
rect 6280 387 6491 406
rect 6280 341 6315 387
rect 6455 341 6491 387
rect 6280 322 6491 341
rect 7662 387 7873 406
rect 7662 341 7697 387
rect 7837 341 7873 387
rect 7662 322 7873 341
rect 8049 387 8260 406
rect 8049 341 8084 387
rect 8224 341 8260 387
rect 8049 322 8260 341
rect 9428 387 9639 406
rect 9428 341 9463 387
rect 9603 341 9639 387
rect 9428 322 9639 341
rect 9815 387 10026 406
rect 9815 341 9850 387
rect 9990 341 10026 387
rect 9815 322 10026 341
rect 11201 387 11412 406
rect 11201 341 11236 387
rect 11376 341 11412 387
rect 11201 322 11412 341
<< polycontact >>
rect 1009 12621 1149 12667
rect 2395 12621 2535 12667
rect 2781 12621 2921 12667
rect 4155 12621 4295 12667
rect 4541 12621 4681 12667
rect 5927 12621 6067 12667
rect 6315 12621 6455 12667
rect 7701 12621 7841 12667
rect 8087 12621 8227 12667
rect 9461 12621 9601 12667
rect 9847 12621 9987 12667
rect 11233 12621 11373 12667
rect 1009 341 1149 387
rect 2395 341 2535 387
rect 2781 341 2921 387
rect 4155 341 4295 387
rect 4546 341 4686 387
rect 5927 341 6067 387
rect 6315 341 6455 387
rect 7697 341 7837 387
rect 8084 341 8224 387
rect 9463 341 9603 387
rect 9850 341 9990 387
rect 11236 341 11376 387
<< metal1 >>
rect -964 15234 804 15245
rect -964 14588 -953 15234
rect 793 14588 804 15234
rect -964 14577 804 14588
rect 1279 15239 2247 15250
rect 1279 14593 1290 15239
rect 2236 14593 2247 15239
rect 1279 14582 2247 14593
rect 3049 15233 4017 15244
rect 3049 14587 3060 15233
rect 4006 14587 4017 15233
rect -964 14481 -64 14577
rect 3049 14576 4017 14587
rect 4817 15235 5785 15246
rect 4817 14589 4828 15235
rect 5774 14589 5785 15235
rect 4817 14578 5785 14589
rect 6593 15238 7561 15249
rect 6593 14592 6604 15238
rect 7550 14592 7561 15238
rect 6593 14581 7561 14592
rect 8357 15227 9325 15238
rect 8357 14581 8368 15227
rect 9314 14581 9325 15227
rect 11476 15227 13344 15238
rect 8357 14570 9325 14581
rect 10130 15214 11098 15225
rect 10130 14568 10141 15214
rect 11087 14568 11098 15214
rect 11476 14782 11487 15227
rect 11468 14770 11487 14782
rect 11468 14718 11480 14770
rect 11468 14662 11487 14718
rect 11468 14610 11480 14662
rect 11468 14598 11487 14610
rect 11476 14581 11487 14598
rect 13333 14581 13344 15227
rect 11476 14570 13344 14581
rect 10130 14557 11098 14568
rect -964 -865 -953 14481
rect -907 -865 -849 14481
rect -803 -865 -745 14481
rect -699 -865 -641 14481
rect -595 -865 -537 14481
rect -491 -865 -433 14481
rect -387 -865 -329 14481
rect -283 -865 -225 14481
rect -179 -865 -121 14481
rect -75 -865 -64 14481
rect 12444 14516 13344 14570
rect 107 14279 875 14290
rect 107 13933 118 14279
rect 864 13933 875 14279
rect 107 13922 875 13933
rect 11520 14279 12288 14290
rect 11520 13933 11531 14279
rect 12277 13933 12288 14279
rect 11520 13922 12288 13933
rect 107 13829 765 13922
rect 172 13818 765 13829
rect 172 546 183 13818
rect 107 272 183 546
rect 429 13120 765 13818
rect 429 10260 467 13120
rect 727 10260 765 13120
rect 11617 13818 12288 13922
rect 11617 13437 11953 13818
rect 998 12667 1160 12678
rect 998 12621 1009 12667
rect 1149 12621 1160 12667
rect 998 12610 1160 12621
rect 2384 12667 2546 12678
rect 2384 12621 2395 12667
rect 2535 12621 2546 12667
rect 2384 12610 2546 12621
rect 2770 12667 2932 12678
rect 2770 12621 2781 12667
rect 2921 12621 2932 12667
rect 2770 12610 2932 12621
rect 4144 12667 4306 12678
rect 4144 12621 4155 12667
rect 4295 12621 4306 12667
rect 4144 12610 4306 12621
rect 4530 12667 4692 12678
rect 4530 12621 4541 12667
rect 4681 12621 4692 12667
rect 4530 12610 4692 12621
rect 5916 12667 6078 12678
rect 5916 12621 5927 12667
rect 6067 12621 6078 12667
rect 5916 12610 6078 12621
rect 6304 12667 6466 12678
rect 6304 12621 6315 12667
rect 6455 12621 6466 12667
rect 6304 12610 6466 12621
rect 7690 12667 7852 12678
rect 7690 12621 7701 12667
rect 7841 12621 7852 12667
rect 7690 12610 7852 12621
rect 8076 12667 8238 12678
rect 8076 12621 8087 12667
rect 8227 12621 8238 12667
rect 8076 12610 8238 12621
rect 9450 12667 9612 12678
rect 9450 12621 9461 12667
rect 9601 12621 9612 12667
rect 9450 12610 9612 12621
rect 9836 12667 9998 12678
rect 9836 12621 9847 12667
rect 9987 12621 9998 12667
rect 9836 12610 9998 12621
rect 11222 12667 11384 12678
rect 11222 12621 11233 12667
rect 11373 12621 11384 12667
rect 11222 12610 11384 12621
rect 429 9920 765 10260
rect 429 7060 467 9920
rect 727 7060 765 9920
rect 429 6720 765 7060
rect 429 3860 467 6720
rect 727 3860 765 6720
rect 429 3535 765 3860
rect 429 675 467 3535
rect 727 675 765 3535
rect 429 496 765 675
rect 429 272 475 496
rect 1055 398 1101 12610
rect 2441 398 2487 12610
rect 2823 398 2869 12610
rect 4209 398 4255 12610
rect 4591 398 4637 12610
rect 5977 398 6023 12610
rect 6359 398 6405 12610
rect 7745 398 7791 12610
rect 8127 398 8173 12610
rect 9513 398 9559 12610
rect 9895 398 9941 12610
rect 11281 398 11327 12610
rect 11617 10265 11682 13437
rect 11942 10265 11953 13437
rect 11617 9915 11953 10265
rect 11617 7055 11682 9915
rect 11942 7055 11953 9915
rect 11617 6715 11953 7055
rect 11617 3855 11682 6715
rect 11942 3855 11953 6715
rect 11617 3515 11953 3855
rect 11617 655 11682 3515
rect 11942 655 11953 3515
rect 11617 497 11953 655
rect 998 387 1160 398
rect 998 341 1009 387
rect 1149 341 1160 387
rect 998 330 1160 341
rect 2384 387 2546 398
rect 2384 341 2395 387
rect 2535 341 2546 387
rect 2384 330 2546 341
rect 2770 387 2932 398
rect 2770 341 2781 387
rect 2921 341 2932 387
rect 2770 330 2932 341
rect 4144 387 4306 398
rect 4144 341 4155 387
rect 4295 341 4306 387
rect 4144 330 4306 341
rect 4535 387 4697 398
rect 4535 341 4546 387
rect 4686 341 4697 387
rect 4535 330 4697 341
rect 5916 387 6078 398
rect 5916 341 5927 387
rect 6067 341 6078 387
rect 5916 330 6078 341
rect 6304 387 6466 398
rect 6304 341 6315 387
rect 6455 341 6466 387
rect 6304 330 6466 341
rect 7686 387 7848 398
rect 7686 341 7697 387
rect 7837 341 7848 387
rect 7686 330 7848 341
rect 8073 387 8235 398
rect 8073 341 8084 387
rect 8224 341 8235 387
rect 8073 330 8235 341
rect 9452 387 9614 398
rect 9452 341 9463 387
rect 9603 341 9614 387
rect 9452 330 9614 341
rect 9839 387 10001 398
rect 9839 341 9850 387
rect 9990 341 10001 387
rect 9839 330 10001 341
rect 11225 387 11387 398
rect 11225 341 11236 387
rect 11376 341 11387 387
rect 11225 330 11387 341
rect 107 43 475 272
rect 11920 272 11953 497
rect 12199 272 12288 13818
rect 11920 43 12288 272
rect 107 32 12288 43
rect 107 -714 118 32
rect 12264 -714 12288 32
rect 107 -725 12288 -714
rect -964 -921 -64 -865
rect 12444 -830 12455 14516
rect 12501 -830 12559 14516
rect 12605 -830 12663 14516
rect 12709 -830 12767 14516
rect 12813 -830 12871 14516
rect 12917 -830 12975 14516
rect 13021 -830 13079 14516
rect 13125 -830 13183 14516
rect 13229 -830 13287 14516
rect 13333 -830 13344 14516
rect 12444 -921 13344 -830
rect -964 -932 13344 -921
rect -964 -978 -913 -932
rect 13333 -978 13344 -932
rect -964 -1036 13344 -978
rect -964 -1082 -913 -1036
rect 13333 -1082 13344 -1036
rect -964 -1140 13344 -1082
rect -964 -1186 -913 -1140
rect 13333 -1186 13344 -1140
rect -964 -1244 13344 -1186
rect -964 -1290 -913 -1244
rect 13333 -1290 13344 -1244
rect -964 -1301 13344 -1290
<< via1 >>
rect -719 14707 -667 14759
rect -611 14707 -559 14759
rect -503 14707 -451 14759
rect 524 14718 576 14770
rect 632 14718 684 14770
rect 740 14718 792 14770
rect -719 14599 -667 14651
rect -611 14599 -559 14651
rect -503 14599 -451 14651
rect 524 14610 576 14662
rect 632 14610 684 14662
rect 740 14610 792 14662
rect 1309 14718 1361 14770
rect 1417 14718 1469 14770
rect 1525 14718 1577 14770
rect 1633 14718 1685 14770
rect 1741 14718 1793 14770
rect 1849 14718 1901 14770
rect 1957 14718 2009 14770
rect 2065 14718 2117 14770
rect 2173 14718 2225 14770
rect 1309 14610 1361 14662
rect 1417 14610 1469 14662
rect 1525 14610 1577 14662
rect 1633 14610 1685 14662
rect 1741 14610 1793 14662
rect 1849 14610 1901 14662
rect 1957 14610 2009 14662
rect 2065 14610 2117 14662
rect 2173 14610 2225 14662
rect 3076 14718 3128 14770
rect 3184 14718 3236 14770
rect 3292 14718 3344 14770
rect 3400 14718 3452 14770
rect 3508 14718 3560 14770
rect 3616 14718 3668 14770
rect 3724 14718 3776 14770
rect 3832 14718 3884 14770
rect 3940 14718 3992 14770
rect 3076 14610 3128 14662
rect 3184 14610 3236 14662
rect 3292 14610 3344 14662
rect 3400 14610 3452 14662
rect 3508 14610 3560 14662
rect 3616 14610 3668 14662
rect 3724 14610 3776 14662
rect 3832 14610 3884 14662
rect 3940 14610 3992 14662
rect 4843 14718 4895 14770
rect 4951 14718 5003 14770
rect 5059 14718 5111 14770
rect 5167 14718 5219 14770
rect 5275 14718 5327 14770
rect 5383 14718 5435 14770
rect 5491 14718 5543 14770
rect 5599 14718 5651 14770
rect 5707 14718 5759 14770
rect 4843 14610 4895 14662
rect 4951 14610 5003 14662
rect 5059 14610 5111 14662
rect 5167 14610 5219 14662
rect 5275 14610 5327 14662
rect 5383 14610 5435 14662
rect 5491 14610 5543 14662
rect 5599 14610 5651 14662
rect 5707 14610 5759 14662
rect 6617 14718 6669 14770
rect 6725 14718 6777 14770
rect 6833 14718 6885 14770
rect 6941 14718 6993 14770
rect 7049 14718 7101 14770
rect 7157 14718 7209 14770
rect 7265 14718 7317 14770
rect 7373 14718 7425 14770
rect 7481 14718 7533 14770
rect 6617 14610 6669 14662
rect 6725 14610 6777 14662
rect 6833 14610 6885 14662
rect 6941 14610 6993 14662
rect 7049 14610 7101 14662
rect 7157 14610 7209 14662
rect 7265 14610 7317 14662
rect 7373 14610 7425 14662
rect 7481 14610 7533 14662
rect 8381 14718 8433 14770
rect 8489 14718 8541 14770
rect 8597 14718 8649 14770
rect 8705 14718 8757 14770
rect 8813 14718 8865 14770
rect 8921 14718 8973 14770
rect 9029 14718 9081 14770
rect 9137 14718 9189 14770
rect 9245 14718 9297 14770
rect 8381 14610 8433 14662
rect 8489 14610 8541 14662
rect 8597 14610 8649 14662
rect 8705 14610 8757 14662
rect 8813 14610 8865 14662
rect 8921 14610 8973 14662
rect 9029 14610 9081 14662
rect 9137 14610 9189 14662
rect 9245 14610 9297 14662
rect 10151 14718 10203 14770
rect 10259 14718 10311 14770
rect 10367 14718 10419 14770
rect 10475 14718 10527 14770
rect 10583 14718 10635 14770
rect 10691 14718 10743 14770
rect 10799 14718 10851 14770
rect 10907 14718 10959 14770
rect 11015 14718 11067 14770
rect 10151 14610 10203 14662
rect 10259 14610 10311 14662
rect 10367 14610 10419 14662
rect 10475 14610 10527 14662
rect 10583 14610 10635 14662
rect 10691 14610 10743 14662
rect 10799 14610 10851 14662
rect 10907 14610 10959 14662
rect 11015 14610 11067 14662
rect 11480 14718 11487 14770
rect 11487 14718 11532 14770
rect 11588 14718 11640 14770
rect 11696 14718 11748 14770
rect 11804 14718 11856 14770
rect 11912 14718 11964 14770
rect 11480 14610 11487 14662
rect 11487 14610 11532 14662
rect 11588 14610 11640 14662
rect 11696 14610 11748 14662
rect 11804 14610 11856 14662
rect 11912 14610 11964 14662
rect 467 10260 727 13120
rect 467 7060 727 9920
rect 467 3860 727 6720
rect 467 675 727 3535
rect 11682 10265 11942 13437
rect 11682 7055 11942 9915
rect 11682 3855 11942 6715
rect 11682 655 11942 3515
<< metal2 >>
rect -756 14778 -439 14820
rect -756 14759 -684 14778
rect -628 14759 -542 14778
rect -486 14759 -439 14778
rect -756 14707 -719 14759
rect -628 14722 -611 14759
rect -667 14707 -611 14722
rect -559 14722 -542 14759
rect -559 14707 -503 14722
rect -451 14707 -439 14759
rect -756 14651 -439 14707
rect -756 14599 -719 14651
rect -667 14636 -611 14651
rect -628 14599 -611 14636
rect -559 14636 -503 14651
rect -559 14599 -542 14636
rect -451 14599 -439 14651
rect -756 14580 -684 14599
rect -628 14580 -542 14599
rect -486 14580 -439 14599
rect -756 14563 -439 14580
rect 404 14778 912 14820
rect 404 14722 488 14778
rect 544 14770 630 14778
rect 686 14770 772 14778
rect 576 14722 630 14770
rect 686 14722 740 14770
rect 828 14722 912 14778
rect 404 14718 524 14722
rect 576 14718 632 14722
rect 684 14718 740 14722
rect 792 14718 912 14722
rect 404 14662 912 14718
rect 404 14636 524 14662
rect 576 14636 632 14662
rect 684 14636 740 14662
rect 792 14636 912 14662
rect 404 14580 488 14636
rect 576 14610 630 14636
rect 686 14610 740 14636
rect 544 14580 630 14610
rect 686 14580 772 14610
rect 828 14580 912 14636
rect 404 14563 912 14580
rect 1297 14778 2237 14820
rect 1297 14770 1313 14778
rect 1369 14770 1455 14778
rect 1511 14770 1597 14778
rect 1653 14770 1739 14778
rect 1795 14770 1881 14778
rect 1937 14770 2023 14778
rect 2079 14770 2165 14778
rect 2221 14770 2237 14778
rect 1297 14718 1309 14770
rect 1369 14722 1417 14770
rect 1511 14722 1525 14770
rect 1361 14718 1417 14722
rect 1469 14718 1525 14722
rect 1577 14722 1597 14770
rect 1685 14722 1739 14770
rect 1795 14722 1849 14770
rect 1937 14722 1957 14770
rect 1577 14718 1633 14722
rect 1685 14718 1741 14722
rect 1793 14718 1849 14722
rect 1901 14718 1957 14722
rect 2009 14722 2023 14770
rect 2117 14722 2165 14770
rect 2009 14718 2065 14722
rect 2117 14718 2173 14722
rect 2225 14718 2237 14770
rect 1297 14662 2237 14718
rect 1297 14610 1309 14662
rect 1361 14636 1417 14662
rect 1469 14636 1525 14662
rect 1369 14610 1417 14636
rect 1511 14610 1525 14636
rect 1577 14636 1633 14662
rect 1685 14636 1741 14662
rect 1793 14636 1849 14662
rect 1901 14636 1957 14662
rect 1577 14610 1597 14636
rect 1685 14610 1739 14636
rect 1795 14610 1849 14636
rect 1937 14610 1957 14636
rect 2009 14636 2065 14662
rect 2117 14636 2173 14662
rect 2009 14610 2023 14636
rect 2117 14610 2165 14636
rect 2225 14610 2237 14662
rect 1297 14580 1313 14610
rect 1369 14580 1455 14610
rect 1511 14580 1597 14610
rect 1653 14580 1739 14610
rect 1795 14580 1881 14610
rect 1937 14580 2023 14610
rect 2079 14580 2165 14610
rect 2221 14580 2237 14610
rect 1297 14563 2237 14580
rect 3064 14778 4004 14820
rect 3064 14770 3080 14778
rect 3136 14770 3222 14778
rect 3278 14770 3364 14778
rect 3420 14770 3506 14778
rect 3562 14770 3648 14778
rect 3704 14770 3790 14778
rect 3846 14770 3932 14778
rect 3988 14770 4004 14778
rect 3064 14718 3076 14770
rect 3136 14722 3184 14770
rect 3278 14722 3292 14770
rect 3128 14718 3184 14722
rect 3236 14718 3292 14722
rect 3344 14722 3364 14770
rect 3452 14722 3506 14770
rect 3562 14722 3616 14770
rect 3704 14722 3724 14770
rect 3344 14718 3400 14722
rect 3452 14718 3508 14722
rect 3560 14718 3616 14722
rect 3668 14718 3724 14722
rect 3776 14722 3790 14770
rect 3884 14722 3932 14770
rect 3776 14718 3832 14722
rect 3884 14718 3940 14722
rect 3992 14718 4004 14770
rect 3064 14662 4004 14718
rect 3064 14610 3076 14662
rect 3128 14636 3184 14662
rect 3236 14636 3292 14662
rect 3136 14610 3184 14636
rect 3278 14610 3292 14636
rect 3344 14636 3400 14662
rect 3452 14636 3508 14662
rect 3560 14636 3616 14662
rect 3668 14636 3724 14662
rect 3344 14610 3364 14636
rect 3452 14610 3506 14636
rect 3562 14610 3616 14636
rect 3704 14610 3724 14636
rect 3776 14636 3832 14662
rect 3884 14636 3940 14662
rect 3776 14610 3790 14636
rect 3884 14610 3932 14636
rect 3992 14610 4004 14662
rect 3064 14580 3080 14610
rect 3136 14580 3222 14610
rect 3278 14580 3364 14610
rect 3420 14580 3506 14610
rect 3562 14580 3648 14610
rect 3704 14580 3790 14610
rect 3846 14580 3932 14610
rect 3988 14580 4004 14610
rect 3064 14563 4004 14580
rect 4831 14778 5771 14820
rect 4831 14770 4847 14778
rect 4903 14770 4989 14778
rect 5045 14770 5131 14778
rect 5187 14770 5273 14778
rect 5329 14770 5415 14778
rect 5471 14770 5557 14778
rect 5613 14770 5699 14778
rect 5755 14770 5771 14778
rect 4831 14718 4843 14770
rect 4903 14722 4951 14770
rect 5045 14722 5059 14770
rect 4895 14718 4951 14722
rect 5003 14718 5059 14722
rect 5111 14722 5131 14770
rect 5219 14722 5273 14770
rect 5329 14722 5383 14770
rect 5471 14722 5491 14770
rect 5111 14718 5167 14722
rect 5219 14718 5275 14722
rect 5327 14718 5383 14722
rect 5435 14718 5491 14722
rect 5543 14722 5557 14770
rect 5651 14722 5699 14770
rect 5543 14718 5599 14722
rect 5651 14718 5707 14722
rect 5759 14718 5771 14770
rect 4831 14662 5771 14718
rect 4831 14610 4843 14662
rect 4895 14636 4951 14662
rect 5003 14636 5059 14662
rect 4903 14610 4951 14636
rect 5045 14610 5059 14636
rect 5111 14636 5167 14662
rect 5219 14636 5275 14662
rect 5327 14636 5383 14662
rect 5435 14636 5491 14662
rect 5111 14610 5131 14636
rect 5219 14610 5273 14636
rect 5329 14610 5383 14636
rect 5471 14610 5491 14636
rect 5543 14636 5599 14662
rect 5651 14636 5707 14662
rect 5543 14610 5557 14636
rect 5651 14610 5699 14636
rect 5759 14610 5771 14662
rect 4831 14580 4847 14610
rect 4903 14580 4989 14610
rect 5045 14580 5131 14610
rect 5187 14580 5273 14610
rect 5329 14580 5415 14610
rect 5471 14580 5557 14610
rect 5613 14580 5699 14610
rect 5755 14580 5771 14610
rect 4831 14563 5771 14580
rect 6605 14778 7545 14820
rect 6605 14770 6621 14778
rect 6677 14770 6763 14778
rect 6819 14770 6905 14778
rect 6961 14770 7047 14778
rect 7103 14770 7189 14778
rect 7245 14770 7331 14778
rect 7387 14770 7473 14778
rect 7529 14770 7545 14778
rect 6605 14718 6617 14770
rect 6677 14722 6725 14770
rect 6819 14722 6833 14770
rect 6669 14718 6725 14722
rect 6777 14718 6833 14722
rect 6885 14722 6905 14770
rect 6993 14722 7047 14770
rect 7103 14722 7157 14770
rect 7245 14722 7265 14770
rect 6885 14718 6941 14722
rect 6993 14718 7049 14722
rect 7101 14718 7157 14722
rect 7209 14718 7265 14722
rect 7317 14722 7331 14770
rect 7425 14722 7473 14770
rect 7317 14718 7373 14722
rect 7425 14718 7481 14722
rect 7533 14718 7545 14770
rect 6605 14662 7545 14718
rect 6605 14610 6617 14662
rect 6669 14636 6725 14662
rect 6777 14636 6833 14662
rect 6677 14610 6725 14636
rect 6819 14610 6833 14636
rect 6885 14636 6941 14662
rect 6993 14636 7049 14662
rect 7101 14636 7157 14662
rect 7209 14636 7265 14662
rect 6885 14610 6905 14636
rect 6993 14610 7047 14636
rect 7103 14610 7157 14636
rect 7245 14610 7265 14636
rect 7317 14636 7373 14662
rect 7425 14636 7481 14662
rect 7317 14610 7331 14636
rect 7425 14610 7473 14636
rect 7533 14610 7545 14662
rect 6605 14580 6621 14610
rect 6677 14580 6763 14610
rect 6819 14580 6905 14610
rect 6961 14580 7047 14610
rect 7103 14580 7189 14610
rect 7245 14580 7331 14610
rect 7387 14580 7473 14610
rect 7529 14580 7545 14610
rect 6605 14563 7545 14580
rect 8369 14778 9309 14820
rect 8369 14770 8385 14778
rect 8441 14770 8527 14778
rect 8583 14770 8669 14778
rect 8725 14770 8811 14778
rect 8867 14770 8953 14778
rect 9009 14770 9095 14778
rect 9151 14770 9237 14778
rect 9293 14770 9309 14778
rect 8369 14718 8381 14770
rect 8441 14722 8489 14770
rect 8583 14722 8597 14770
rect 8433 14718 8489 14722
rect 8541 14718 8597 14722
rect 8649 14722 8669 14770
rect 8757 14722 8811 14770
rect 8867 14722 8921 14770
rect 9009 14722 9029 14770
rect 8649 14718 8705 14722
rect 8757 14718 8813 14722
rect 8865 14718 8921 14722
rect 8973 14718 9029 14722
rect 9081 14722 9095 14770
rect 9189 14722 9237 14770
rect 9081 14718 9137 14722
rect 9189 14718 9245 14722
rect 9297 14718 9309 14770
rect 8369 14662 9309 14718
rect 8369 14610 8381 14662
rect 8433 14636 8489 14662
rect 8541 14636 8597 14662
rect 8441 14610 8489 14636
rect 8583 14610 8597 14636
rect 8649 14636 8705 14662
rect 8757 14636 8813 14662
rect 8865 14636 8921 14662
rect 8973 14636 9029 14662
rect 8649 14610 8669 14636
rect 8757 14610 8811 14636
rect 8867 14610 8921 14636
rect 9009 14610 9029 14636
rect 9081 14636 9137 14662
rect 9189 14636 9245 14662
rect 9081 14610 9095 14636
rect 9189 14610 9237 14636
rect 9297 14610 9309 14662
rect 8369 14580 8385 14610
rect 8441 14580 8527 14610
rect 8583 14580 8669 14610
rect 8725 14580 8811 14610
rect 8867 14580 8953 14610
rect 9009 14580 9095 14610
rect 9151 14580 9237 14610
rect 9293 14580 9309 14610
rect 8369 14563 9309 14580
rect 10139 14789 11079 14820
rect 10139 14770 10155 14789
rect 10211 14770 10297 14789
rect 10353 14770 10439 14789
rect 10495 14770 10581 14789
rect 10637 14770 10723 14789
rect 10779 14770 10865 14789
rect 10921 14770 11007 14789
rect 11063 14770 11079 14789
rect 10139 14718 10151 14770
rect 10211 14733 10259 14770
rect 10353 14733 10367 14770
rect 10203 14718 10259 14733
rect 10311 14718 10367 14733
rect 10419 14733 10439 14770
rect 10527 14733 10581 14770
rect 10637 14733 10691 14770
rect 10779 14733 10799 14770
rect 10419 14718 10475 14733
rect 10527 14718 10583 14733
rect 10635 14718 10691 14733
rect 10743 14718 10799 14733
rect 10851 14733 10865 14770
rect 10959 14733 11007 14770
rect 10851 14718 10907 14733
rect 10959 14718 11015 14733
rect 11067 14718 11079 14770
rect 10139 14662 11079 14718
rect 10139 14610 10151 14662
rect 10203 14647 10259 14662
rect 10311 14647 10367 14662
rect 10211 14610 10259 14647
rect 10353 14610 10367 14647
rect 10419 14647 10475 14662
rect 10527 14647 10583 14662
rect 10635 14647 10691 14662
rect 10743 14647 10799 14662
rect 10419 14610 10439 14647
rect 10527 14610 10581 14647
rect 10637 14610 10691 14647
rect 10779 14610 10799 14647
rect 10851 14647 10907 14662
rect 10959 14647 11015 14662
rect 10851 14610 10865 14647
rect 10959 14610 11007 14647
rect 11067 14610 11079 14662
rect 10139 14591 10155 14610
rect 10211 14591 10297 14610
rect 10353 14591 10439 14610
rect 10495 14591 10581 14610
rect 10637 14591 10723 14610
rect 10779 14591 10865 14610
rect 10921 14591 11007 14610
rect 11063 14591 11079 14610
rect 10139 14563 11079 14591
rect 11468 14778 11976 14820
rect 11468 14770 11481 14778
rect 11537 14770 11623 14778
rect 11679 14770 11765 14778
rect 11821 14770 11907 14778
rect 11963 14770 11976 14778
rect 11468 14718 11480 14770
rect 11537 14722 11588 14770
rect 11679 14722 11696 14770
rect 11532 14718 11588 14722
rect 11640 14718 11696 14722
rect 11748 14722 11765 14770
rect 11856 14722 11907 14770
rect 11748 14718 11804 14722
rect 11856 14718 11912 14722
rect 11964 14718 11976 14770
rect 11468 14662 11976 14718
rect 11468 14610 11480 14662
rect 11532 14636 11588 14662
rect 11640 14636 11696 14662
rect 11537 14610 11588 14636
rect 11679 14610 11696 14636
rect 11748 14636 11804 14662
rect 11856 14636 11912 14662
rect 11748 14610 11765 14636
rect 11856 14610 11907 14636
rect 11964 14610 11976 14662
rect 11468 14580 11481 14610
rect 11537 14580 11623 14610
rect 11679 14580 11765 14610
rect 11821 14580 11907 14610
rect 11963 14580 11976 14610
rect 11468 14563 11976 14580
rect 11617 13437 12003 13496
rect 393 13138 779 13173
rect 393 13120 498 13138
rect 554 13120 640 13138
rect 696 13120 779 13138
rect 393 10260 467 13120
rect 727 10260 779 13120
rect 393 10242 498 10260
rect 554 10242 640 10260
rect 696 10242 779 10260
rect 393 10188 779 10242
rect 11617 13133 11682 13437
rect 11942 13133 12003 13437
rect 11617 13077 11653 13133
rect 11993 13077 12003 13133
rect 11617 12991 11682 13077
rect 11942 12991 12003 13077
rect 11617 12935 11653 12991
rect 11993 12935 12003 12991
rect 11617 12849 11682 12935
rect 11942 12849 12003 12935
rect 11617 12793 11653 12849
rect 11993 12793 12003 12849
rect 11617 12707 11682 12793
rect 11942 12707 12003 12793
rect 11617 12651 11653 12707
rect 11993 12651 12003 12707
rect 11617 12565 11682 12651
rect 11942 12565 12003 12651
rect 11617 12509 11653 12565
rect 11993 12509 12003 12565
rect 11617 12423 11682 12509
rect 11942 12423 12003 12509
rect 11617 12367 11653 12423
rect 11993 12367 12003 12423
rect 11617 12281 11682 12367
rect 11942 12281 12003 12367
rect 11617 12225 11653 12281
rect 11993 12225 12003 12281
rect 11617 12139 11682 12225
rect 11942 12139 12003 12225
rect 11617 12083 11653 12139
rect 11993 12083 12003 12139
rect 11617 11997 11682 12083
rect 11942 11997 12003 12083
rect 11617 11941 11653 11997
rect 11993 11941 12003 11997
rect 11617 11855 11682 11941
rect 11942 11855 12003 11941
rect 11617 11799 11653 11855
rect 11993 11799 12003 11855
rect 11617 11713 11682 11799
rect 11942 11713 12003 11799
rect 11617 11657 11653 11713
rect 11993 11657 12003 11713
rect 11617 11571 11682 11657
rect 11942 11571 12003 11657
rect 11617 11515 11653 11571
rect 11993 11515 12003 11571
rect 11617 11429 11682 11515
rect 11942 11429 12003 11515
rect 11617 11373 11653 11429
rect 11993 11373 12003 11429
rect 11617 11287 11682 11373
rect 11942 11287 12003 11373
rect 11617 11231 11653 11287
rect 11993 11231 12003 11287
rect 11617 11145 11682 11231
rect 11942 11145 12003 11231
rect 11617 11089 11653 11145
rect 11993 11089 12003 11145
rect 11617 11003 11682 11089
rect 11942 11003 12003 11089
rect 11617 10947 11653 11003
rect 11993 10947 12003 11003
rect 11617 10861 11682 10947
rect 11942 10861 12003 10947
rect 11617 10805 11653 10861
rect 11993 10805 12003 10861
rect 11617 10719 11682 10805
rect 11942 10719 12003 10805
rect 11617 10663 11653 10719
rect 11993 10663 12003 10719
rect 11617 10577 11682 10663
rect 11942 10577 12003 10663
rect 11617 10521 11653 10577
rect 11993 10521 12003 10577
rect 11617 10435 11682 10521
rect 11942 10435 12003 10521
rect 11617 10379 11653 10435
rect 11993 10379 12003 10435
rect 11617 10293 11682 10379
rect 11942 10293 12003 10379
rect 11617 10237 11653 10293
rect 11709 10237 11795 10265
rect 11851 10237 11937 10265
rect 11993 10237 12003 10293
rect 11617 10188 12003 10237
rect 393 9938 779 9973
rect 393 9920 498 9938
rect 554 9920 640 9938
rect 696 9920 779 9938
rect 393 7060 467 9920
rect 727 7060 779 9920
rect 393 7042 498 7060
rect 554 7042 640 7060
rect 696 7042 779 7060
rect 393 6988 779 7042
rect 11617 9933 12003 9988
rect 11617 9877 11653 9933
rect 11709 9915 11795 9933
rect 11851 9915 11937 9933
rect 11993 9877 12003 9933
rect 11617 9791 11682 9877
rect 11942 9791 12003 9877
rect 11617 9735 11653 9791
rect 11993 9735 12003 9791
rect 11617 9649 11682 9735
rect 11942 9649 12003 9735
rect 11617 9593 11653 9649
rect 11993 9593 12003 9649
rect 11617 9507 11682 9593
rect 11942 9507 12003 9593
rect 11617 9451 11653 9507
rect 11993 9451 12003 9507
rect 11617 9365 11682 9451
rect 11942 9365 12003 9451
rect 11617 9309 11653 9365
rect 11993 9309 12003 9365
rect 11617 9223 11682 9309
rect 11942 9223 12003 9309
rect 11617 9167 11653 9223
rect 11993 9167 12003 9223
rect 11617 9081 11682 9167
rect 11942 9081 12003 9167
rect 11617 9025 11653 9081
rect 11993 9025 12003 9081
rect 11617 8939 11682 9025
rect 11942 8939 12003 9025
rect 11617 8883 11653 8939
rect 11993 8883 12003 8939
rect 11617 8797 11682 8883
rect 11942 8797 12003 8883
rect 11617 8741 11653 8797
rect 11993 8741 12003 8797
rect 11617 8655 11682 8741
rect 11942 8655 12003 8741
rect 11617 8599 11653 8655
rect 11993 8599 12003 8655
rect 11617 8513 11682 8599
rect 11942 8513 12003 8599
rect 11617 8457 11653 8513
rect 11993 8457 12003 8513
rect 11617 8371 11682 8457
rect 11942 8371 12003 8457
rect 11617 8315 11653 8371
rect 11993 8315 12003 8371
rect 11617 8229 11682 8315
rect 11942 8229 12003 8315
rect 11617 8173 11653 8229
rect 11993 8173 12003 8229
rect 11617 8087 11682 8173
rect 11942 8087 12003 8173
rect 11617 8031 11653 8087
rect 11993 8031 12003 8087
rect 11617 7945 11682 8031
rect 11942 7945 12003 8031
rect 11617 7889 11653 7945
rect 11993 7889 12003 7945
rect 11617 7803 11682 7889
rect 11942 7803 12003 7889
rect 11617 7747 11653 7803
rect 11993 7747 12003 7803
rect 11617 7661 11682 7747
rect 11942 7661 12003 7747
rect 11617 7605 11653 7661
rect 11993 7605 12003 7661
rect 11617 7519 11682 7605
rect 11942 7519 12003 7605
rect 11617 7463 11653 7519
rect 11993 7463 12003 7519
rect 11617 7377 11682 7463
rect 11942 7377 12003 7463
rect 11617 7321 11653 7377
rect 11993 7321 12003 7377
rect 11617 7235 11682 7321
rect 11942 7235 12003 7321
rect 11617 7179 11653 7235
rect 11993 7179 12003 7235
rect 11617 7093 11682 7179
rect 11942 7093 12003 7179
rect 11617 7037 11653 7093
rect 11709 7037 11795 7055
rect 11851 7037 11937 7055
rect 11993 7037 12003 7093
rect 11617 6988 12003 7037
rect 393 6738 779 6773
rect 393 6720 498 6738
rect 554 6720 640 6738
rect 696 6720 779 6738
rect 393 3860 467 6720
rect 727 3860 779 6720
rect 393 3842 498 3860
rect 554 3842 640 3860
rect 696 3842 779 3860
rect 393 3788 779 3842
rect 11617 6733 12003 6788
rect 11617 6677 11653 6733
rect 11709 6715 11795 6733
rect 11851 6715 11937 6733
rect 11993 6677 12003 6733
rect 11617 6591 11682 6677
rect 11942 6591 12003 6677
rect 11617 6535 11653 6591
rect 11993 6535 12003 6591
rect 11617 6449 11682 6535
rect 11942 6449 12003 6535
rect 11617 6393 11653 6449
rect 11993 6393 12003 6449
rect 11617 6307 11682 6393
rect 11942 6307 12003 6393
rect 11617 6251 11653 6307
rect 11993 6251 12003 6307
rect 11617 6165 11682 6251
rect 11942 6165 12003 6251
rect 11617 6109 11653 6165
rect 11993 6109 12003 6165
rect 11617 6023 11682 6109
rect 11942 6023 12003 6109
rect 11617 5967 11653 6023
rect 11993 5967 12003 6023
rect 11617 5881 11682 5967
rect 11942 5881 12003 5967
rect 11617 5825 11653 5881
rect 11993 5825 12003 5881
rect 11617 5739 11682 5825
rect 11942 5739 12003 5825
rect 11617 5683 11653 5739
rect 11993 5683 12003 5739
rect 11617 5597 11682 5683
rect 11942 5597 12003 5683
rect 11617 5541 11653 5597
rect 11993 5541 12003 5597
rect 11617 5455 11682 5541
rect 11942 5455 12003 5541
rect 11617 5399 11653 5455
rect 11993 5399 12003 5455
rect 11617 5313 11682 5399
rect 11942 5313 12003 5399
rect 11617 5257 11653 5313
rect 11993 5257 12003 5313
rect 11617 5171 11682 5257
rect 11942 5171 12003 5257
rect 11617 5115 11653 5171
rect 11993 5115 12003 5171
rect 11617 5029 11682 5115
rect 11942 5029 12003 5115
rect 11617 4973 11653 5029
rect 11993 4973 12003 5029
rect 11617 4887 11682 4973
rect 11942 4887 12003 4973
rect 11617 4831 11653 4887
rect 11993 4831 12003 4887
rect 11617 4745 11682 4831
rect 11942 4745 12003 4831
rect 11617 4689 11653 4745
rect 11993 4689 12003 4745
rect 11617 4603 11682 4689
rect 11942 4603 12003 4689
rect 11617 4547 11653 4603
rect 11993 4547 12003 4603
rect 11617 4461 11682 4547
rect 11942 4461 12003 4547
rect 11617 4405 11653 4461
rect 11993 4405 12003 4461
rect 11617 4319 11682 4405
rect 11942 4319 12003 4405
rect 11617 4263 11653 4319
rect 11993 4263 12003 4319
rect 11617 4177 11682 4263
rect 11942 4177 12003 4263
rect 11617 4121 11653 4177
rect 11993 4121 12003 4177
rect 11617 4035 11682 4121
rect 11942 4035 12003 4121
rect 11617 3979 11653 4035
rect 11993 3979 12003 4035
rect 11617 3893 11682 3979
rect 11942 3893 12003 3979
rect 11617 3837 11653 3893
rect 11709 3837 11795 3855
rect 11851 3837 11937 3855
rect 11993 3837 12003 3893
rect 11617 3788 12003 3837
rect 393 3553 779 3588
rect 393 3535 498 3553
rect 554 3535 640 3553
rect 696 3535 779 3553
rect 393 675 467 3535
rect 727 675 779 3535
rect 393 657 498 675
rect 554 657 640 675
rect 696 657 779 675
rect 393 496 779 657
rect 11617 3533 12003 3588
rect 11617 3477 11653 3533
rect 11709 3515 11795 3533
rect 11851 3515 11937 3533
rect 11993 3477 12003 3533
rect 11617 3391 11682 3477
rect 11942 3391 12003 3477
rect 11617 3335 11653 3391
rect 11993 3335 12003 3391
rect 11617 3249 11682 3335
rect 11942 3249 12003 3335
rect 11617 3193 11653 3249
rect 11993 3193 12003 3249
rect 11617 3107 11682 3193
rect 11942 3107 12003 3193
rect 11617 3051 11653 3107
rect 11993 3051 12003 3107
rect 11617 2965 11682 3051
rect 11942 2965 12003 3051
rect 11617 2909 11653 2965
rect 11993 2909 12003 2965
rect 11617 2823 11682 2909
rect 11942 2823 12003 2909
rect 11617 2767 11653 2823
rect 11993 2767 12003 2823
rect 11617 2681 11682 2767
rect 11942 2681 12003 2767
rect 11617 2625 11653 2681
rect 11993 2625 12003 2681
rect 11617 2539 11682 2625
rect 11942 2539 12003 2625
rect 11617 2483 11653 2539
rect 11993 2483 12003 2539
rect 11617 2397 11682 2483
rect 11942 2397 12003 2483
rect 11617 2341 11653 2397
rect 11993 2341 12003 2397
rect 11617 2255 11682 2341
rect 11942 2255 12003 2341
rect 11617 2199 11653 2255
rect 11993 2199 12003 2255
rect 11617 2113 11682 2199
rect 11942 2113 12003 2199
rect 11617 2057 11653 2113
rect 11993 2057 12003 2113
rect 11617 1971 11682 2057
rect 11942 1971 12003 2057
rect 11617 1915 11653 1971
rect 11993 1915 12003 1971
rect 11617 1829 11682 1915
rect 11942 1829 12003 1915
rect 11617 1773 11653 1829
rect 11993 1773 12003 1829
rect 11617 1687 11682 1773
rect 11942 1687 12003 1773
rect 11617 1631 11653 1687
rect 11993 1631 12003 1687
rect 11617 1545 11682 1631
rect 11942 1545 12003 1631
rect 11617 1489 11653 1545
rect 11993 1489 12003 1545
rect 11617 1403 11682 1489
rect 11942 1403 12003 1489
rect 11617 1347 11653 1403
rect 11993 1347 12003 1403
rect 11617 1261 11682 1347
rect 11942 1261 12003 1347
rect 11617 1205 11653 1261
rect 11993 1205 12003 1261
rect 11617 1119 11682 1205
rect 11942 1119 12003 1205
rect 11617 1063 11653 1119
rect 11993 1063 12003 1119
rect 11617 977 11682 1063
rect 11942 977 12003 1063
rect 11617 921 11653 977
rect 11993 921 12003 977
rect 11617 835 11682 921
rect 11942 835 12003 921
rect 11617 779 11653 835
rect 11993 779 12003 835
rect 11617 693 11682 779
rect 11942 693 12003 779
rect 11617 637 11653 693
rect 11709 637 11795 655
rect 11851 637 11937 655
rect 11993 637 12003 693
rect 11617 496 12003 637
<< via2 >>
rect -684 14759 -628 14778
rect -542 14759 -486 14778
rect -684 14722 -667 14759
rect -667 14722 -628 14759
rect -542 14722 -503 14759
rect -503 14722 -486 14759
rect -684 14599 -667 14636
rect -667 14599 -628 14636
rect -542 14599 -503 14636
rect -503 14599 -486 14636
rect -684 14580 -628 14599
rect -542 14580 -486 14599
rect 488 14770 544 14778
rect 630 14770 686 14778
rect 772 14770 828 14778
rect 488 14722 524 14770
rect 524 14722 544 14770
rect 630 14722 632 14770
rect 632 14722 684 14770
rect 684 14722 686 14770
rect 772 14722 792 14770
rect 792 14722 828 14770
rect 488 14610 524 14636
rect 524 14610 544 14636
rect 630 14610 632 14636
rect 632 14610 684 14636
rect 684 14610 686 14636
rect 772 14610 792 14636
rect 792 14610 828 14636
rect 488 14580 544 14610
rect 630 14580 686 14610
rect 772 14580 828 14610
rect 1313 14770 1369 14778
rect 1455 14770 1511 14778
rect 1597 14770 1653 14778
rect 1739 14770 1795 14778
rect 1881 14770 1937 14778
rect 2023 14770 2079 14778
rect 2165 14770 2221 14778
rect 1313 14722 1361 14770
rect 1361 14722 1369 14770
rect 1455 14722 1469 14770
rect 1469 14722 1511 14770
rect 1597 14722 1633 14770
rect 1633 14722 1653 14770
rect 1739 14722 1741 14770
rect 1741 14722 1793 14770
rect 1793 14722 1795 14770
rect 1881 14722 1901 14770
rect 1901 14722 1937 14770
rect 2023 14722 2065 14770
rect 2065 14722 2079 14770
rect 2165 14722 2173 14770
rect 2173 14722 2221 14770
rect 1313 14610 1361 14636
rect 1361 14610 1369 14636
rect 1455 14610 1469 14636
rect 1469 14610 1511 14636
rect 1597 14610 1633 14636
rect 1633 14610 1653 14636
rect 1739 14610 1741 14636
rect 1741 14610 1793 14636
rect 1793 14610 1795 14636
rect 1881 14610 1901 14636
rect 1901 14610 1937 14636
rect 2023 14610 2065 14636
rect 2065 14610 2079 14636
rect 2165 14610 2173 14636
rect 2173 14610 2221 14636
rect 1313 14580 1369 14610
rect 1455 14580 1511 14610
rect 1597 14580 1653 14610
rect 1739 14580 1795 14610
rect 1881 14580 1937 14610
rect 2023 14580 2079 14610
rect 2165 14580 2221 14610
rect 3080 14770 3136 14778
rect 3222 14770 3278 14778
rect 3364 14770 3420 14778
rect 3506 14770 3562 14778
rect 3648 14770 3704 14778
rect 3790 14770 3846 14778
rect 3932 14770 3988 14778
rect 3080 14722 3128 14770
rect 3128 14722 3136 14770
rect 3222 14722 3236 14770
rect 3236 14722 3278 14770
rect 3364 14722 3400 14770
rect 3400 14722 3420 14770
rect 3506 14722 3508 14770
rect 3508 14722 3560 14770
rect 3560 14722 3562 14770
rect 3648 14722 3668 14770
rect 3668 14722 3704 14770
rect 3790 14722 3832 14770
rect 3832 14722 3846 14770
rect 3932 14722 3940 14770
rect 3940 14722 3988 14770
rect 3080 14610 3128 14636
rect 3128 14610 3136 14636
rect 3222 14610 3236 14636
rect 3236 14610 3278 14636
rect 3364 14610 3400 14636
rect 3400 14610 3420 14636
rect 3506 14610 3508 14636
rect 3508 14610 3560 14636
rect 3560 14610 3562 14636
rect 3648 14610 3668 14636
rect 3668 14610 3704 14636
rect 3790 14610 3832 14636
rect 3832 14610 3846 14636
rect 3932 14610 3940 14636
rect 3940 14610 3988 14636
rect 3080 14580 3136 14610
rect 3222 14580 3278 14610
rect 3364 14580 3420 14610
rect 3506 14580 3562 14610
rect 3648 14580 3704 14610
rect 3790 14580 3846 14610
rect 3932 14580 3988 14610
rect 4847 14770 4903 14778
rect 4989 14770 5045 14778
rect 5131 14770 5187 14778
rect 5273 14770 5329 14778
rect 5415 14770 5471 14778
rect 5557 14770 5613 14778
rect 5699 14770 5755 14778
rect 4847 14722 4895 14770
rect 4895 14722 4903 14770
rect 4989 14722 5003 14770
rect 5003 14722 5045 14770
rect 5131 14722 5167 14770
rect 5167 14722 5187 14770
rect 5273 14722 5275 14770
rect 5275 14722 5327 14770
rect 5327 14722 5329 14770
rect 5415 14722 5435 14770
rect 5435 14722 5471 14770
rect 5557 14722 5599 14770
rect 5599 14722 5613 14770
rect 5699 14722 5707 14770
rect 5707 14722 5755 14770
rect 4847 14610 4895 14636
rect 4895 14610 4903 14636
rect 4989 14610 5003 14636
rect 5003 14610 5045 14636
rect 5131 14610 5167 14636
rect 5167 14610 5187 14636
rect 5273 14610 5275 14636
rect 5275 14610 5327 14636
rect 5327 14610 5329 14636
rect 5415 14610 5435 14636
rect 5435 14610 5471 14636
rect 5557 14610 5599 14636
rect 5599 14610 5613 14636
rect 5699 14610 5707 14636
rect 5707 14610 5755 14636
rect 4847 14580 4903 14610
rect 4989 14580 5045 14610
rect 5131 14580 5187 14610
rect 5273 14580 5329 14610
rect 5415 14580 5471 14610
rect 5557 14580 5613 14610
rect 5699 14580 5755 14610
rect 6621 14770 6677 14778
rect 6763 14770 6819 14778
rect 6905 14770 6961 14778
rect 7047 14770 7103 14778
rect 7189 14770 7245 14778
rect 7331 14770 7387 14778
rect 7473 14770 7529 14778
rect 6621 14722 6669 14770
rect 6669 14722 6677 14770
rect 6763 14722 6777 14770
rect 6777 14722 6819 14770
rect 6905 14722 6941 14770
rect 6941 14722 6961 14770
rect 7047 14722 7049 14770
rect 7049 14722 7101 14770
rect 7101 14722 7103 14770
rect 7189 14722 7209 14770
rect 7209 14722 7245 14770
rect 7331 14722 7373 14770
rect 7373 14722 7387 14770
rect 7473 14722 7481 14770
rect 7481 14722 7529 14770
rect 6621 14610 6669 14636
rect 6669 14610 6677 14636
rect 6763 14610 6777 14636
rect 6777 14610 6819 14636
rect 6905 14610 6941 14636
rect 6941 14610 6961 14636
rect 7047 14610 7049 14636
rect 7049 14610 7101 14636
rect 7101 14610 7103 14636
rect 7189 14610 7209 14636
rect 7209 14610 7245 14636
rect 7331 14610 7373 14636
rect 7373 14610 7387 14636
rect 7473 14610 7481 14636
rect 7481 14610 7529 14636
rect 6621 14580 6677 14610
rect 6763 14580 6819 14610
rect 6905 14580 6961 14610
rect 7047 14580 7103 14610
rect 7189 14580 7245 14610
rect 7331 14580 7387 14610
rect 7473 14580 7529 14610
rect 8385 14770 8441 14778
rect 8527 14770 8583 14778
rect 8669 14770 8725 14778
rect 8811 14770 8867 14778
rect 8953 14770 9009 14778
rect 9095 14770 9151 14778
rect 9237 14770 9293 14778
rect 8385 14722 8433 14770
rect 8433 14722 8441 14770
rect 8527 14722 8541 14770
rect 8541 14722 8583 14770
rect 8669 14722 8705 14770
rect 8705 14722 8725 14770
rect 8811 14722 8813 14770
rect 8813 14722 8865 14770
rect 8865 14722 8867 14770
rect 8953 14722 8973 14770
rect 8973 14722 9009 14770
rect 9095 14722 9137 14770
rect 9137 14722 9151 14770
rect 9237 14722 9245 14770
rect 9245 14722 9293 14770
rect 8385 14610 8433 14636
rect 8433 14610 8441 14636
rect 8527 14610 8541 14636
rect 8541 14610 8583 14636
rect 8669 14610 8705 14636
rect 8705 14610 8725 14636
rect 8811 14610 8813 14636
rect 8813 14610 8865 14636
rect 8865 14610 8867 14636
rect 8953 14610 8973 14636
rect 8973 14610 9009 14636
rect 9095 14610 9137 14636
rect 9137 14610 9151 14636
rect 9237 14610 9245 14636
rect 9245 14610 9293 14636
rect 8385 14580 8441 14610
rect 8527 14580 8583 14610
rect 8669 14580 8725 14610
rect 8811 14580 8867 14610
rect 8953 14580 9009 14610
rect 9095 14580 9151 14610
rect 9237 14580 9293 14610
rect 10155 14770 10211 14789
rect 10297 14770 10353 14789
rect 10439 14770 10495 14789
rect 10581 14770 10637 14789
rect 10723 14770 10779 14789
rect 10865 14770 10921 14789
rect 11007 14770 11063 14789
rect 10155 14733 10203 14770
rect 10203 14733 10211 14770
rect 10297 14733 10311 14770
rect 10311 14733 10353 14770
rect 10439 14733 10475 14770
rect 10475 14733 10495 14770
rect 10581 14733 10583 14770
rect 10583 14733 10635 14770
rect 10635 14733 10637 14770
rect 10723 14733 10743 14770
rect 10743 14733 10779 14770
rect 10865 14733 10907 14770
rect 10907 14733 10921 14770
rect 11007 14733 11015 14770
rect 11015 14733 11063 14770
rect 10155 14610 10203 14647
rect 10203 14610 10211 14647
rect 10297 14610 10311 14647
rect 10311 14610 10353 14647
rect 10439 14610 10475 14647
rect 10475 14610 10495 14647
rect 10581 14610 10583 14647
rect 10583 14610 10635 14647
rect 10635 14610 10637 14647
rect 10723 14610 10743 14647
rect 10743 14610 10779 14647
rect 10865 14610 10907 14647
rect 10907 14610 10921 14647
rect 11007 14610 11015 14647
rect 11015 14610 11063 14647
rect 10155 14591 10211 14610
rect 10297 14591 10353 14610
rect 10439 14591 10495 14610
rect 10581 14591 10637 14610
rect 10723 14591 10779 14610
rect 10865 14591 10921 14610
rect 11007 14591 11063 14610
rect 11481 14770 11537 14778
rect 11623 14770 11679 14778
rect 11765 14770 11821 14778
rect 11907 14770 11963 14778
rect 11481 14722 11532 14770
rect 11532 14722 11537 14770
rect 11623 14722 11640 14770
rect 11640 14722 11679 14770
rect 11765 14722 11804 14770
rect 11804 14722 11821 14770
rect 11907 14722 11912 14770
rect 11912 14722 11963 14770
rect 11481 14610 11532 14636
rect 11532 14610 11537 14636
rect 11623 14610 11640 14636
rect 11640 14610 11679 14636
rect 11765 14610 11804 14636
rect 11804 14610 11821 14636
rect 11907 14610 11912 14636
rect 11912 14610 11963 14636
rect 11481 14580 11537 14610
rect 11623 14580 11679 14610
rect 11765 14580 11821 14610
rect 11907 14580 11963 14610
rect 498 13120 554 13138
rect 640 13120 696 13138
rect 498 13082 554 13120
rect 640 13082 696 13120
rect 498 12940 554 12996
rect 640 12940 696 12996
rect 498 12798 554 12854
rect 640 12798 696 12854
rect 498 12656 554 12712
rect 640 12656 696 12712
rect 498 12514 554 12570
rect 640 12514 696 12570
rect 498 12372 554 12428
rect 640 12372 696 12428
rect 498 12230 554 12286
rect 640 12230 696 12286
rect 498 12088 554 12144
rect 640 12088 696 12144
rect 498 11946 554 12002
rect 640 11946 696 12002
rect 498 11804 554 11860
rect 640 11804 696 11860
rect 498 11662 554 11718
rect 640 11662 696 11718
rect 498 11520 554 11576
rect 640 11520 696 11576
rect 498 11378 554 11434
rect 640 11378 696 11434
rect 498 11236 554 11292
rect 640 11236 696 11292
rect 498 11094 554 11150
rect 640 11094 696 11150
rect 498 10952 554 11008
rect 640 10952 696 11008
rect 498 10810 554 10866
rect 640 10810 696 10866
rect 498 10668 554 10724
rect 640 10668 696 10724
rect 498 10526 554 10582
rect 640 10526 696 10582
rect 498 10384 554 10440
rect 640 10384 696 10440
rect 498 10260 554 10298
rect 640 10260 696 10298
rect 498 10242 554 10260
rect 640 10242 696 10260
rect 11653 13077 11682 13133
rect 11682 13077 11709 13133
rect 11795 13077 11851 13133
rect 11937 13077 11942 13133
rect 11942 13077 11993 13133
rect 11653 12935 11682 12991
rect 11682 12935 11709 12991
rect 11795 12935 11851 12991
rect 11937 12935 11942 12991
rect 11942 12935 11993 12991
rect 11653 12793 11682 12849
rect 11682 12793 11709 12849
rect 11795 12793 11851 12849
rect 11937 12793 11942 12849
rect 11942 12793 11993 12849
rect 11653 12651 11682 12707
rect 11682 12651 11709 12707
rect 11795 12651 11851 12707
rect 11937 12651 11942 12707
rect 11942 12651 11993 12707
rect 11653 12509 11682 12565
rect 11682 12509 11709 12565
rect 11795 12509 11851 12565
rect 11937 12509 11942 12565
rect 11942 12509 11993 12565
rect 11653 12367 11682 12423
rect 11682 12367 11709 12423
rect 11795 12367 11851 12423
rect 11937 12367 11942 12423
rect 11942 12367 11993 12423
rect 11653 12225 11682 12281
rect 11682 12225 11709 12281
rect 11795 12225 11851 12281
rect 11937 12225 11942 12281
rect 11942 12225 11993 12281
rect 11653 12083 11682 12139
rect 11682 12083 11709 12139
rect 11795 12083 11851 12139
rect 11937 12083 11942 12139
rect 11942 12083 11993 12139
rect 11653 11941 11682 11997
rect 11682 11941 11709 11997
rect 11795 11941 11851 11997
rect 11937 11941 11942 11997
rect 11942 11941 11993 11997
rect 11653 11799 11682 11855
rect 11682 11799 11709 11855
rect 11795 11799 11851 11855
rect 11937 11799 11942 11855
rect 11942 11799 11993 11855
rect 11653 11657 11682 11713
rect 11682 11657 11709 11713
rect 11795 11657 11851 11713
rect 11937 11657 11942 11713
rect 11942 11657 11993 11713
rect 11653 11515 11682 11571
rect 11682 11515 11709 11571
rect 11795 11515 11851 11571
rect 11937 11515 11942 11571
rect 11942 11515 11993 11571
rect 11653 11373 11682 11429
rect 11682 11373 11709 11429
rect 11795 11373 11851 11429
rect 11937 11373 11942 11429
rect 11942 11373 11993 11429
rect 11653 11231 11682 11287
rect 11682 11231 11709 11287
rect 11795 11231 11851 11287
rect 11937 11231 11942 11287
rect 11942 11231 11993 11287
rect 11653 11089 11682 11145
rect 11682 11089 11709 11145
rect 11795 11089 11851 11145
rect 11937 11089 11942 11145
rect 11942 11089 11993 11145
rect 11653 10947 11682 11003
rect 11682 10947 11709 11003
rect 11795 10947 11851 11003
rect 11937 10947 11942 11003
rect 11942 10947 11993 11003
rect 11653 10805 11682 10861
rect 11682 10805 11709 10861
rect 11795 10805 11851 10861
rect 11937 10805 11942 10861
rect 11942 10805 11993 10861
rect 11653 10663 11682 10719
rect 11682 10663 11709 10719
rect 11795 10663 11851 10719
rect 11937 10663 11942 10719
rect 11942 10663 11993 10719
rect 11653 10521 11682 10577
rect 11682 10521 11709 10577
rect 11795 10521 11851 10577
rect 11937 10521 11942 10577
rect 11942 10521 11993 10577
rect 11653 10379 11682 10435
rect 11682 10379 11709 10435
rect 11795 10379 11851 10435
rect 11937 10379 11942 10435
rect 11942 10379 11993 10435
rect 11653 10265 11682 10293
rect 11682 10265 11709 10293
rect 11795 10265 11851 10293
rect 11937 10265 11942 10293
rect 11942 10265 11993 10293
rect 11653 10237 11709 10265
rect 11795 10237 11851 10265
rect 11937 10237 11993 10265
rect 498 9920 554 9938
rect 640 9920 696 9938
rect 498 9882 554 9920
rect 640 9882 696 9920
rect 498 9740 554 9796
rect 640 9740 696 9796
rect 498 9598 554 9654
rect 640 9598 696 9654
rect 498 9456 554 9512
rect 640 9456 696 9512
rect 498 9314 554 9370
rect 640 9314 696 9370
rect 498 9172 554 9228
rect 640 9172 696 9228
rect 498 9030 554 9086
rect 640 9030 696 9086
rect 498 8888 554 8944
rect 640 8888 696 8944
rect 498 8746 554 8802
rect 640 8746 696 8802
rect 498 8604 554 8660
rect 640 8604 696 8660
rect 498 8462 554 8518
rect 640 8462 696 8518
rect 498 8320 554 8376
rect 640 8320 696 8376
rect 498 8178 554 8234
rect 640 8178 696 8234
rect 498 8036 554 8092
rect 640 8036 696 8092
rect 498 7894 554 7950
rect 640 7894 696 7950
rect 498 7752 554 7808
rect 640 7752 696 7808
rect 498 7610 554 7666
rect 640 7610 696 7666
rect 498 7468 554 7524
rect 640 7468 696 7524
rect 498 7326 554 7382
rect 640 7326 696 7382
rect 498 7184 554 7240
rect 640 7184 696 7240
rect 498 7060 554 7098
rect 640 7060 696 7098
rect 498 7042 554 7060
rect 640 7042 696 7060
rect 11653 9915 11709 9933
rect 11795 9915 11851 9933
rect 11937 9915 11993 9933
rect 11653 9877 11682 9915
rect 11682 9877 11709 9915
rect 11795 9877 11851 9915
rect 11937 9877 11942 9915
rect 11942 9877 11993 9915
rect 11653 9735 11682 9791
rect 11682 9735 11709 9791
rect 11795 9735 11851 9791
rect 11937 9735 11942 9791
rect 11942 9735 11993 9791
rect 11653 9593 11682 9649
rect 11682 9593 11709 9649
rect 11795 9593 11851 9649
rect 11937 9593 11942 9649
rect 11942 9593 11993 9649
rect 11653 9451 11682 9507
rect 11682 9451 11709 9507
rect 11795 9451 11851 9507
rect 11937 9451 11942 9507
rect 11942 9451 11993 9507
rect 11653 9309 11682 9365
rect 11682 9309 11709 9365
rect 11795 9309 11851 9365
rect 11937 9309 11942 9365
rect 11942 9309 11993 9365
rect 11653 9167 11682 9223
rect 11682 9167 11709 9223
rect 11795 9167 11851 9223
rect 11937 9167 11942 9223
rect 11942 9167 11993 9223
rect 11653 9025 11682 9081
rect 11682 9025 11709 9081
rect 11795 9025 11851 9081
rect 11937 9025 11942 9081
rect 11942 9025 11993 9081
rect 11653 8883 11682 8939
rect 11682 8883 11709 8939
rect 11795 8883 11851 8939
rect 11937 8883 11942 8939
rect 11942 8883 11993 8939
rect 11653 8741 11682 8797
rect 11682 8741 11709 8797
rect 11795 8741 11851 8797
rect 11937 8741 11942 8797
rect 11942 8741 11993 8797
rect 11653 8599 11682 8655
rect 11682 8599 11709 8655
rect 11795 8599 11851 8655
rect 11937 8599 11942 8655
rect 11942 8599 11993 8655
rect 11653 8457 11682 8513
rect 11682 8457 11709 8513
rect 11795 8457 11851 8513
rect 11937 8457 11942 8513
rect 11942 8457 11993 8513
rect 11653 8315 11682 8371
rect 11682 8315 11709 8371
rect 11795 8315 11851 8371
rect 11937 8315 11942 8371
rect 11942 8315 11993 8371
rect 11653 8173 11682 8229
rect 11682 8173 11709 8229
rect 11795 8173 11851 8229
rect 11937 8173 11942 8229
rect 11942 8173 11993 8229
rect 11653 8031 11682 8087
rect 11682 8031 11709 8087
rect 11795 8031 11851 8087
rect 11937 8031 11942 8087
rect 11942 8031 11993 8087
rect 11653 7889 11682 7945
rect 11682 7889 11709 7945
rect 11795 7889 11851 7945
rect 11937 7889 11942 7945
rect 11942 7889 11993 7945
rect 11653 7747 11682 7803
rect 11682 7747 11709 7803
rect 11795 7747 11851 7803
rect 11937 7747 11942 7803
rect 11942 7747 11993 7803
rect 11653 7605 11682 7661
rect 11682 7605 11709 7661
rect 11795 7605 11851 7661
rect 11937 7605 11942 7661
rect 11942 7605 11993 7661
rect 11653 7463 11682 7519
rect 11682 7463 11709 7519
rect 11795 7463 11851 7519
rect 11937 7463 11942 7519
rect 11942 7463 11993 7519
rect 11653 7321 11682 7377
rect 11682 7321 11709 7377
rect 11795 7321 11851 7377
rect 11937 7321 11942 7377
rect 11942 7321 11993 7377
rect 11653 7179 11682 7235
rect 11682 7179 11709 7235
rect 11795 7179 11851 7235
rect 11937 7179 11942 7235
rect 11942 7179 11993 7235
rect 11653 7055 11682 7093
rect 11682 7055 11709 7093
rect 11795 7055 11851 7093
rect 11937 7055 11942 7093
rect 11942 7055 11993 7093
rect 11653 7037 11709 7055
rect 11795 7037 11851 7055
rect 11937 7037 11993 7055
rect 498 6720 554 6738
rect 640 6720 696 6738
rect 498 6682 554 6720
rect 640 6682 696 6720
rect 498 6540 554 6596
rect 640 6540 696 6596
rect 498 6398 554 6454
rect 640 6398 696 6454
rect 498 6256 554 6312
rect 640 6256 696 6312
rect 498 6114 554 6170
rect 640 6114 696 6170
rect 498 5972 554 6028
rect 640 5972 696 6028
rect 498 5830 554 5886
rect 640 5830 696 5886
rect 498 5688 554 5744
rect 640 5688 696 5744
rect 498 5546 554 5602
rect 640 5546 696 5602
rect 498 5404 554 5460
rect 640 5404 696 5460
rect 498 5262 554 5318
rect 640 5262 696 5318
rect 498 5120 554 5176
rect 640 5120 696 5176
rect 498 4978 554 5034
rect 640 4978 696 5034
rect 498 4836 554 4892
rect 640 4836 696 4892
rect 498 4694 554 4750
rect 640 4694 696 4750
rect 498 4552 554 4608
rect 640 4552 696 4608
rect 498 4410 554 4466
rect 640 4410 696 4466
rect 498 4268 554 4324
rect 640 4268 696 4324
rect 498 4126 554 4182
rect 640 4126 696 4182
rect 498 3984 554 4040
rect 640 3984 696 4040
rect 498 3860 554 3898
rect 640 3860 696 3898
rect 498 3842 554 3860
rect 640 3842 696 3860
rect 11653 6715 11709 6733
rect 11795 6715 11851 6733
rect 11937 6715 11993 6733
rect 11653 6677 11682 6715
rect 11682 6677 11709 6715
rect 11795 6677 11851 6715
rect 11937 6677 11942 6715
rect 11942 6677 11993 6715
rect 11653 6535 11682 6591
rect 11682 6535 11709 6591
rect 11795 6535 11851 6591
rect 11937 6535 11942 6591
rect 11942 6535 11993 6591
rect 11653 6393 11682 6449
rect 11682 6393 11709 6449
rect 11795 6393 11851 6449
rect 11937 6393 11942 6449
rect 11942 6393 11993 6449
rect 11653 6251 11682 6307
rect 11682 6251 11709 6307
rect 11795 6251 11851 6307
rect 11937 6251 11942 6307
rect 11942 6251 11993 6307
rect 11653 6109 11682 6165
rect 11682 6109 11709 6165
rect 11795 6109 11851 6165
rect 11937 6109 11942 6165
rect 11942 6109 11993 6165
rect 11653 5967 11682 6023
rect 11682 5967 11709 6023
rect 11795 5967 11851 6023
rect 11937 5967 11942 6023
rect 11942 5967 11993 6023
rect 11653 5825 11682 5881
rect 11682 5825 11709 5881
rect 11795 5825 11851 5881
rect 11937 5825 11942 5881
rect 11942 5825 11993 5881
rect 11653 5683 11682 5739
rect 11682 5683 11709 5739
rect 11795 5683 11851 5739
rect 11937 5683 11942 5739
rect 11942 5683 11993 5739
rect 11653 5541 11682 5597
rect 11682 5541 11709 5597
rect 11795 5541 11851 5597
rect 11937 5541 11942 5597
rect 11942 5541 11993 5597
rect 11653 5399 11682 5455
rect 11682 5399 11709 5455
rect 11795 5399 11851 5455
rect 11937 5399 11942 5455
rect 11942 5399 11993 5455
rect 11653 5257 11682 5313
rect 11682 5257 11709 5313
rect 11795 5257 11851 5313
rect 11937 5257 11942 5313
rect 11942 5257 11993 5313
rect 11653 5115 11682 5171
rect 11682 5115 11709 5171
rect 11795 5115 11851 5171
rect 11937 5115 11942 5171
rect 11942 5115 11993 5171
rect 11653 4973 11682 5029
rect 11682 4973 11709 5029
rect 11795 4973 11851 5029
rect 11937 4973 11942 5029
rect 11942 4973 11993 5029
rect 11653 4831 11682 4887
rect 11682 4831 11709 4887
rect 11795 4831 11851 4887
rect 11937 4831 11942 4887
rect 11942 4831 11993 4887
rect 11653 4689 11682 4745
rect 11682 4689 11709 4745
rect 11795 4689 11851 4745
rect 11937 4689 11942 4745
rect 11942 4689 11993 4745
rect 11653 4547 11682 4603
rect 11682 4547 11709 4603
rect 11795 4547 11851 4603
rect 11937 4547 11942 4603
rect 11942 4547 11993 4603
rect 11653 4405 11682 4461
rect 11682 4405 11709 4461
rect 11795 4405 11851 4461
rect 11937 4405 11942 4461
rect 11942 4405 11993 4461
rect 11653 4263 11682 4319
rect 11682 4263 11709 4319
rect 11795 4263 11851 4319
rect 11937 4263 11942 4319
rect 11942 4263 11993 4319
rect 11653 4121 11682 4177
rect 11682 4121 11709 4177
rect 11795 4121 11851 4177
rect 11937 4121 11942 4177
rect 11942 4121 11993 4177
rect 11653 3979 11682 4035
rect 11682 3979 11709 4035
rect 11795 3979 11851 4035
rect 11937 3979 11942 4035
rect 11942 3979 11993 4035
rect 11653 3855 11682 3893
rect 11682 3855 11709 3893
rect 11795 3855 11851 3893
rect 11937 3855 11942 3893
rect 11942 3855 11993 3893
rect 11653 3837 11709 3855
rect 11795 3837 11851 3855
rect 11937 3837 11993 3855
rect 498 3535 554 3553
rect 640 3535 696 3553
rect 498 3497 554 3535
rect 640 3497 696 3535
rect 498 3355 554 3411
rect 640 3355 696 3411
rect 498 3213 554 3269
rect 640 3213 696 3269
rect 498 3071 554 3127
rect 640 3071 696 3127
rect 498 2929 554 2985
rect 640 2929 696 2985
rect 498 2787 554 2843
rect 640 2787 696 2843
rect 498 2645 554 2701
rect 640 2645 696 2701
rect 498 2503 554 2559
rect 640 2503 696 2559
rect 498 2361 554 2417
rect 640 2361 696 2417
rect 498 2219 554 2275
rect 640 2219 696 2275
rect 498 2077 554 2133
rect 640 2077 696 2133
rect 498 1935 554 1991
rect 640 1935 696 1991
rect 498 1793 554 1849
rect 640 1793 696 1849
rect 498 1651 554 1707
rect 640 1651 696 1707
rect 498 1509 554 1565
rect 640 1509 696 1565
rect 498 1367 554 1423
rect 640 1367 696 1423
rect 498 1225 554 1281
rect 640 1225 696 1281
rect 498 1083 554 1139
rect 640 1083 696 1139
rect 498 941 554 997
rect 640 941 696 997
rect 498 799 554 855
rect 640 799 696 855
rect 498 675 554 713
rect 640 675 696 713
rect 498 657 554 675
rect 640 657 696 675
rect 11653 3515 11709 3533
rect 11795 3515 11851 3533
rect 11937 3515 11993 3533
rect 11653 3477 11682 3515
rect 11682 3477 11709 3515
rect 11795 3477 11851 3515
rect 11937 3477 11942 3515
rect 11942 3477 11993 3515
rect 11653 3335 11682 3391
rect 11682 3335 11709 3391
rect 11795 3335 11851 3391
rect 11937 3335 11942 3391
rect 11942 3335 11993 3391
rect 11653 3193 11682 3249
rect 11682 3193 11709 3249
rect 11795 3193 11851 3249
rect 11937 3193 11942 3249
rect 11942 3193 11993 3249
rect 11653 3051 11682 3107
rect 11682 3051 11709 3107
rect 11795 3051 11851 3107
rect 11937 3051 11942 3107
rect 11942 3051 11993 3107
rect 11653 2909 11682 2965
rect 11682 2909 11709 2965
rect 11795 2909 11851 2965
rect 11937 2909 11942 2965
rect 11942 2909 11993 2965
rect 11653 2767 11682 2823
rect 11682 2767 11709 2823
rect 11795 2767 11851 2823
rect 11937 2767 11942 2823
rect 11942 2767 11993 2823
rect 11653 2625 11682 2681
rect 11682 2625 11709 2681
rect 11795 2625 11851 2681
rect 11937 2625 11942 2681
rect 11942 2625 11993 2681
rect 11653 2483 11682 2539
rect 11682 2483 11709 2539
rect 11795 2483 11851 2539
rect 11937 2483 11942 2539
rect 11942 2483 11993 2539
rect 11653 2341 11682 2397
rect 11682 2341 11709 2397
rect 11795 2341 11851 2397
rect 11937 2341 11942 2397
rect 11942 2341 11993 2397
rect 11653 2199 11682 2255
rect 11682 2199 11709 2255
rect 11795 2199 11851 2255
rect 11937 2199 11942 2255
rect 11942 2199 11993 2255
rect 11653 2057 11682 2113
rect 11682 2057 11709 2113
rect 11795 2057 11851 2113
rect 11937 2057 11942 2113
rect 11942 2057 11993 2113
rect 11653 1915 11682 1971
rect 11682 1915 11709 1971
rect 11795 1915 11851 1971
rect 11937 1915 11942 1971
rect 11942 1915 11993 1971
rect 11653 1773 11682 1829
rect 11682 1773 11709 1829
rect 11795 1773 11851 1829
rect 11937 1773 11942 1829
rect 11942 1773 11993 1829
rect 11653 1631 11682 1687
rect 11682 1631 11709 1687
rect 11795 1631 11851 1687
rect 11937 1631 11942 1687
rect 11942 1631 11993 1687
rect 11653 1489 11682 1545
rect 11682 1489 11709 1545
rect 11795 1489 11851 1545
rect 11937 1489 11942 1545
rect 11942 1489 11993 1545
rect 11653 1347 11682 1403
rect 11682 1347 11709 1403
rect 11795 1347 11851 1403
rect 11937 1347 11942 1403
rect 11942 1347 11993 1403
rect 11653 1205 11682 1261
rect 11682 1205 11709 1261
rect 11795 1205 11851 1261
rect 11937 1205 11942 1261
rect 11942 1205 11993 1261
rect 11653 1063 11682 1119
rect 11682 1063 11709 1119
rect 11795 1063 11851 1119
rect 11937 1063 11942 1119
rect 11942 1063 11993 1119
rect 11653 921 11682 977
rect 11682 921 11709 977
rect 11795 921 11851 977
rect 11937 921 11942 977
rect 11942 921 11993 977
rect 11653 779 11682 835
rect 11682 779 11709 835
rect 11795 779 11851 835
rect 11937 779 11942 835
rect 11942 779 11993 835
rect 11653 655 11682 693
rect 11682 655 11709 693
rect 11795 655 11851 693
rect 11937 655 11942 693
rect 11942 655 11993 693
rect 11653 637 11709 655
rect 11795 637 11851 655
rect 11937 637 11993 655
<< metal3 >>
rect 10145 14789 11073 14799
rect -694 14778 -476 14788
rect -694 14722 -684 14778
rect -628 14722 -542 14778
rect -486 14722 -476 14778
rect -694 14636 -476 14722
rect -694 14580 -684 14636
rect -628 14580 -542 14636
rect -486 14580 -476 14636
rect -694 14570 -476 14580
rect 478 14778 838 14788
rect 478 14722 488 14778
rect 544 14722 630 14778
rect 686 14722 772 14778
rect 828 14722 838 14778
rect 478 14636 838 14722
rect 478 14580 488 14636
rect 544 14580 630 14636
rect 686 14580 772 14636
rect 828 14580 838 14636
rect 478 14570 838 14580
rect 1303 14778 2231 14788
rect 1303 14722 1313 14778
rect 1369 14722 1455 14778
rect 1511 14722 1597 14778
rect 1653 14722 1739 14778
rect 1795 14722 1881 14778
rect 1937 14722 2023 14778
rect 2079 14722 2165 14778
rect 2221 14722 2231 14778
rect 1303 14636 2231 14722
rect 1303 14580 1313 14636
rect 1369 14580 1455 14636
rect 1511 14580 1597 14636
rect 1653 14580 1739 14636
rect 1795 14580 1881 14636
rect 1937 14580 2023 14636
rect 2079 14580 2165 14636
rect 2221 14580 2231 14636
rect 1303 14570 2231 14580
rect 3070 14778 3998 14788
rect 3070 14722 3080 14778
rect 3136 14722 3222 14778
rect 3278 14722 3364 14778
rect 3420 14722 3506 14778
rect 3562 14722 3648 14778
rect 3704 14722 3790 14778
rect 3846 14722 3932 14778
rect 3988 14722 3998 14778
rect 3070 14636 3998 14722
rect 3070 14580 3080 14636
rect 3136 14580 3222 14636
rect 3278 14580 3364 14636
rect 3420 14580 3506 14636
rect 3562 14580 3648 14636
rect 3704 14580 3790 14636
rect 3846 14580 3932 14636
rect 3988 14580 3998 14636
rect 3070 14570 3998 14580
rect 4837 14778 5765 14788
rect 4837 14722 4847 14778
rect 4903 14722 4989 14778
rect 5045 14722 5131 14778
rect 5187 14722 5273 14778
rect 5329 14722 5415 14778
rect 5471 14722 5557 14778
rect 5613 14722 5699 14778
rect 5755 14722 5765 14778
rect 4837 14636 5765 14722
rect 4837 14580 4847 14636
rect 4903 14580 4989 14636
rect 5045 14580 5131 14636
rect 5187 14580 5273 14636
rect 5329 14580 5415 14636
rect 5471 14580 5557 14636
rect 5613 14580 5699 14636
rect 5755 14580 5765 14636
rect 4837 14570 5765 14580
rect 6611 14778 7539 14788
rect 6611 14722 6621 14778
rect 6677 14722 6763 14778
rect 6819 14722 6905 14778
rect 6961 14722 7047 14778
rect 7103 14722 7189 14778
rect 7245 14722 7331 14778
rect 7387 14722 7473 14778
rect 7529 14722 7539 14778
rect 6611 14636 7539 14722
rect 6611 14580 6621 14636
rect 6677 14580 6763 14636
rect 6819 14580 6905 14636
rect 6961 14580 7047 14636
rect 7103 14580 7189 14636
rect 7245 14580 7331 14636
rect 7387 14580 7473 14636
rect 7529 14580 7539 14636
rect 6611 14570 7539 14580
rect 8375 14778 9303 14788
rect 8375 14722 8385 14778
rect 8441 14722 8527 14778
rect 8583 14722 8669 14778
rect 8725 14722 8811 14778
rect 8867 14722 8953 14778
rect 9009 14722 9095 14778
rect 9151 14722 9237 14778
rect 9293 14722 9303 14778
rect 8375 14636 9303 14722
rect 8375 14580 8385 14636
rect 8441 14580 8527 14636
rect 8583 14580 8669 14636
rect 8725 14580 8811 14636
rect 8867 14580 8953 14636
rect 9009 14580 9095 14636
rect 9151 14580 9237 14636
rect 9293 14580 9303 14636
rect 10145 14733 10155 14789
rect 10211 14733 10297 14789
rect 10353 14733 10439 14789
rect 10495 14733 10581 14789
rect 10637 14733 10723 14789
rect 10779 14733 10865 14789
rect 10921 14733 11007 14789
rect 11063 14733 11073 14789
rect 10145 14647 11073 14733
rect 10145 14591 10155 14647
rect 10211 14591 10297 14647
rect 10353 14591 10439 14647
rect 10495 14591 10581 14647
rect 10637 14591 10723 14647
rect 10779 14591 10865 14647
rect 10921 14591 11007 14647
rect 11063 14591 11073 14647
rect 10145 14581 11073 14591
rect 11471 14778 11973 14788
rect 11471 14722 11481 14778
rect 11537 14722 11623 14778
rect 11679 14722 11765 14778
rect 11821 14722 11907 14778
rect 11963 14722 11973 14778
rect 11471 14636 11973 14722
rect 8375 14570 9303 14580
rect 11471 14580 11481 14636
rect 11537 14580 11623 14636
rect 11679 14580 11765 14636
rect 11821 14580 11907 14636
rect 11963 14580 11973 14636
rect 11471 14570 11973 14580
rect 488 13138 706 13148
rect 488 13082 498 13138
rect 554 13082 640 13138
rect 696 13082 706 13138
rect 488 12996 706 13082
rect 488 12940 498 12996
rect 554 12940 640 12996
rect 696 12940 706 12996
rect 488 12854 706 12940
rect 488 12798 498 12854
rect 554 12798 640 12854
rect 696 12798 706 12854
rect 488 12712 706 12798
rect 488 12656 498 12712
rect 554 12656 640 12712
rect 696 12656 706 12712
rect 488 12570 706 12656
rect 488 12514 498 12570
rect 554 12514 640 12570
rect 696 12514 706 12570
rect 488 12428 706 12514
rect 488 12372 498 12428
rect 554 12372 640 12428
rect 696 12372 706 12428
rect 488 12286 706 12372
rect 488 12230 498 12286
rect 554 12230 640 12286
rect 696 12230 706 12286
rect 488 12144 706 12230
rect 488 12088 498 12144
rect 554 12088 640 12144
rect 696 12088 706 12144
rect 488 12002 706 12088
rect 488 11946 498 12002
rect 554 11946 640 12002
rect 696 11946 706 12002
rect 488 11860 706 11946
rect 488 11804 498 11860
rect 554 11804 640 11860
rect 696 11804 706 11860
rect 488 11718 706 11804
rect 488 11662 498 11718
rect 554 11662 640 11718
rect 696 11662 706 11718
rect 488 11576 706 11662
rect 488 11520 498 11576
rect 554 11520 640 11576
rect 696 11520 706 11576
rect 488 11434 706 11520
rect 488 11378 498 11434
rect 554 11378 640 11434
rect 696 11378 706 11434
rect 488 11292 706 11378
rect 488 11236 498 11292
rect 554 11236 640 11292
rect 696 11236 706 11292
rect 488 11150 706 11236
rect 488 11094 498 11150
rect 554 11094 640 11150
rect 696 11094 706 11150
rect 488 11008 706 11094
rect 488 10952 498 11008
rect 554 10952 640 11008
rect 696 10952 706 11008
rect 488 10866 706 10952
rect 488 10810 498 10866
rect 554 10810 640 10866
rect 696 10810 706 10866
rect 488 10724 706 10810
rect 488 10668 498 10724
rect 554 10668 640 10724
rect 696 10668 706 10724
rect 488 10582 706 10668
rect 488 10526 498 10582
rect 554 10526 640 10582
rect 696 10526 706 10582
rect 488 10440 706 10526
rect 488 10384 498 10440
rect 554 10384 640 10440
rect 696 10384 706 10440
rect 488 10298 706 10384
rect 488 10242 498 10298
rect 554 10242 640 10298
rect 696 10242 706 10298
rect 488 10232 706 10242
rect 11643 13133 12003 13143
rect 11643 13077 11653 13133
rect 11709 13077 11795 13133
rect 11851 13077 11937 13133
rect 11993 13077 12003 13133
rect 11643 12991 12003 13077
rect 11643 12935 11653 12991
rect 11709 12935 11795 12991
rect 11851 12935 11937 12991
rect 11993 12935 12003 12991
rect 11643 12849 12003 12935
rect 11643 12793 11653 12849
rect 11709 12793 11795 12849
rect 11851 12793 11937 12849
rect 11993 12793 12003 12849
rect 11643 12707 12003 12793
rect 11643 12651 11653 12707
rect 11709 12651 11795 12707
rect 11851 12651 11937 12707
rect 11993 12651 12003 12707
rect 11643 12565 12003 12651
rect 11643 12509 11653 12565
rect 11709 12509 11795 12565
rect 11851 12509 11937 12565
rect 11993 12509 12003 12565
rect 11643 12423 12003 12509
rect 11643 12367 11653 12423
rect 11709 12367 11795 12423
rect 11851 12367 11937 12423
rect 11993 12367 12003 12423
rect 11643 12281 12003 12367
rect 11643 12225 11653 12281
rect 11709 12225 11795 12281
rect 11851 12225 11937 12281
rect 11993 12225 12003 12281
rect 11643 12139 12003 12225
rect 11643 12083 11653 12139
rect 11709 12083 11795 12139
rect 11851 12083 11937 12139
rect 11993 12083 12003 12139
rect 11643 11997 12003 12083
rect 11643 11941 11653 11997
rect 11709 11941 11795 11997
rect 11851 11941 11937 11997
rect 11993 11941 12003 11997
rect 11643 11855 12003 11941
rect 11643 11799 11653 11855
rect 11709 11799 11795 11855
rect 11851 11799 11937 11855
rect 11993 11799 12003 11855
rect 11643 11713 12003 11799
rect 11643 11657 11653 11713
rect 11709 11657 11795 11713
rect 11851 11657 11937 11713
rect 11993 11657 12003 11713
rect 11643 11571 12003 11657
rect 11643 11515 11653 11571
rect 11709 11515 11795 11571
rect 11851 11515 11937 11571
rect 11993 11515 12003 11571
rect 11643 11429 12003 11515
rect 11643 11373 11653 11429
rect 11709 11373 11795 11429
rect 11851 11373 11937 11429
rect 11993 11373 12003 11429
rect 11643 11287 12003 11373
rect 11643 11231 11653 11287
rect 11709 11231 11795 11287
rect 11851 11231 11937 11287
rect 11993 11231 12003 11287
rect 11643 11145 12003 11231
rect 11643 11089 11653 11145
rect 11709 11089 11795 11145
rect 11851 11089 11937 11145
rect 11993 11089 12003 11145
rect 11643 11003 12003 11089
rect 11643 10947 11653 11003
rect 11709 10947 11795 11003
rect 11851 10947 11937 11003
rect 11993 10947 12003 11003
rect 11643 10861 12003 10947
rect 11643 10805 11653 10861
rect 11709 10805 11795 10861
rect 11851 10805 11937 10861
rect 11993 10805 12003 10861
rect 11643 10719 12003 10805
rect 11643 10663 11653 10719
rect 11709 10663 11795 10719
rect 11851 10663 11937 10719
rect 11993 10663 12003 10719
rect 11643 10577 12003 10663
rect 11643 10521 11653 10577
rect 11709 10521 11795 10577
rect 11851 10521 11937 10577
rect 11993 10521 12003 10577
rect 11643 10435 12003 10521
rect 11643 10379 11653 10435
rect 11709 10379 11795 10435
rect 11851 10379 11937 10435
rect 11993 10379 12003 10435
rect 11643 10293 12003 10379
rect 11643 10237 11653 10293
rect 11709 10237 11795 10293
rect 11851 10237 11937 10293
rect 11993 10237 12003 10293
rect 11643 10227 12003 10237
rect 488 9938 706 9948
rect 488 9882 498 9938
rect 554 9882 640 9938
rect 696 9882 706 9938
rect 488 9796 706 9882
rect 488 9740 498 9796
rect 554 9740 640 9796
rect 696 9740 706 9796
rect 488 9654 706 9740
rect 488 9598 498 9654
rect 554 9598 640 9654
rect 696 9598 706 9654
rect 488 9512 706 9598
rect 488 9456 498 9512
rect 554 9456 640 9512
rect 696 9456 706 9512
rect 488 9370 706 9456
rect 488 9314 498 9370
rect 554 9314 640 9370
rect 696 9314 706 9370
rect 488 9228 706 9314
rect 488 9172 498 9228
rect 554 9172 640 9228
rect 696 9172 706 9228
rect 488 9086 706 9172
rect 488 9030 498 9086
rect 554 9030 640 9086
rect 696 9030 706 9086
rect 488 8944 706 9030
rect 488 8888 498 8944
rect 554 8888 640 8944
rect 696 8888 706 8944
rect 488 8802 706 8888
rect 488 8746 498 8802
rect 554 8746 640 8802
rect 696 8746 706 8802
rect 488 8660 706 8746
rect 488 8604 498 8660
rect 554 8604 640 8660
rect 696 8604 706 8660
rect 488 8518 706 8604
rect 488 8462 498 8518
rect 554 8462 640 8518
rect 696 8462 706 8518
rect 488 8376 706 8462
rect 488 8320 498 8376
rect 554 8320 640 8376
rect 696 8320 706 8376
rect 488 8234 706 8320
rect 488 8178 498 8234
rect 554 8178 640 8234
rect 696 8178 706 8234
rect 488 8092 706 8178
rect 488 8036 498 8092
rect 554 8036 640 8092
rect 696 8036 706 8092
rect 488 7950 706 8036
rect 488 7894 498 7950
rect 554 7894 640 7950
rect 696 7894 706 7950
rect 488 7808 706 7894
rect 488 7752 498 7808
rect 554 7752 640 7808
rect 696 7752 706 7808
rect 488 7666 706 7752
rect 488 7610 498 7666
rect 554 7610 640 7666
rect 696 7610 706 7666
rect 488 7524 706 7610
rect 488 7468 498 7524
rect 554 7468 640 7524
rect 696 7468 706 7524
rect 488 7382 706 7468
rect 488 7326 498 7382
rect 554 7326 640 7382
rect 696 7326 706 7382
rect 488 7240 706 7326
rect 488 7184 498 7240
rect 554 7184 640 7240
rect 696 7184 706 7240
rect 488 7098 706 7184
rect 488 7042 498 7098
rect 554 7042 640 7098
rect 696 7042 706 7098
rect 488 7032 706 7042
rect 11643 9933 12003 9943
rect 11643 9877 11653 9933
rect 11709 9877 11795 9933
rect 11851 9877 11937 9933
rect 11993 9877 12003 9933
rect 11643 9791 12003 9877
rect 11643 9735 11653 9791
rect 11709 9735 11795 9791
rect 11851 9735 11937 9791
rect 11993 9735 12003 9791
rect 11643 9649 12003 9735
rect 11643 9593 11653 9649
rect 11709 9593 11795 9649
rect 11851 9593 11937 9649
rect 11993 9593 12003 9649
rect 11643 9507 12003 9593
rect 11643 9451 11653 9507
rect 11709 9451 11795 9507
rect 11851 9451 11937 9507
rect 11993 9451 12003 9507
rect 11643 9365 12003 9451
rect 11643 9309 11653 9365
rect 11709 9309 11795 9365
rect 11851 9309 11937 9365
rect 11993 9309 12003 9365
rect 11643 9223 12003 9309
rect 11643 9167 11653 9223
rect 11709 9167 11795 9223
rect 11851 9167 11937 9223
rect 11993 9167 12003 9223
rect 11643 9081 12003 9167
rect 11643 9025 11653 9081
rect 11709 9025 11795 9081
rect 11851 9025 11937 9081
rect 11993 9025 12003 9081
rect 11643 8939 12003 9025
rect 11643 8883 11653 8939
rect 11709 8883 11795 8939
rect 11851 8883 11937 8939
rect 11993 8883 12003 8939
rect 11643 8797 12003 8883
rect 11643 8741 11653 8797
rect 11709 8741 11795 8797
rect 11851 8741 11937 8797
rect 11993 8741 12003 8797
rect 11643 8655 12003 8741
rect 11643 8599 11653 8655
rect 11709 8599 11795 8655
rect 11851 8599 11937 8655
rect 11993 8599 12003 8655
rect 11643 8513 12003 8599
rect 11643 8457 11653 8513
rect 11709 8457 11795 8513
rect 11851 8457 11937 8513
rect 11993 8457 12003 8513
rect 11643 8371 12003 8457
rect 11643 8315 11653 8371
rect 11709 8315 11795 8371
rect 11851 8315 11937 8371
rect 11993 8315 12003 8371
rect 11643 8229 12003 8315
rect 11643 8173 11653 8229
rect 11709 8173 11795 8229
rect 11851 8173 11937 8229
rect 11993 8173 12003 8229
rect 11643 8087 12003 8173
rect 11643 8031 11653 8087
rect 11709 8031 11795 8087
rect 11851 8031 11937 8087
rect 11993 8031 12003 8087
rect 11643 7945 12003 8031
rect 11643 7889 11653 7945
rect 11709 7889 11795 7945
rect 11851 7889 11937 7945
rect 11993 7889 12003 7945
rect 11643 7803 12003 7889
rect 11643 7747 11653 7803
rect 11709 7747 11795 7803
rect 11851 7747 11937 7803
rect 11993 7747 12003 7803
rect 11643 7661 12003 7747
rect 11643 7605 11653 7661
rect 11709 7605 11795 7661
rect 11851 7605 11937 7661
rect 11993 7605 12003 7661
rect 11643 7519 12003 7605
rect 11643 7463 11653 7519
rect 11709 7463 11795 7519
rect 11851 7463 11937 7519
rect 11993 7463 12003 7519
rect 11643 7377 12003 7463
rect 11643 7321 11653 7377
rect 11709 7321 11795 7377
rect 11851 7321 11937 7377
rect 11993 7321 12003 7377
rect 11643 7235 12003 7321
rect 11643 7179 11653 7235
rect 11709 7179 11795 7235
rect 11851 7179 11937 7235
rect 11993 7179 12003 7235
rect 11643 7093 12003 7179
rect 11643 7037 11653 7093
rect 11709 7037 11795 7093
rect 11851 7037 11937 7093
rect 11993 7037 12003 7093
rect 11643 7027 12003 7037
rect 488 6738 706 6748
rect 488 6682 498 6738
rect 554 6682 640 6738
rect 696 6682 706 6738
rect 488 6596 706 6682
rect 488 6540 498 6596
rect 554 6540 640 6596
rect 696 6540 706 6596
rect 488 6454 706 6540
rect 488 6398 498 6454
rect 554 6398 640 6454
rect 696 6398 706 6454
rect 488 6312 706 6398
rect 488 6256 498 6312
rect 554 6256 640 6312
rect 696 6256 706 6312
rect 488 6170 706 6256
rect 488 6114 498 6170
rect 554 6114 640 6170
rect 696 6114 706 6170
rect 488 6028 706 6114
rect 488 5972 498 6028
rect 554 5972 640 6028
rect 696 5972 706 6028
rect 488 5886 706 5972
rect 488 5830 498 5886
rect 554 5830 640 5886
rect 696 5830 706 5886
rect 488 5744 706 5830
rect 488 5688 498 5744
rect 554 5688 640 5744
rect 696 5688 706 5744
rect 488 5602 706 5688
rect 488 5546 498 5602
rect 554 5546 640 5602
rect 696 5546 706 5602
rect 488 5460 706 5546
rect 488 5404 498 5460
rect 554 5404 640 5460
rect 696 5404 706 5460
rect 488 5318 706 5404
rect 488 5262 498 5318
rect 554 5262 640 5318
rect 696 5262 706 5318
rect 488 5176 706 5262
rect 488 5120 498 5176
rect 554 5120 640 5176
rect 696 5120 706 5176
rect 488 5034 706 5120
rect 488 4978 498 5034
rect 554 4978 640 5034
rect 696 4978 706 5034
rect 488 4892 706 4978
rect 488 4836 498 4892
rect 554 4836 640 4892
rect 696 4836 706 4892
rect 488 4750 706 4836
rect 488 4694 498 4750
rect 554 4694 640 4750
rect 696 4694 706 4750
rect 488 4608 706 4694
rect 488 4552 498 4608
rect 554 4552 640 4608
rect 696 4552 706 4608
rect 488 4466 706 4552
rect 488 4410 498 4466
rect 554 4410 640 4466
rect 696 4410 706 4466
rect 488 4324 706 4410
rect 488 4268 498 4324
rect 554 4268 640 4324
rect 696 4268 706 4324
rect 488 4182 706 4268
rect 488 4126 498 4182
rect 554 4126 640 4182
rect 696 4126 706 4182
rect 488 4040 706 4126
rect 488 3984 498 4040
rect 554 3984 640 4040
rect 696 3984 706 4040
rect 488 3898 706 3984
rect 488 3842 498 3898
rect 554 3842 640 3898
rect 696 3842 706 3898
rect 488 3832 706 3842
rect 11643 6733 12003 6743
rect 11643 6677 11653 6733
rect 11709 6677 11795 6733
rect 11851 6677 11937 6733
rect 11993 6677 12003 6733
rect 11643 6591 12003 6677
rect 11643 6535 11653 6591
rect 11709 6535 11795 6591
rect 11851 6535 11937 6591
rect 11993 6535 12003 6591
rect 11643 6449 12003 6535
rect 11643 6393 11653 6449
rect 11709 6393 11795 6449
rect 11851 6393 11937 6449
rect 11993 6393 12003 6449
rect 11643 6307 12003 6393
rect 11643 6251 11653 6307
rect 11709 6251 11795 6307
rect 11851 6251 11937 6307
rect 11993 6251 12003 6307
rect 11643 6165 12003 6251
rect 11643 6109 11653 6165
rect 11709 6109 11795 6165
rect 11851 6109 11937 6165
rect 11993 6109 12003 6165
rect 11643 6023 12003 6109
rect 11643 5967 11653 6023
rect 11709 5967 11795 6023
rect 11851 5967 11937 6023
rect 11993 5967 12003 6023
rect 11643 5881 12003 5967
rect 11643 5825 11653 5881
rect 11709 5825 11795 5881
rect 11851 5825 11937 5881
rect 11993 5825 12003 5881
rect 11643 5739 12003 5825
rect 11643 5683 11653 5739
rect 11709 5683 11795 5739
rect 11851 5683 11937 5739
rect 11993 5683 12003 5739
rect 11643 5597 12003 5683
rect 11643 5541 11653 5597
rect 11709 5541 11795 5597
rect 11851 5541 11937 5597
rect 11993 5541 12003 5597
rect 11643 5455 12003 5541
rect 11643 5399 11653 5455
rect 11709 5399 11795 5455
rect 11851 5399 11937 5455
rect 11993 5399 12003 5455
rect 11643 5313 12003 5399
rect 11643 5257 11653 5313
rect 11709 5257 11795 5313
rect 11851 5257 11937 5313
rect 11993 5257 12003 5313
rect 11643 5171 12003 5257
rect 11643 5115 11653 5171
rect 11709 5115 11795 5171
rect 11851 5115 11937 5171
rect 11993 5115 12003 5171
rect 11643 5029 12003 5115
rect 11643 4973 11653 5029
rect 11709 4973 11795 5029
rect 11851 4973 11937 5029
rect 11993 4973 12003 5029
rect 11643 4887 12003 4973
rect 11643 4831 11653 4887
rect 11709 4831 11795 4887
rect 11851 4831 11937 4887
rect 11993 4831 12003 4887
rect 11643 4745 12003 4831
rect 11643 4689 11653 4745
rect 11709 4689 11795 4745
rect 11851 4689 11937 4745
rect 11993 4689 12003 4745
rect 11643 4603 12003 4689
rect 11643 4547 11653 4603
rect 11709 4547 11795 4603
rect 11851 4547 11937 4603
rect 11993 4547 12003 4603
rect 11643 4461 12003 4547
rect 11643 4405 11653 4461
rect 11709 4405 11795 4461
rect 11851 4405 11937 4461
rect 11993 4405 12003 4461
rect 11643 4319 12003 4405
rect 11643 4263 11653 4319
rect 11709 4263 11795 4319
rect 11851 4263 11937 4319
rect 11993 4263 12003 4319
rect 11643 4177 12003 4263
rect 11643 4121 11653 4177
rect 11709 4121 11795 4177
rect 11851 4121 11937 4177
rect 11993 4121 12003 4177
rect 11643 4035 12003 4121
rect 11643 3979 11653 4035
rect 11709 3979 11795 4035
rect 11851 3979 11937 4035
rect 11993 3979 12003 4035
rect 11643 3893 12003 3979
rect 11643 3837 11653 3893
rect 11709 3837 11795 3893
rect 11851 3837 11937 3893
rect 11993 3837 12003 3893
rect 11643 3827 12003 3837
rect 488 3553 706 3563
rect 488 3497 498 3553
rect 554 3497 640 3553
rect 696 3497 706 3553
rect 488 3411 706 3497
rect 488 3355 498 3411
rect 554 3355 640 3411
rect 696 3355 706 3411
rect 488 3269 706 3355
rect 488 3213 498 3269
rect 554 3213 640 3269
rect 696 3213 706 3269
rect 488 3127 706 3213
rect 488 3071 498 3127
rect 554 3071 640 3127
rect 696 3071 706 3127
rect 488 2985 706 3071
rect 488 2929 498 2985
rect 554 2929 640 2985
rect 696 2929 706 2985
rect 488 2843 706 2929
rect 488 2787 498 2843
rect 554 2787 640 2843
rect 696 2787 706 2843
rect 488 2701 706 2787
rect 488 2645 498 2701
rect 554 2645 640 2701
rect 696 2645 706 2701
rect 488 2559 706 2645
rect 488 2503 498 2559
rect 554 2503 640 2559
rect 696 2503 706 2559
rect 488 2417 706 2503
rect 488 2361 498 2417
rect 554 2361 640 2417
rect 696 2361 706 2417
rect 488 2275 706 2361
rect 488 2219 498 2275
rect 554 2219 640 2275
rect 696 2219 706 2275
rect 488 2133 706 2219
rect 488 2077 498 2133
rect 554 2077 640 2133
rect 696 2077 706 2133
rect 488 1991 706 2077
rect 488 1935 498 1991
rect 554 1935 640 1991
rect 696 1935 706 1991
rect 488 1849 706 1935
rect 488 1793 498 1849
rect 554 1793 640 1849
rect 696 1793 706 1849
rect 488 1707 706 1793
rect 488 1651 498 1707
rect 554 1651 640 1707
rect 696 1651 706 1707
rect 488 1565 706 1651
rect 488 1509 498 1565
rect 554 1509 640 1565
rect 696 1509 706 1565
rect 488 1423 706 1509
rect 488 1367 498 1423
rect 554 1367 640 1423
rect 696 1367 706 1423
rect 488 1281 706 1367
rect 488 1225 498 1281
rect 554 1225 640 1281
rect 696 1225 706 1281
rect 488 1139 706 1225
rect 488 1083 498 1139
rect 554 1083 640 1139
rect 696 1083 706 1139
rect 488 997 706 1083
rect 488 941 498 997
rect 554 941 640 997
rect 696 941 706 997
rect 488 855 706 941
rect 488 799 498 855
rect 554 799 640 855
rect 696 799 706 855
rect 488 713 706 799
rect 488 657 498 713
rect 554 657 640 713
rect 696 657 706 713
rect 488 647 706 657
rect 11643 3533 12003 3543
rect 11643 3477 11653 3533
rect 11709 3477 11795 3533
rect 11851 3477 11937 3533
rect 11993 3477 12003 3533
rect 11643 3391 12003 3477
rect 11643 3335 11653 3391
rect 11709 3335 11795 3391
rect 11851 3335 11937 3391
rect 11993 3335 12003 3391
rect 11643 3249 12003 3335
rect 11643 3193 11653 3249
rect 11709 3193 11795 3249
rect 11851 3193 11937 3249
rect 11993 3193 12003 3249
rect 11643 3107 12003 3193
rect 11643 3051 11653 3107
rect 11709 3051 11795 3107
rect 11851 3051 11937 3107
rect 11993 3051 12003 3107
rect 11643 2965 12003 3051
rect 11643 2909 11653 2965
rect 11709 2909 11795 2965
rect 11851 2909 11937 2965
rect 11993 2909 12003 2965
rect 11643 2823 12003 2909
rect 11643 2767 11653 2823
rect 11709 2767 11795 2823
rect 11851 2767 11937 2823
rect 11993 2767 12003 2823
rect 11643 2681 12003 2767
rect 11643 2625 11653 2681
rect 11709 2625 11795 2681
rect 11851 2625 11937 2681
rect 11993 2625 12003 2681
rect 11643 2539 12003 2625
rect 11643 2483 11653 2539
rect 11709 2483 11795 2539
rect 11851 2483 11937 2539
rect 11993 2483 12003 2539
rect 11643 2397 12003 2483
rect 11643 2341 11653 2397
rect 11709 2341 11795 2397
rect 11851 2341 11937 2397
rect 11993 2341 12003 2397
rect 11643 2255 12003 2341
rect 11643 2199 11653 2255
rect 11709 2199 11795 2255
rect 11851 2199 11937 2255
rect 11993 2199 12003 2255
rect 11643 2113 12003 2199
rect 11643 2057 11653 2113
rect 11709 2057 11795 2113
rect 11851 2057 11937 2113
rect 11993 2057 12003 2113
rect 11643 1971 12003 2057
rect 11643 1915 11653 1971
rect 11709 1915 11795 1971
rect 11851 1915 11937 1971
rect 11993 1915 12003 1971
rect 11643 1829 12003 1915
rect 11643 1773 11653 1829
rect 11709 1773 11795 1829
rect 11851 1773 11937 1829
rect 11993 1773 12003 1829
rect 11643 1687 12003 1773
rect 11643 1631 11653 1687
rect 11709 1631 11795 1687
rect 11851 1631 11937 1687
rect 11993 1631 12003 1687
rect 11643 1545 12003 1631
rect 11643 1489 11653 1545
rect 11709 1489 11795 1545
rect 11851 1489 11937 1545
rect 11993 1489 12003 1545
rect 11643 1403 12003 1489
rect 11643 1347 11653 1403
rect 11709 1347 11795 1403
rect 11851 1347 11937 1403
rect 11993 1347 12003 1403
rect 11643 1261 12003 1347
rect 11643 1205 11653 1261
rect 11709 1205 11795 1261
rect 11851 1205 11937 1261
rect 11993 1205 12003 1261
rect 11643 1119 12003 1205
rect 11643 1063 11653 1119
rect 11709 1063 11795 1119
rect 11851 1063 11937 1119
rect 11993 1063 12003 1119
rect 11643 977 12003 1063
rect 11643 921 11653 977
rect 11709 921 11795 977
rect 11851 921 11937 977
rect 11993 921 12003 977
rect 11643 835 12003 921
rect 11643 779 11653 835
rect 11709 779 11795 835
rect 11851 779 11937 835
rect 11993 779 12003 835
rect 11643 693 12003 779
rect 11643 637 11653 693
rect 11709 637 11795 693
rect 11851 637 11937 693
rect 11993 637 12003 693
rect 11643 627 12003 637
use comp018green_out_drv_pleg_6T_X  comp018green_out_drv_pleg_6T_X_0
timestamp 1758724778
transform -1 0 11651 0 1 364
box 0 12 2080 12252
use comp018green_out_drv_pleg_6T_X  comp018green_out_drv_pleg_6T_X_1
timestamp 1758724778
transform -1 0 6347 0 1 364
box 0 12 2080 12252
use comp018green_out_drv_pleg_6T_X  comp018green_out_drv_pleg_6T_X_2
timestamp 1758724778
transform 1 0 6035 0 1 364
box 0 12 2080 12252
use comp018green_out_drv_pleg_6T_X  comp018green_out_drv_pleg_6T_X_3
timestamp 1758724778
transform 1 0 731 0 1 364
box 0 12 2080 12252
use comp018green_out_drv_pleg_6T_Y  comp018green_out_drv_pleg_6T_Y_0
timestamp 1758724778
transform -1 0 9883 0 1 364
box 0 12 1196 12252
use comp018green_out_drv_pleg_6T_Y  comp018green_out_drv_pleg_6T_Y_1
timestamp 1758724778
transform -1 0 4579 0 1 364
box 0 12 1196 12252
use comp018green_out_drv_pleg_6T_Y  comp018green_out_drv_pleg_6T_Y_2
timestamp 1758724778
transform 1 0 7803 0 1 364
box 0 12 1196 12252
use comp018green_out_drv_pleg_6T_Y  comp018green_out_drv_pleg_6T_Y_3
timestamp 1758724778
transform 1 0 2499 0 1 364
box 0 12 1196 12252
use PMOS_metal_stack  PMOS_metal_stack_0
timestamp 1758724778
transform -1 0 11573 0 1 496
box -44 0 1584 12000
use PMOS_metal_stack  PMOS_metal_stack_1
timestamp 1758724778
transform 1 0 9649 0 1 496
box -44 0 1584 12000
use PMOS_metal_stack  PMOS_metal_stack_2
timestamp 1758724778
transform 1 0 6113 0 1 496
box -44 0 1584 12000
use PMOS_metal_stack  PMOS_metal_stack_3
timestamp 1758724778
transform 1 0 7881 0 1 496
box -44 0 1584 12000
use PMOS_metal_stack  PMOS_metal_stack_4
timestamp 1758724778
transform 1 0 4345 0 1 496
box -44 0 1584 12000
use PMOS_metal_stack  PMOS_metal_stack_5
timestamp 1758724778
transform 1 0 2577 0 1 496
box -44 0 1584 12000
use PMOS_metal_stack  PMOS_metal_stack_6
timestamp 1758724778
transform 1 0 809 0 1 496
box -44 0 1584 12000
<< end >>
