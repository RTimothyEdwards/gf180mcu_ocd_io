magic
tech gf180mcuD
magscale 1 10
timestamp 1484609607
<< metal4 >>
rect 118 64944 298 64954
rect 118 64888 128 64944
rect 288 64888 298 64944
rect 118 64832 298 64888
rect 118 64776 128 64832
rect 288 64776 298 64832
rect 118 64720 298 64776
rect 118 64664 128 64720
rect 288 64664 298 64720
rect 118 64608 298 64664
rect 118 64552 128 64608
rect 288 64552 298 64608
rect 118 64496 298 64552
rect 118 64440 128 64496
rect 288 64440 298 64496
rect 118 64384 298 64440
rect 118 64328 128 64384
rect 288 64328 298 64384
rect 118 64272 298 64328
rect 118 64216 128 64272
rect 288 64216 298 64272
rect 118 64160 298 64216
rect 118 64104 128 64160
rect 288 64104 298 64160
rect 118 64048 298 64104
rect 118 63992 128 64048
rect 288 63992 298 64048
rect 118 63936 298 63992
rect 118 63880 128 63936
rect 288 63880 298 63936
rect 118 63824 298 63880
rect 118 63768 128 63824
rect 288 63768 298 63824
rect 118 63712 298 63768
rect 118 63656 128 63712
rect 288 63656 298 63712
rect 118 63646 298 63656
rect 115 50538 303 50548
rect 115 50482 125 50538
rect 181 50482 237 50538
rect 293 50482 303 50538
rect 115 50426 303 50482
rect 115 50370 125 50426
rect 181 50370 237 50426
rect 293 50370 303 50426
rect 115 50314 303 50370
rect 115 50258 125 50314
rect 181 50258 237 50314
rect 293 50258 303 50314
rect 115 50202 303 50258
rect 115 50146 125 50202
rect 181 50146 237 50202
rect 293 50146 303 50202
rect 115 50090 303 50146
rect 115 50034 125 50090
rect 181 50034 237 50090
rect 293 50034 303 50090
rect 115 49978 303 50034
rect 115 49922 125 49978
rect 181 49922 237 49978
rect 293 49922 303 49978
rect 115 49866 303 49922
rect 115 49810 125 49866
rect 181 49810 237 49866
rect 293 49810 303 49866
rect 115 49754 303 49810
rect 115 49698 125 49754
rect 181 49698 237 49754
rect 293 49698 303 49754
rect 115 49642 303 49698
rect 115 49586 125 49642
rect 181 49586 237 49642
rect 293 49586 303 49642
rect 115 49530 303 49586
rect 115 49474 125 49530
rect 181 49474 237 49530
rect 293 49474 303 49530
rect 115 49418 303 49474
rect 115 49362 125 49418
rect 181 49362 237 49418
rect 293 49362 303 49418
rect 115 49306 303 49362
rect 115 49250 125 49306
rect 181 49250 237 49306
rect 293 49250 303 49306
rect 115 49240 303 49250
<< via4 >>
rect 128 64888 288 64944
rect 128 64776 288 64832
rect 128 64664 288 64720
rect 128 64552 288 64608
rect 128 64440 288 64496
rect 128 64328 288 64384
rect 128 64216 288 64272
rect 128 64104 288 64160
rect 128 63992 288 64048
rect 128 63880 288 63936
rect 128 63768 288 63824
rect 128 63656 288 63712
rect 125 50482 181 50538
rect 237 50482 293 50538
rect 125 50370 181 50426
rect 237 50370 293 50426
rect 125 50258 181 50314
rect 237 50258 293 50314
rect 125 50146 181 50202
rect 237 50146 293 50202
rect 125 50034 181 50090
rect 237 50034 293 50090
rect 125 49922 181 49978
rect 237 49922 293 49978
rect 125 49810 181 49866
rect 237 49810 293 49866
rect 125 49698 181 49754
rect 237 49698 293 49754
rect 125 49586 181 49642
rect 237 49586 293 49642
rect 125 49474 181 49530
rect 237 49474 293 49530
rect 125 49362 181 49418
rect 237 49362 293 49418
rect 125 49250 181 49306
rect 237 49250 293 49306
<< metal5 >>
rect 0 64944 400 65000
rect 0 64888 128 64944
rect 288 64888 400 64944
rect 0 64832 400 64888
rect 0 64776 128 64832
rect 288 64776 400 64832
rect 0 64720 400 64776
rect 0 64664 128 64720
rect 288 64664 400 64720
rect 0 64608 400 64664
rect 0 64552 128 64608
rect 288 64552 400 64608
rect 0 64496 400 64552
rect 0 64440 128 64496
rect 288 64440 400 64496
rect 0 64384 400 64440
rect 0 64328 128 64384
rect 288 64328 400 64384
rect 0 64272 400 64328
rect 0 64216 128 64272
rect 288 64216 400 64272
rect 0 64160 400 64216
rect 0 64104 128 64160
rect 288 64104 400 64160
rect 0 64048 400 64104
rect 0 63992 128 64048
rect 288 63992 400 64048
rect 0 63936 400 63992
rect 0 63880 128 63936
rect 288 63880 400 63936
rect 0 63824 400 63880
rect 0 63768 128 63824
rect 288 63768 400 63824
rect 0 63712 400 63768
rect 0 63656 128 63712
rect 288 63656 400 63712
rect 0 63600 400 63656
rect 0 50538 400 50600
rect 0 50482 125 50538
rect 181 50482 237 50538
rect 293 50482 400 50538
rect 0 50426 400 50482
rect 0 50370 125 50426
rect 181 50370 237 50426
rect 293 50370 400 50426
rect 0 50314 400 50370
rect 0 50258 125 50314
rect 181 50258 237 50314
rect 293 50258 400 50314
rect 0 50202 400 50258
rect 0 50146 125 50202
rect 181 50146 237 50202
rect 293 50146 400 50202
rect 0 50090 400 50146
rect 0 50034 125 50090
rect 181 50034 237 50090
rect 293 50034 400 50090
rect 0 49978 400 50034
rect 0 49922 125 49978
rect 181 49922 237 49978
rect 293 49922 400 49978
rect 0 49866 400 49922
rect 0 49810 125 49866
rect 181 49810 237 49866
rect 293 49810 400 49866
rect 0 49754 400 49810
rect 0 49698 125 49754
rect 181 49698 237 49754
rect 293 49698 400 49754
rect 0 49642 400 49698
rect 0 49586 125 49642
rect 181 49586 237 49642
rect 293 49586 400 49642
rect 0 49530 400 49586
rect 0 49474 125 49530
rect 181 49474 237 49530
rect 293 49474 400 49530
rect 0 49418 400 49474
rect 0 49362 125 49418
rect 181 49362 237 49418
rect 293 49362 400 49418
rect 0 49306 400 49362
rect 0 49250 125 49306
rect 181 49250 237 49306
rect 293 49250 400 49306
rect 0 49200 400 49250
use GF_NI_BRK2_0  GF_NI_BRK2_0_0
timestamp 1484609607
transform 1 0 0 0 1 0
box -32 13097 432 69968
<< labels >>
rlabel metal3 s 207 64258 207 64258 4 VSS
port 1 nsew
rlabel metal3 s 208 50023 208 50023 4 VSS
port 1 nsew
rlabel metal4 s 207 64258 207 64258 4 VSS
port 1 nsew
rlabel metal4 s 208 50023 208 50023 4 VSS
port 1 nsew
rlabel metal5 s 207 64258 207 64258 4 VSS
port 1 nsew
rlabel metal5 s 208 50023 208 50023 4 VSS
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 400 70000
<< end >>
