magic
tech gf180mcuD
magscale 1 10
timestamp 1758892345
<< isosubstrate >>
rect -496 -83 2202 2575
<< nwell >>
rect -247 1551 2202 2575
rect 633 1281 2202 1551
rect 2741 1281 4189 2004
<< nmos >>
rect 3011 747 3067 867
rect 3175 747 3231 867
rect 3339 747 3395 867
rect 3503 747 3559 867
rect 3667 747 3723 867
rect 3831 747 3887 867
<< pmos >>
rect 3011 1523 3067 1803
rect 3175 1523 3231 1803
rect 3339 1523 3395 1803
rect 3503 1523 3559 1803
rect 3667 1523 3723 1803
rect 3831 1523 3887 1803
<< mvnmos >>
rect -92 263 48 1063
rect 152 263 292 1063
rect 1255 270 1395 520
rect 1499 270 1639 520
<< mvpmos >>
rect 152 1811 292 2211
rect 1011 1522 1151 2022
rect 1255 1522 1395 2022
rect 1499 1522 1639 2022
rect 1743 1522 1883 2022
<< ndiff >>
rect 2919 854 3011 867
rect 2919 760 2932 854
rect 2982 760 3011 854
rect 2919 747 3011 760
rect 3067 854 3175 867
rect 3067 760 3096 854
rect 3146 760 3175 854
rect 3067 747 3175 760
rect 3231 854 3339 867
rect 3231 760 3260 854
rect 3310 760 3339 854
rect 3231 747 3339 760
rect 3395 854 3503 867
rect 3395 760 3424 854
rect 3474 760 3503 854
rect 3395 747 3503 760
rect 3559 854 3667 867
rect 3559 760 3588 854
rect 3638 760 3667 854
rect 3559 747 3667 760
rect 3723 854 3831 867
rect 3723 760 3752 854
rect 3802 760 3831 854
rect 3723 747 3831 760
rect 3887 854 3979 867
rect 3887 760 3916 854
rect 3966 760 3979 854
rect 3887 747 3979 760
<< pdiff >>
rect 2919 1790 3011 1803
rect 2919 1536 2932 1790
rect 2982 1536 3011 1790
rect 2919 1523 3011 1536
rect 3067 1790 3175 1803
rect 3067 1536 3096 1790
rect 3146 1536 3175 1790
rect 3067 1523 3175 1536
rect 3231 1790 3339 1803
rect 3231 1536 3260 1790
rect 3310 1536 3339 1790
rect 3231 1523 3339 1536
rect 3395 1790 3503 1803
rect 3395 1536 3424 1790
rect 3474 1536 3503 1790
rect 3395 1523 3503 1536
rect 3559 1790 3667 1803
rect 3559 1536 3588 1790
rect 3638 1536 3667 1790
rect 3559 1523 3667 1536
rect 3723 1790 3831 1803
rect 3723 1536 3752 1790
rect 3802 1536 3831 1790
rect 3723 1523 3831 1536
rect 3887 1790 3979 1803
rect 3887 1536 3916 1790
rect 3966 1536 3979 1790
rect 3887 1523 3979 1536
<< mvndiff >>
rect -180 1050 -92 1063
rect -180 1004 -167 1050
rect -121 1004 -92 1050
rect -180 946 -92 1004
rect -180 900 -167 946
rect -121 900 -92 946
rect -180 842 -92 900
rect -180 796 -167 842
rect -121 796 -92 842
rect -180 738 -92 796
rect -180 692 -167 738
rect -121 692 -92 738
rect -180 634 -92 692
rect -180 588 -167 634
rect -121 588 -92 634
rect -180 530 -92 588
rect -180 484 -167 530
rect -121 484 -92 530
rect -180 426 -92 484
rect -180 380 -167 426
rect -121 380 -92 426
rect -180 322 -92 380
rect -180 276 -167 322
rect -121 276 -92 322
rect -180 263 -92 276
rect 48 1050 152 1063
rect 48 1004 77 1050
rect 123 1004 152 1050
rect 48 946 152 1004
rect 48 900 77 946
rect 123 900 152 946
rect 48 842 152 900
rect 48 796 77 842
rect 123 796 152 842
rect 48 738 152 796
rect 48 692 77 738
rect 123 692 152 738
rect 48 634 152 692
rect 48 588 77 634
rect 123 588 152 634
rect 48 530 152 588
rect 48 484 77 530
rect 123 484 152 530
rect 48 426 152 484
rect 48 380 77 426
rect 123 380 152 426
rect 48 322 152 380
rect 48 276 77 322
rect 123 276 152 322
rect 48 263 152 276
rect 292 1050 380 1063
rect 292 1004 321 1050
rect 367 1004 380 1050
rect 292 946 380 1004
rect 292 900 321 946
rect 367 900 380 946
rect 292 842 380 900
rect 292 796 321 842
rect 367 796 380 842
rect 292 738 380 796
rect 292 692 321 738
rect 367 692 380 738
rect 292 634 380 692
rect 292 588 321 634
rect 367 588 380 634
rect 292 530 380 588
rect 292 484 321 530
rect 367 484 380 530
rect 292 426 380 484
rect 292 380 321 426
rect 367 380 380 426
rect 292 322 380 380
rect 292 276 321 322
rect 367 276 380 322
rect 292 263 380 276
rect 1167 507 1255 520
rect 1167 461 1180 507
rect 1226 461 1255 507
rect 1167 329 1255 461
rect 1167 283 1180 329
rect 1226 283 1255 329
rect 1167 270 1255 283
rect 1395 507 1499 520
rect 1395 461 1424 507
rect 1470 461 1499 507
rect 1395 329 1499 461
rect 1395 283 1424 329
rect 1470 283 1499 329
rect 1395 270 1499 283
rect 1639 507 1727 520
rect 1639 461 1668 507
rect 1714 461 1727 507
rect 1639 329 1727 461
rect 1639 283 1668 329
rect 1714 283 1727 329
rect 1639 270 1727 283
<< mvpdiff >>
rect 64 2198 152 2211
rect 64 2152 77 2198
rect 123 2152 152 2198
rect 64 2089 152 2152
rect 64 2043 77 2089
rect 123 2043 152 2089
rect 64 1980 152 2043
rect 64 1934 77 1980
rect 123 1934 152 1980
rect 64 1870 152 1934
rect 64 1824 77 1870
rect 123 1824 152 1870
rect 64 1811 152 1824
rect 292 2198 380 2211
rect 292 2152 321 2198
rect 367 2152 380 2198
rect 292 2089 380 2152
rect 292 2043 321 2089
rect 367 2043 380 2089
rect 292 1980 380 2043
rect 292 1934 321 1980
rect 367 1934 380 1980
rect 292 1870 380 1934
rect 292 1824 321 1870
rect 367 1824 380 1870
rect 292 1811 380 1824
rect 923 2009 1011 2022
rect 923 1963 936 2009
rect 982 1963 1011 2009
rect 923 1902 1011 1963
rect 923 1856 936 1902
rect 982 1856 1011 1902
rect 923 1795 1011 1856
rect 923 1749 936 1795
rect 982 1749 1011 1795
rect 923 1688 1011 1749
rect 923 1642 936 1688
rect 982 1642 1011 1688
rect 923 1581 1011 1642
rect 923 1535 936 1581
rect 982 1535 1011 1581
rect 923 1522 1011 1535
rect 1151 2009 1255 2022
rect 1151 1963 1180 2009
rect 1226 1963 1255 2009
rect 1151 1902 1255 1963
rect 1151 1856 1180 1902
rect 1226 1856 1255 1902
rect 1151 1795 1255 1856
rect 1151 1749 1180 1795
rect 1226 1749 1255 1795
rect 1151 1688 1255 1749
rect 1151 1642 1180 1688
rect 1226 1642 1255 1688
rect 1151 1581 1255 1642
rect 1151 1535 1180 1581
rect 1226 1535 1255 1581
rect 1151 1522 1255 1535
rect 1395 2009 1499 2022
rect 1395 1963 1424 2009
rect 1470 1963 1499 2009
rect 1395 1902 1499 1963
rect 1395 1856 1424 1902
rect 1470 1856 1499 1902
rect 1395 1795 1499 1856
rect 1395 1749 1424 1795
rect 1470 1749 1499 1795
rect 1395 1688 1499 1749
rect 1395 1642 1424 1688
rect 1470 1642 1499 1688
rect 1395 1581 1499 1642
rect 1395 1535 1424 1581
rect 1470 1535 1499 1581
rect 1395 1522 1499 1535
rect 1639 2009 1743 2022
rect 1639 1963 1668 2009
rect 1714 1963 1743 2009
rect 1639 1902 1743 1963
rect 1639 1856 1668 1902
rect 1714 1856 1743 1902
rect 1639 1795 1743 1856
rect 1639 1749 1668 1795
rect 1714 1749 1743 1795
rect 1639 1688 1743 1749
rect 1639 1642 1668 1688
rect 1714 1642 1743 1688
rect 1639 1581 1743 1642
rect 1639 1535 1668 1581
rect 1714 1535 1743 1581
rect 1639 1522 1743 1535
rect 1883 2009 1971 2022
rect 1883 1963 1912 2009
rect 1958 1963 1971 2009
rect 1883 1902 1971 1963
rect 1883 1856 1912 1902
rect 1958 1856 1971 1902
rect 1883 1795 1971 1856
rect 1883 1749 1912 1795
rect 1958 1749 1971 1795
rect 1883 1688 1971 1749
rect 1883 1642 1912 1688
rect 1958 1642 1971 1688
rect 1883 1581 1971 1642
rect 1883 1535 1912 1581
rect 1958 1535 1971 1581
rect 1883 1522 1971 1535
<< ndiffc >>
rect 2932 760 2982 854
rect 3096 760 3146 854
rect 3260 760 3310 854
rect 3424 760 3474 854
rect 3588 760 3638 854
rect 3752 760 3802 854
rect 3916 760 3966 854
<< pdiffc >>
rect 2932 1536 2982 1790
rect 3096 1536 3146 1790
rect 3260 1536 3310 1790
rect 3424 1536 3474 1790
rect 3588 1536 3638 1790
rect 3752 1536 3802 1790
rect 3916 1536 3966 1790
<< mvndiffc >>
rect -167 1004 -121 1050
rect -167 900 -121 946
rect -167 796 -121 842
rect -167 692 -121 738
rect -167 588 -121 634
rect -167 484 -121 530
rect -167 380 -121 426
rect -167 276 -121 322
rect 77 1004 123 1050
rect 77 900 123 946
rect 77 796 123 842
rect 77 692 123 738
rect 77 588 123 634
rect 77 484 123 530
rect 77 380 123 426
rect 77 276 123 322
rect 321 1004 367 1050
rect 321 900 367 946
rect 321 796 367 842
rect 321 692 367 738
rect 321 588 367 634
rect 321 484 367 530
rect 321 380 367 426
rect 321 276 367 322
rect 1180 461 1226 507
rect 1180 283 1226 329
rect 1424 461 1470 507
rect 1424 283 1470 329
rect 1668 461 1714 507
rect 1668 283 1714 329
<< mvpdiffc >>
rect 77 2152 123 2198
rect 77 2043 123 2089
rect 77 1934 123 1980
rect 77 1824 123 1870
rect 321 2152 367 2198
rect 321 2043 367 2089
rect 321 1934 367 1980
rect 321 1824 367 1870
rect 936 1963 982 2009
rect 936 1856 982 1902
rect 936 1749 982 1795
rect 936 1642 982 1688
rect 936 1535 982 1581
rect 1180 1963 1226 2009
rect 1180 1856 1226 1902
rect 1180 1749 1226 1795
rect 1180 1642 1226 1688
rect 1180 1535 1226 1581
rect 1424 1963 1470 2009
rect 1424 1856 1470 1902
rect 1424 1749 1470 1795
rect 1424 1642 1470 1688
rect 1424 1535 1470 1581
rect 1668 1963 1714 2009
rect 1668 1856 1714 1902
rect 1668 1749 1714 1795
rect 1668 1642 1714 1688
rect 1668 1535 1714 1581
rect 1912 1963 1958 2009
rect 1912 1856 1958 1902
rect 1912 1749 1958 1795
rect 1912 1642 1958 1688
rect 1912 1535 1958 1581
<< psubdiff >>
rect -443 1196 -353 1218
rect -443 22 -421 1196
rect -375 90 -353 1196
rect 520 1196 610 1218
rect 520 90 542 1196
rect -375 68 542 90
rect 471 22 542 68
rect 588 22 610 1196
rect -443 0 610 22
rect 716 1008 806 1030
rect 716 22 738 1008
rect 784 90 806 1008
rect 4064 1041 4154 1055
rect 2771 840 2861 854
rect 1998 810 2088 832
rect 1998 90 2020 810
rect 784 68 2020 90
rect 784 22 892 68
rect 1962 22 2020 68
rect 2066 22 2088 810
rect 2771 602 2793 840
rect 2839 670 2861 840
rect 4064 670 4086 1041
rect 2839 648 4086 670
rect 2839 602 2887 648
rect 4032 602 4086 648
rect 4132 602 4154 1041
rect 2771 580 4154 602
rect 716 0 2088 22
<< nsubdiff >>
rect -164 2470 610 2492
rect -164 1766 -142 2470
rect -96 2424 12 2470
rect 434 2424 542 2470
rect -96 2402 542 2424
rect -96 1766 -74 2402
rect -164 1744 -74 1766
rect 520 1766 542 2402
rect 588 1766 610 2470
rect 520 1744 610 1766
rect 716 2470 2178 2492
rect 716 1484 738 2470
rect 784 2424 860 2470
rect 1970 2424 2110 2470
rect 784 2402 2110 2424
rect 784 1484 806 2402
rect 716 1462 806 1484
rect 2088 1519 2110 2402
rect 2156 1519 2178 2470
rect 2765 1950 4160 1972
rect 2765 1544 2787 1950
rect 2833 1904 2894 1950
rect 4041 1904 4092 1950
rect 2833 1882 4092 1904
rect 2833 1544 2855 1882
rect 2765 1522 2855 1544
rect 2088 1497 2178 1519
rect 4070 1484 4092 1882
rect 4138 1484 4160 1950
rect 4070 1462 4160 1484
<< psubdiffcont >>
rect -421 68 -375 1196
rect -421 22 471 68
rect 542 22 588 1196
rect 738 22 784 1008
rect 892 22 1962 68
rect 2020 22 2066 810
rect 2793 602 2839 840
rect 2887 602 4032 648
rect 4086 602 4132 1041
<< nsubdiffcont >>
rect -142 1766 -96 2470
rect 12 2424 434 2470
rect 542 1766 588 2470
rect 738 1484 784 2470
rect 860 2424 1970 2470
rect 2110 1519 2156 2470
rect 2787 1544 2833 1950
rect 2894 1904 4041 1950
rect 4092 1484 4138 1950
<< polysilicon >>
rect 152 2211 292 2255
rect -92 1412 48 1431
rect -92 1272 -47 1412
rect -1 1272 48 1412
rect -92 1063 48 1272
rect 152 1412 292 1811
rect 1011 2022 1151 2066
rect 1255 2022 1395 2066
rect 1499 2022 1639 2066
rect 1743 2022 1883 2066
rect 152 1272 199 1412
rect 245 1272 292 1412
rect 152 1063 292 1272
rect 1011 1265 1151 1522
rect -92 219 48 263
rect 152 219 292 263
rect 1011 1125 1058 1265
rect 1104 1125 1151 1265
rect 1011 1106 1151 1125
rect 1255 1265 1395 1522
rect 1255 1125 1302 1265
rect 1348 1125 1395 1265
rect 1255 520 1395 1125
rect 1499 1265 1639 1522
rect 1499 1125 1546 1265
rect 1592 1125 1639 1265
rect 1499 520 1639 1125
rect 1743 1265 1883 1522
rect 3011 1803 3067 1857
rect 3175 1803 3231 1857
rect 3339 1803 3395 1857
rect 3503 1803 3559 1857
rect 3667 1803 3723 1857
rect 3831 1803 3887 1857
rect 3011 1279 3067 1523
rect 3175 1279 3231 1523
rect 3339 1279 3395 1523
rect 3503 1279 3559 1523
rect 3667 1279 3723 1523
rect 3831 1279 3887 1523
rect 1743 1125 1790 1265
rect 1836 1125 1883 1265
rect 1743 1106 1883 1125
rect 3001 1265 3075 1279
rect 3001 1125 3016 1265
rect 3062 1125 3075 1265
rect 3001 1111 3075 1125
rect 3165 1265 3241 1279
rect 3165 1125 3180 1265
rect 3226 1125 3241 1265
rect 3165 1111 3241 1125
rect 3329 1265 3403 1279
rect 3329 1125 3344 1265
rect 3390 1125 3403 1265
rect 3329 1111 3403 1125
rect 3493 1265 3567 1279
rect 3493 1125 3508 1265
rect 3554 1125 3567 1265
rect 3493 1111 3567 1125
rect 3657 1265 3733 1279
rect 3657 1125 3672 1265
rect 3718 1125 3733 1265
rect 3657 1111 3733 1125
rect 3821 1265 3897 1279
rect 3821 1125 3836 1265
rect 3882 1125 3897 1265
rect 3821 1111 3897 1125
rect 3011 867 3067 1111
rect 3175 867 3231 1111
rect 3339 867 3395 1111
rect 3503 867 3559 1111
rect 3667 867 3723 1111
rect 3831 867 3887 1111
rect 1255 226 1395 270
rect 1499 226 1639 270
rect 3011 700 3067 747
rect 3175 700 3231 747
rect 3339 700 3395 747
rect 3503 700 3559 747
rect 3667 700 3723 747
rect 3831 700 3887 747
<< polycontact >>
rect -47 1272 -1 1412
rect 199 1272 245 1412
rect 1058 1125 1104 1265
rect 1302 1125 1348 1265
rect 1546 1125 1592 1265
rect 1790 1125 1836 1265
rect 3016 1125 3062 1265
rect 3180 1125 3226 1265
rect 3344 1125 3390 1265
rect 3508 1125 3554 1265
rect 3672 1125 3718 1265
rect 3836 1125 3882 1265
<< metal1 >>
rect -153 2470 599 2481
rect -153 1766 -142 2470
rect -96 2424 12 2470
rect 434 2424 542 2470
rect -96 2413 542 2424
rect -96 1766 -85 2413
rect 62 2198 138 2413
rect 62 2152 77 2198
rect 123 2152 138 2198
rect 62 2089 138 2152
rect 62 2043 77 2089
rect 123 2043 138 2089
rect 62 1980 138 2043
rect 62 1934 77 1980
rect 123 1934 138 1980
rect 62 1870 138 1934
rect 62 1824 77 1870
rect 123 1824 138 1870
rect 62 1811 138 1824
rect 306 2198 382 2211
rect 306 2152 321 2198
rect 367 2152 382 2198
rect 306 2089 382 2152
rect 306 2043 321 2089
rect 367 2043 382 2089
rect 306 1980 382 2043
rect 306 1934 321 1980
rect 367 1934 382 1980
rect 306 1870 382 1934
rect 306 1824 321 1870
rect 367 1824 382 1870
rect -153 1755 -85 1766
rect -58 1412 10 1423
rect -58 1272 -47 1412
rect -1 1272 10 1412
rect -58 1261 10 1272
rect 188 1412 256 1423
rect 188 1272 199 1412
rect 245 1272 256 1412
rect 188 1261 256 1272
rect 306 1391 382 1824
rect 531 1766 542 2413
rect 588 1766 599 2470
rect 531 1755 599 1766
rect 727 2470 2167 2481
rect 727 1484 738 2470
rect 784 2424 860 2470
rect 1970 2424 2110 2470
rect 784 2413 2110 2424
rect 784 1484 795 2413
rect 921 2177 1973 2321
rect 921 2009 997 2177
rect 921 1963 936 2009
rect 982 1963 997 2009
rect 921 1902 997 1963
rect 1180 2009 1226 2022
rect 1180 1958 1226 1963
rect 1409 2009 1485 2177
rect 1409 1963 1424 2009
rect 1470 1963 1485 2009
rect 921 1856 936 1902
rect 982 1856 997 1902
rect 921 1795 997 1856
rect 921 1749 936 1795
rect 982 1749 997 1795
rect 921 1688 997 1749
rect 921 1642 936 1688
rect 982 1642 997 1688
rect 921 1581 997 1642
rect 921 1535 936 1581
rect 982 1535 997 1581
rect 921 1522 997 1535
rect 1165 1902 1241 1958
rect 1165 1856 1180 1902
rect 1226 1856 1241 1902
rect 1165 1795 1241 1856
rect 1165 1749 1180 1795
rect 1226 1749 1241 1795
rect 1165 1688 1241 1749
rect 1165 1642 1180 1688
rect 1226 1642 1241 1688
rect 1165 1581 1241 1642
rect 1165 1535 1180 1581
rect 1226 1535 1241 1581
rect 727 1473 795 1484
rect 1165 1442 1241 1535
rect 1409 1902 1485 1963
rect 1668 2009 1714 2022
rect 1668 1958 1714 1963
rect 1897 2009 1973 2177
rect 1897 1963 1912 2009
rect 1958 1963 1973 2009
rect 1409 1856 1424 1902
rect 1470 1856 1485 1902
rect 1409 1795 1485 1856
rect 1409 1749 1424 1795
rect 1470 1749 1485 1795
rect 1409 1688 1485 1749
rect 1409 1642 1424 1688
rect 1470 1642 1485 1688
rect 1409 1581 1485 1642
rect 1409 1535 1424 1581
rect 1470 1535 1485 1581
rect 1409 1522 1485 1535
rect 1653 1902 1729 1958
rect 1653 1856 1668 1902
rect 1714 1856 1729 1902
rect 1653 1795 1729 1856
rect 1653 1749 1668 1795
rect 1714 1749 1729 1795
rect 1653 1688 1729 1749
rect 1653 1642 1668 1688
rect 1714 1642 1729 1688
rect 1653 1581 1729 1642
rect 1653 1535 1668 1581
rect 1714 1535 1729 1581
rect 1653 1442 1729 1535
rect 1897 1902 1973 1963
rect 1897 1856 1912 1902
rect 1958 1856 1973 1902
rect 1897 1795 1973 1856
rect 1897 1749 1912 1795
rect 1958 1749 1973 1795
rect 1897 1688 1973 1749
rect 1897 1642 1912 1688
rect 1958 1642 1973 1688
rect 1897 1581 1973 1642
rect 1897 1535 1912 1581
rect 1958 1535 1973 1581
rect 1897 1522 1973 1535
rect 2099 1519 2110 2413
rect 2156 1519 2167 2470
rect 2776 1950 4149 1961
rect 2776 1544 2787 1950
rect 2833 1904 2894 1950
rect 4041 1904 4092 1950
rect 2833 1893 4092 1904
rect 2833 1544 2844 1893
rect 2776 1533 2844 1544
rect 2919 1790 2995 1893
rect 2919 1536 2932 1790
rect 2982 1536 2995 1790
rect 2919 1523 2995 1536
rect 3083 1790 3159 1803
rect 3083 1536 3096 1790
rect 3146 1536 3159 1790
rect 2099 1503 2167 1519
rect 3083 1445 3159 1536
rect 3247 1790 3323 1893
rect 3247 1536 3260 1790
rect 3310 1536 3323 1790
rect 3247 1523 3323 1536
rect 3411 1790 3487 1803
rect 3411 1536 3424 1790
rect 3474 1536 3487 1790
rect 3084 1442 3159 1445
rect 3411 1442 3487 1536
rect 3575 1790 3651 1893
rect 3575 1536 3588 1790
rect 3638 1536 3651 1790
rect 3575 1523 3651 1536
rect 3739 1790 3815 1803
rect 3739 1536 3752 1790
rect 3802 1536 3815 1790
rect 3739 1442 3815 1536
rect 3903 1790 3979 1893
rect 3903 1536 3916 1790
rect 3966 1536 3979 1790
rect 3903 1523 3979 1536
rect 4081 1484 4092 1893
rect 4138 1484 4149 1950
rect 4081 1473 4149 1484
rect 306 1291 917 1391
rect 1165 1366 2073 1442
rect 3084 1366 4028 1442
rect -432 1196 -364 1207
rect -432 22 -421 1196
rect -375 79 -364 1196
rect -167 1050 -121 1063
rect -167 946 -121 1004
rect 77 1050 123 1063
rect 77 990 123 1004
rect 306 1050 382 1291
rect 817 1276 917 1291
rect 1997 1276 2073 1366
rect 817 1265 1847 1276
rect 306 1004 321 1050
rect 367 1004 382 1050
rect -167 842 -121 900
rect -167 738 -121 796
rect -182 696 -167 708
rect 62 946 138 990
rect 62 900 77 946
rect 123 900 138 946
rect 62 842 138 900
rect 62 796 77 842
rect 123 796 138 842
rect 62 738 138 796
rect -121 696 -106 708
rect -182 332 -170 696
rect -118 332 -106 696
rect -182 322 -106 332
rect -182 320 -167 322
rect -121 320 -106 322
rect 62 692 77 738
rect 123 692 138 738
rect 62 634 138 692
rect 62 588 77 634
rect 123 588 138 634
rect 62 530 138 588
rect 62 484 77 530
rect 123 484 138 530
rect 62 426 138 484
rect 62 380 77 426
rect 123 380 138 426
rect 62 322 138 380
rect -167 263 -121 276
rect 62 276 77 322
rect 123 276 138 322
rect 62 79 138 276
rect 306 946 382 1004
rect 306 900 321 946
rect 367 900 382 946
rect 306 842 382 900
rect 306 796 321 842
rect 367 796 382 842
rect 306 738 382 796
rect 306 696 321 738
rect 367 696 382 738
rect 306 332 318 696
rect 370 332 382 696
rect 306 322 382 332
rect 306 276 321 322
rect 367 276 382 322
rect 306 263 382 276
rect 531 1196 599 1207
rect 531 79 542 1196
rect -375 68 542 79
rect 471 22 542 68
rect 588 22 599 1196
rect 817 1125 1058 1265
rect 1104 1125 1302 1265
rect 1348 1125 1546 1265
rect 1592 1125 1790 1265
rect 1836 1125 1847 1265
rect 817 1114 1847 1125
rect 1997 1265 3893 1276
rect 1997 1125 3016 1265
rect 3062 1125 3180 1265
rect 3226 1125 3344 1265
rect 3390 1125 3508 1265
rect 3554 1125 3672 1265
rect 3718 1125 3836 1265
rect 3882 1125 3893 1265
rect 1997 1114 3893 1125
rect 1997 1019 2073 1114
rect 3952 1019 4028 1366
rect -432 11 599 22
rect 727 1008 795 1019
rect 727 22 738 1008
rect 784 79 795 1008
rect 1409 943 2073 1019
rect 3083 943 4028 1019
rect 4075 1041 4143 1053
rect 1165 507 1241 520
rect 1165 461 1180 507
rect 1226 461 1241 507
rect 1165 329 1241 461
rect 1165 283 1180 329
rect 1226 283 1241 329
rect 1165 204 1241 283
rect 1409 507 1485 943
rect 2919 854 2995 867
rect 2782 840 2850 852
rect 2009 810 2077 821
rect 1409 461 1424 507
rect 1470 461 1485 507
rect 1409 329 1485 461
rect 1409 283 1424 329
rect 1470 283 1485 329
rect 1409 270 1485 283
rect 1653 507 1729 520
rect 1653 461 1668 507
rect 1714 461 1729 507
rect 1653 329 1729 461
rect 1653 283 1668 329
rect 1714 283 1729 329
rect 1653 204 1729 283
rect 1165 134 1729 204
rect 2009 79 2020 810
rect 784 68 2020 79
rect 784 22 892 68
rect 1962 22 2020 68
rect 2066 22 2077 810
rect 2782 602 2793 840
rect 2839 659 2850 840
rect 2919 760 2932 854
rect 2982 760 2995 854
rect 2919 659 2995 760
rect 3083 854 3159 943
rect 3083 760 3096 854
rect 3146 760 3159 854
rect 3083 748 3159 760
rect 3247 854 3323 867
rect 3247 760 3260 854
rect 3310 760 3323 854
rect 3247 659 3323 760
rect 3411 854 3487 943
rect 3411 760 3424 854
rect 3474 760 3487 854
rect 3411 748 3487 760
rect 3575 854 3651 867
rect 3575 760 3588 854
rect 3638 760 3651 854
rect 3575 659 3651 760
rect 3739 854 3815 943
rect 3739 760 3752 854
rect 3802 760 3815 854
rect 3739 748 3815 760
rect 3901 854 3977 867
rect 3901 760 3916 854
rect 3966 760 3977 854
rect 3901 659 3977 760
rect 4075 659 4086 1041
rect 2839 648 4086 659
rect 2839 602 2887 648
rect 4032 602 4086 648
rect 4132 602 4143 1041
rect 2782 591 4143 602
rect 727 11 2077 22
<< via1 >>
rect -170 692 -167 696
rect -167 692 -121 696
rect -121 692 -118 696
rect -170 634 -118 692
rect -170 588 -167 634
rect -167 588 -121 634
rect -121 588 -118 634
rect -170 530 -118 588
rect -170 484 -167 530
rect -167 484 -121 530
rect -121 484 -118 530
rect -170 426 -118 484
rect -170 380 -167 426
rect -167 380 -121 426
rect -121 380 -118 426
rect -170 332 -118 380
rect 318 692 321 696
rect 321 692 367 696
rect 367 692 370 696
rect 318 634 370 692
rect 318 588 321 634
rect 321 588 367 634
rect 367 588 370 634
rect 318 530 370 588
rect 318 484 321 530
rect 321 484 367 530
rect 367 484 370 530
rect 318 426 370 484
rect 318 380 321 426
rect 321 380 367 426
rect 367 380 370 426
rect 318 332 370 380
<< metal2 >>
rect -182 696 -106 708
rect -182 332 -170 696
rect -118 573 -106 696
rect 306 696 382 708
rect 306 573 318 696
rect -118 435 318 573
rect -118 332 -106 435
rect -182 320 -106 332
rect 306 332 318 435
rect 370 332 382 696
rect 306 320 382 332
<< labels >>
rlabel metal1 s 2 2452 2 2452 4 DVDD
port 1 nsew
rlabel metal1 s 225 1326 225 1326 4 A
port 2 nsew
rlabel metal1 s 80 45 80 45 4 DVSS
port 3 nsew
rlabel metal1 s -21 1326 -21 1326 4 A
port 2 nsew
rlabel metal1 s 1452 2452 1452 2452 4 VDD
port 4 nsew
rlabel metal1 s 1082 45 1082 45 4 VSS
port 5 nsew
rlabel metal1 s 3642 1200 3642 1200 4 Z
port 6 nsew
<< end >>
