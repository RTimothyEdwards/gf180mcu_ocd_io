* NGSPICE file created from gf180mcu_ocd_io__fill5.ext - technology: gf180mcuD

.subckt POLY_SUB_FILL a_1165_n91# a_1077_1#
X0 a_1165_n91# a_1077_1# cap_nmos_06v0 c_width=1.5u c_length=1.5u
X1 a_1165_n91# a_1077_1# cap_nmos_06v0 c_width=1.5u c_length=1.5u
.ends

.subckt GF_NI_FILL5_1 VSS VDD DVSS DVDD
XPOLY_SUB_FILL_0[0] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[1] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[2] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[3] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[4] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[5] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[6] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[7] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[8] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[9] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[10] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[11] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[12] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[13] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[14] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[15] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[16] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[17] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[18] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[19] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[20] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[21] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[22] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[23] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[24] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[25] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[26] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[27] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[28] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[29] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[30] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[31] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[32] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[33] VDD VSS POLY_SUB_FILL
XPOLY_SUB_FILL_0[34] VDD VSS POLY_SUB_FILL
.ends

.subckt GF_NI_FILL5_0 DVSS DVDD VDD VSS
XGF_NI_FILL5_1_0 VSS VDD DVSS DVDD GF_NI_FILL5_1
.ends

.subckt gf180mcu_ocd_io__fill5 DVDD DVSS VDD VSS
XGF_NI_FILL5_0_0 DVSS DVDD VDD VSS GF_NI_FILL5_0
.ends

