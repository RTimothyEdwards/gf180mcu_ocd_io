VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_ocd_io__vdd
  CLASS PAD POWER ;
  FOREIGN gf180mcu_ocd_io__vdd ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 350.000 ;
  SYMMETRY X Y R90 ;
  SITE GF_IO_Site ;
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 334.000 75.000 341.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 294.000 75.000 301.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 278.000 75.000 285.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 270.000 75.000 277.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 262.000 75.000 269.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 206.000 75.000 213.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 214.000 75.000 229.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 182.000 75.000 197.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 166.000 75.000 181.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 150.000 75.000 165.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 134.000 75.000 149.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 118.000 75.000 125.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 86.000 75.000 101.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 70.000 75.000 85.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 230.000 75.000 245.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 198.000 75.000 205.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 126.000 75.000 133.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 102.000 75.000 117.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 286.000 75.000 293.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 302.000 75.000 309.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 326.000 75.000 333.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 342.000 75.000 348.390 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal2 ;
        RECT 1.360 345.345 10.860 350.000 ;
    END
    PORT
      LAYER Metal2 ;
        RECT 13.760 345.345 24.010 350.000 ;
    END
    PORT
      LAYER Metal2 ;
        RECT 25.610 345.345 35.860 350.000 ;
    END
    PORT
      LAYER Metal2 ;
        RECT 39.140 345.345 49.390 350.000 ;
    END
    PORT
      LAYER Metal2 ;
        RECT 50.990 345.345 61.240 350.000 ;
    END
    PORT
      LAYER Metal2 ;
        RECT 64.140 345.345 73.640 350.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 7.500 2.000 67.500 62.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 310.000 5.000 317.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 254.000 5.000 261.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 70.000 310.000 75.000 317.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 70.000 254.000 75.000 261.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 246.000 5.000 253.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 318.000 5.000 325.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 70.000 246.000 75.000 253.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 70.000 318.000 75.000 325.000 ;
    END
  END VSS
  OBS
      LAYER Nwell ;
        RECT 3.060 67.480 71.940 345.275 ;
      LAYER Metal1 ;
        RECT -0.160 65.540 75.160 349.785 ;
      LAYER Metal2 ;
        RECT 0.000 345.045 1.060 348.390 ;
        RECT 11.160 345.045 13.460 348.390 ;
        RECT 24.310 345.045 25.310 348.390 ;
        RECT 36.160 345.045 38.840 348.390 ;
        RECT 49.690 345.045 50.690 348.390 ;
        RECT 61.540 345.045 63.840 348.390 ;
        RECT 73.940 345.045 75.000 348.390 ;
        RECT 0.000 0.000 75.000 345.045 ;
      LAYER Metal3 ;
        RECT 6.800 310.800 68.200 324.200 ;
        RECT 6.800 246.800 68.200 260.200 ;
        RECT 3.500 63.800 71.500 68.200 ;
        RECT 3.500 0.200 5.700 63.800 ;
        RECT 69.300 0.200 71.500 63.800 ;
        RECT 3.500 0.000 71.500 0.200 ;
  END
END gf180mcu_ocd_io__vdd
END LIBRARY

