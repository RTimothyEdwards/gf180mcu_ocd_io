magic
tech gf180mcuD
magscale 1 10
timestamp 1758724778
<< nwell >>
rect 16038 51147 16457 51634
<< nmos >>
rect 16224 50941 16280 51061
<< pmos >>
rect 16224 51233 16280 51473
<< ndiff >>
rect 16135 51048 16224 51061
rect 16135 50956 16149 51048
rect 16195 50956 16224 51048
rect 16135 50941 16224 50956
rect 16280 51047 16368 51061
rect 16280 50955 16309 51047
rect 16355 50955 16368 51047
rect 16280 50941 16368 50955
<< pdiff >>
rect 16131 51459 16224 51473
rect 16131 51246 16144 51459
rect 16190 51246 16224 51459
rect 16131 51233 16224 51246
rect 16280 51459 16368 51473
rect 16280 51246 16309 51459
rect 16355 51246 16368 51459
rect 16280 51233 16368 51246
<< ndiffc >>
rect 16149 50956 16195 51048
rect 16309 50955 16355 51047
<< pdiffc >>
rect 16144 51246 16190 51459
rect 16309 51246 16355 51459
<< psubdiff >>
rect 16066 50872 16182 50885
rect 16360 50872 16432 50885
rect 16066 50826 16079 50872
rect 16125 50826 16373 50872
rect 16419 50826 16432 50872
rect 16066 50813 16432 50826
<< nsubdiff >>
rect 16066 51588 16432 51601
rect 16066 51542 16079 51588
rect 16125 51547 16373 51588
rect 16125 51542 16184 51547
rect 16066 51529 16184 51542
rect 16359 51542 16373 51547
rect 16419 51542 16432 51588
rect 16359 51529 16432 51542
<< psubdiffcont >>
rect 16079 50826 16125 50872
rect 16373 50826 16419 50872
<< nsubdiffcont >>
rect 16079 51542 16125 51588
rect 16373 51542 16419 51588
<< polysilicon >>
rect 16224 51473 16280 51520
rect 16224 51178 16280 51233
rect 16119 51165 16280 51178
rect 16119 51119 16132 51165
rect 16252 51119 16280 51165
rect 16119 51106 16280 51119
rect 16224 51061 16280 51106
rect 16224 50897 16280 50941
<< polycontact >>
rect 16132 51119 16252 51165
<< metal1 >>
rect 16066 51588 16432 51601
rect 16066 51542 16079 51588
rect 16125 51542 16373 51588
rect 16419 51542 16432 51588
rect 16066 51526 16432 51542
rect 16144 51459 16190 51526
rect 16144 51235 16190 51246
rect 16309 51459 16355 51470
rect 16121 51119 16132 51165
rect 16252 51119 16263 51165
rect 16149 51048 16195 51059
rect 16149 50889 16195 50956
rect 16309 51047 16355 51246
rect 16309 50944 16355 50955
rect 16066 50872 16432 50889
rect 16066 50826 16079 50872
rect 16125 50826 16373 50872
rect 16419 50826 16432 50872
rect 16066 50813 16432 50826
<< end >>
