magic
tech gf180mcuD
magscale 1 10
timestamp 1758724778
<< nwell >>
rect 16932 51136 17513 51623
<< nmos >>
rect 17148 50930 17204 51050
rect 17280 50930 17336 51050
<< pmos >>
rect 17113 51222 17169 51462
rect 17280 51222 17336 51462
<< ndiff >>
rect 17059 51037 17148 51050
rect 17059 50945 17073 51037
rect 17119 50945 17148 51037
rect 17059 50930 17148 50945
rect 17204 50930 17280 51050
rect 17336 51036 17424 51050
rect 17336 50944 17365 51036
rect 17411 50944 17424 51036
rect 17336 50930 17424 50944
<< pdiff >>
rect 17024 51449 17113 51462
rect 17024 51236 17038 51449
rect 17084 51236 17113 51449
rect 17024 51222 17113 51236
rect 17169 51448 17280 51462
rect 17169 51315 17200 51448
rect 17246 51315 17280 51448
rect 17169 51222 17280 51315
rect 17336 51448 17424 51462
rect 17336 51235 17365 51448
rect 17411 51235 17424 51448
rect 17336 51222 17424 51235
<< ndiffc >>
rect 17073 50945 17119 51037
rect 17365 50944 17411 51036
<< pdiffc >>
rect 17038 51236 17084 51449
rect 17200 51315 17246 51448
rect 17365 51235 17411 51448
<< psubdiff >>
rect 16960 50861 17033 50874
rect 17375 50861 17488 50874
rect 16960 50815 16973 50861
rect 17019 50815 17429 50861
rect 17475 50815 17488 50861
rect 16960 50802 17488 50815
<< nsubdiff >>
rect 16956 51577 17488 51590
rect 16956 51531 16973 51577
rect 17019 51536 17429 51577
rect 17019 51531 17035 51536
rect 16956 51518 17035 51531
rect 17374 51531 17429 51536
rect 17475 51531 17488 51577
rect 17374 51518 17488 51531
<< psubdiffcont >>
rect 16973 50815 17019 50861
rect 17429 50815 17475 50861
<< nsubdiffcont >>
rect 16973 51531 17019 51577
rect 17429 51531 17475 51577
<< polysilicon >>
rect 17113 51462 17169 51506
rect 17280 51462 17336 51506
rect 17113 51168 17169 51222
rect 17113 51154 17204 51168
rect 17280 51167 17336 51222
rect 17113 51108 17132 51154
rect 17182 51108 17204 51154
rect 17113 51095 17204 51108
rect 17252 51154 17336 51167
rect 17252 51108 17268 51154
rect 17318 51108 17336 51154
rect 17252 51095 17336 51108
rect 17148 51050 17204 51095
rect 17280 51050 17336 51095
rect 17148 50885 17204 50930
rect 17280 50886 17336 50930
<< polycontact >>
rect 17132 51108 17182 51154
rect 17268 51108 17318 51154
<< metal1 >>
rect 16956 51577 17488 51590
rect 16956 51531 16973 51577
rect 17019 51531 17429 51577
rect 17475 51531 17488 51577
rect 16956 51515 17488 51531
rect 17038 51449 17084 51461
rect 17179 51448 17270 51515
rect 17179 51315 17200 51448
rect 17246 51315 17270 51448
rect 17179 51304 17270 51315
rect 17365 51448 17411 51459
rect 17084 51236 17365 51258
rect 17038 51235 17365 51236
rect 17038 51211 17411 51235
rect 17059 51154 17218 51165
rect 17059 51108 17132 51154
rect 17182 51108 17218 51154
rect 17059 51094 17218 51108
rect 17268 51154 17318 51165
rect 17073 51037 17119 51048
rect 17268 51046 17318 51108
rect 17073 50878 17119 50945
rect 17213 50983 17318 51046
rect 17365 51036 17411 51211
rect 17213 50940 17271 50983
rect 17365 50933 17411 50944
rect 16960 50861 17488 50878
rect 16960 50815 16973 50861
rect 17019 50815 17429 50861
rect 17475 50815 17488 50861
rect 16960 50802 17488 50815
<< end >>
