magic
tech gf180mcuA
magscale 1 10
timestamp 1758828810
<< metal3 >>
rect 0 63600 400 65000
rect 0 49200 400 50600
use GF_NI_BRK2_0  GF_NI_BRK2_0_0 ..
timestamp 1484609607
transform 1 0 0 0 1 0
box -32 13097 432 69968
<< labels >>
flabel metal3 s 0 63600 400 65000 0 FreeSans 1600 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal3 s 0 49200 400 50600 0 FreeSans 1600 90 0 0 VSS
port 1 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 400 70000
string LEFclass PAD SPACER
string LEFsite GF_IO_Site
string LEFsymmetry X Y R90
<< end >>
