magic
tech gf180mcuD
magscale 1 10
timestamp 1758749514
<< isosubstrate >>
rect 13458 69312 69613 70630
rect 13458 56958 70557 69312
rect 13436 56517 70557 56958
rect 13436 44853 52740 56517
tri 13436 13361 44928 44853 ne
rect 44928 41550 52740 44853
rect 44928 13361 56957 41550
<< psubdiff >>
rect 60177 70507 69501 70529
rect 60177 70461 60199 70507
rect 60245 70461 60313 70507
rect 60359 70461 60427 70507
rect 60473 70461 60541 70507
rect 60587 70461 60655 70507
rect 60701 70461 60769 70507
rect 60815 70461 60883 70507
rect 60929 70461 60997 70507
rect 61043 70461 61111 70507
rect 61157 70461 61225 70507
rect 61271 70461 61339 70507
rect 61385 70461 61453 70507
rect 61499 70461 61567 70507
rect 61613 70461 61681 70507
rect 61727 70461 61795 70507
rect 61841 70461 61909 70507
rect 61955 70461 62023 70507
rect 62069 70461 62137 70507
rect 62183 70461 62251 70507
rect 62297 70461 62365 70507
rect 62411 70461 62479 70507
rect 62525 70461 62593 70507
rect 62639 70461 62707 70507
rect 62753 70461 62821 70507
rect 62867 70461 62935 70507
rect 62981 70461 63049 70507
rect 63095 70461 63163 70507
rect 63209 70461 63277 70507
rect 63323 70461 63391 70507
rect 63437 70461 63505 70507
rect 63551 70461 63619 70507
rect 63665 70461 63733 70507
rect 63779 70461 63847 70507
rect 63893 70461 63961 70507
rect 64007 70461 64075 70507
rect 64121 70461 64189 70507
rect 64235 70461 64303 70507
rect 64349 70461 64417 70507
rect 64463 70461 64531 70507
rect 64577 70461 64645 70507
rect 64691 70461 64759 70507
rect 64805 70461 64873 70507
rect 64919 70461 64987 70507
rect 65033 70461 65101 70507
rect 65147 70461 65215 70507
rect 65261 70461 65329 70507
rect 65375 70461 65443 70507
rect 65489 70461 65557 70507
rect 65603 70461 65671 70507
rect 65717 70461 65785 70507
rect 65831 70461 65899 70507
rect 65945 70461 66013 70507
rect 66059 70461 66127 70507
rect 66173 70461 66241 70507
rect 66287 70461 66355 70507
rect 66401 70461 66469 70507
rect 66515 70461 66583 70507
rect 66629 70461 66697 70507
rect 66743 70461 66811 70507
rect 66857 70461 66925 70507
rect 66971 70461 67039 70507
rect 67085 70461 67153 70507
rect 67199 70461 67267 70507
rect 67313 70461 67381 70507
rect 67427 70461 67495 70507
rect 67541 70461 67609 70507
rect 67655 70461 67723 70507
rect 67769 70461 67837 70507
rect 67883 70461 67951 70507
rect 67997 70461 68065 70507
rect 68111 70461 68179 70507
rect 68225 70461 68293 70507
rect 68339 70461 68407 70507
rect 68453 70461 68521 70507
rect 68567 70461 68635 70507
rect 68681 70461 68749 70507
rect 68795 70461 68863 70507
rect 68909 70461 68977 70507
rect 69023 70461 69091 70507
rect 69137 70461 69205 70507
rect 69251 70461 69319 70507
rect 69365 70461 69433 70507
rect 69479 70461 69501 70507
rect 60177 70393 69501 70461
rect 60177 70347 60199 70393
rect 60245 70347 60313 70393
rect 60359 70347 60427 70393
rect 60473 70347 60541 70393
rect 60587 70347 60655 70393
rect 60701 70347 60769 70393
rect 60815 70347 60883 70393
rect 60929 70347 60997 70393
rect 61043 70347 61111 70393
rect 61157 70347 61225 70393
rect 61271 70347 61339 70393
rect 61385 70347 61453 70393
rect 61499 70347 61567 70393
rect 61613 70347 61681 70393
rect 61727 70347 61795 70393
rect 61841 70347 61909 70393
rect 61955 70347 62023 70393
rect 62069 70347 62137 70393
rect 62183 70347 62251 70393
rect 62297 70347 62365 70393
rect 62411 70347 62479 70393
rect 62525 70347 62593 70393
rect 62639 70347 62707 70393
rect 62753 70347 62821 70393
rect 62867 70347 62935 70393
rect 62981 70347 63049 70393
rect 63095 70347 63163 70393
rect 63209 70347 63277 70393
rect 63323 70347 63391 70393
rect 63437 70347 63505 70393
rect 63551 70347 63619 70393
rect 63665 70347 63733 70393
rect 63779 70347 63847 70393
rect 63893 70347 63961 70393
rect 64007 70347 64075 70393
rect 64121 70347 64189 70393
rect 64235 70347 64303 70393
rect 64349 70347 64417 70393
rect 64463 70347 64531 70393
rect 64577 70347 64645 70393
rect 64691 70347 64759 70393
rect 64805 70347 64873 70393
rect 64919 70347 64987 70393
rect 65033 70347 65101 70393
rect 65147 70347 65215 70393
rect 65261 70347 65329 70393
rect 65375 70347 65443 70393
rect 65489 70347 65557 70393
rect 65603 70347 65671 70393
rect 65717 70347 65785 70393
rect 65831 70347 65899 70393
rect 65945 70347 66013 70393
rect 66059 70347 66127 70393
rect 66173 70347 66241 70393
rect 66287 70347 66355 70393
rect 66401 70347 66469 70393
rect 66515 70347 66583 70393
rect 66629 70347 66697 70393
rect 66743 70347 66811 70393
rect 66857 70347 66925 70393
rect 66971 70347 67039 70393
rect 67085 70347 67153 70393
rect 67199 70347 67267 70393
rect 67313 70347 67381 70393
rect 67427 70347 67495 70393
rect 67541 70347 67609 70393
rect 67655 70347 67723 70393
rect 67769 70347 67837 70393
rect 67883 70347 67951 70393
rect 67997 70347 68065 70393
rect 68111 70347 68179 70393
rect 68225 70347 68293 70393
rect 68339 70347 68407 70393
rect 68453 70347 68521 70393
rect 68567 70347 68635 70393
rect 68681 70347 68749 70393
rect 68795 70347 68863 70393
rect 68909 70347 68977 70393
rect 69023 70347 69091 70393
rect 69137 70347 69205 70393
rect 69251 70347 69319 70393
rect 69365 70347 69433 70393
rect 69479 70347 69501 70393
rect 60177 70279 69501 70347
rect 60177 70233 60199 70279
rect 60245 70233 60313 70279
rect 60359 70233 60427 70279
rect 60473 70233 60541 70279
rect 60587 70233 60655 70279
rect 60701 70233 60769 70279
rect 60815 70233 60883 70279
rect 60929 70233 60997 70279
rect 61043 70233 61111 70279
rect 61157 70233 61225 70279
rect 61271 70233 61339 70279
rect 61385 70233 61453 70279
rect 61499 70233 61567 70279
rect 61613 70233 61681 70279
rect 61727 70233 61795 70279
rect 61841 70233 61909 70279
rect 61955 70233 62023 70279
rect 62069 70233 62137 70279
rect 62183 70233 62251 70279
rect 62297 70233 62365 70279
rect 62411 70233 62479 70279
rect 62525 70233 62593 70279
rect 62639 70233 62707 70279
rect 62753 70233 62821 70279
rect 62867 70233 62935 70279
rect 62981 70233 63049 70279
rect 63095 70233 63163 70279
rect 63209 70233 63277 70279
rect 63323 70233 63391 70279
rect 63437 70233 63505 70279
rect 63551 70233 63619 70279
rect 63665 70233 63733 70279
rect 63779 70233 63847 70279
rect 63893 70233 63961 70279
rect 64007 70233 64075 70279
rect 64121 70233 64189 70279
rect 64235 70233 64303 70279
rect 64349 70233 64417 70279
rect 64463 70233 64531 70279
rect 64577 70233 64645 70279
rect 64691 70233 64759 70279
rect 64805 70233 64873 70279
rect 64919 70233 64987 70279
rect 65033 70233 65101 70279
rect 65147 70233 65215 70279
rect 65261 70233 65329 70279
rect 65375 70233 65443 70279
rect 65489 70233 65557 70279
rect 65603 70233 65671 70279
rect 65717 70233 65785 70279
rect 65831 70233 65899 70279
rect 65945 70233 66013 70279
rect 66059 70233 66127 70279
rect 66173 70233 66241 70279
rect 66287 70233 66355 70279
rect 66401 70233 66469 70279
rect 66515 70233 66583 70279
rect 66629 70233 66697 70279
rect 66743 70233 66811 70279
rect 66857 70233 66925 70279
rect 66971 70233 67039 70279
rect 67085 70233 67153 70279
rect 67199 70233 67267 70279
rect 67313 70233 67381 70279
rect 67427 70233 67495 70279
rect 67541 70233 67609 70279
rect 67655 70233 67723 70279
rect 67769 70233 67837 70279
rect 67883 70233 67951 70279
rect 67997 70233 68065 70279
rect 68111 70233 68179 70279
rect 68225 70233 68293 70279
rect 68339 70233 68407 70279
rect 68453 70233 68521 70279
rect 68567 70233 68635 70279
rect 68681 70233 68749 70279
rect 68795 70233 68863 70279
rect 68909 70233 68977 70279
rect 69023 70233 69091 70279
rect 69137 70233 69205 70279
rect 69251 70233 69319 70279
rect 69365 70233 69433 70279
rect 69479 70233 69501 70279
rect 60177 70165 69501 70233
rect 60177 70119 60199 70165
rect 60245 70119 60313 70165
rect 60359 70119 60427 70165
rect 60473 70119 60541 70165
rect 60587 70119 60655 70165
rect 60701 70119 60769 70165
rect 60815 70119 60883 70165
rect 60929 70119 60997 70165
rect 61043 70119 61111 70165
rect 61157 70119 61225 70165
rect 61271 70119 61339 70165
rect 61385 70119 61453 70165
rect 61499 70119 61567 70165
rect 61613 70119 61681 70165
rect 61727 70119 61795 70165
rect 61841 70119 61909 70165
rect 61955 70119 62023 70165
rect 62069 70119 62137 70165
rect 62183 70119 62251 70165
rect 62297 70119 62365 70165
rect 62411 70119 62479 70165
rect 62525 70119 62593 70165
rect 62639 70119 62707 70165
rect 62753 70119 62821 70165
rect 62867 70119 62935 70165
rect 62981 70119 63049 70165
rect 63095 70119 63163 70165
rect 63209 70119 63277 70165
rect 63323 70119 63391 70165
rect 63437 70119 63505 70165
rect 63551 70119 63619 70165
rect 63665 70119 63733 70165
rect 63779 70119 63847 70165
rect 63893 70119 63961 70165
rect 64007 70119 64075 70165
rect 64121 70119 64189 70165
rect 64235 70119 64303 70165
rect 64349 70119 64417 70165
rect 64463 70119 64531 70165
rect 64577 70119 64645 70165
rect 64691 70119 64759 70165
rect 64805 70119 64873 70165
rect 64919 70119 64987 70165
rect 65033 70119 65101 70165
rect 65147 70119 65215 70165
rect 65261 70119 65329 70165
rect 65375 70119 65443 70165
rect 65489 70119 65557 70165
rect 65603 70119 65671 70165
rect 65717 70119 65785 70165
rect 65831 70119 65899 70165
rect 65945 70119 66013 70165
rect 66059 70119 66127 70165
rect 66173 70119 66241 70165
rect 66287 70119 66355 70165
rect 66401 70119 66469 70165
rect 66515 70119 66583 70165
rect 66629 70119 66697 70165
rect 66743 70119 66811 70165
rect 66857 70119 66925 70165
rect 66971 70119 67039 70165
rect 67085 70119 67153 70165
rect 67199 70119 67267 70165
rect 67313 70119 67381 70165
rect 67427 70119 67495 70165
rect 67541 70119 67609 70165
rect 67655 70119 67723 70165
rect 67769 70119 67837 70165
rect 67883 70119 67951 70165
rect 67997 70119 68065 70165
rect 68111 70119 68179 70165
rect 68225 70119 68293 70165
rect 68339 70119 68407 70165
rect 68453 70119 68521 70165
rect 68567 70119 68635 70165
rect 68681 70119 68749 70165
rect 68795 70119 68863 70165
rect 68909 70119 68977 70165
rect 69023 70119 69091 70165
rect 69137 70119 69205 70165
rect 69251 70119 69319 70165
rect 69365 70119 69433 70165
rect 69479 70119 69501 70165
rect 60177 70051 69501 70119
rect 60177 70005 60199 70051
rect 60245 70005 60313 70051
rect 60359 70005 60427 70051
rect 60473 70005 60541 70051
rect 60587 70005 60655 70051
rect 60701 70005 60769 70051
rect 60815 70005 60883 70051
rect 60929 70005 60997 70051
rect 61043 70005 61111 70051
rect 61157 70005 61225 70051
rect 61271 70005 61339 70051
rect 61385 70005 61453 70051
rect 61499 70005 61567 70051
rect 61613 70005 61681 70051
rect 61727 70005 61795 70051
rect 61841 70005 61909 70051
rect 61955 70005 62023 70051
rect 62069 70005 62137 70051
rect 62183 70005 62251 70051
rect 62297 70005 62365 70051
rect 62411 70005 62479 70051
rect 62525 70005 62593 70051
rect 62639 70005 62707 70051
rect 62753 70005 62821 70051
rect 62867 70005 62935 70051
rect 62981 70005 63049 70051
rect 63095 70005 63163 70051
rect 63209 70005 63277 70051
rect 63323 70005 63391 70051
rect 63437 70005 63505 70051
rect 63551 70005 63619 70051
rect 63665 70005 63733 70051
rect 63779 70005 63847 70051
rect 63893 70005 63961 70051
rect 64007 70005 64075 70051
rect 64121 70005 64189 70051
rect 64235 70005 64303 70051
rect 64349 70005 64417 70051
rect 64463 70005 64531 70051
rect 64577 70005 64645 70051
rect 64691 70005 64759 70051
rect 64805 70005 64873 70051
rect 64919 70005 64987 70051
rect 65033 70005 65101 70051
rect 65147 70005 65215 70051
rect 65261 70005 65329 70051
rect 65375 70005 65443 70051
rect 65489 70005 65557 70051
rect 65603 70005 65671 70051
rect 65717 70005 65785 70051
rect 65831 70005 65899 70051
rect 65945 70005 66013 70051
rect 66059 70005 66127 70051
rect 66173 70005 66241 70051
rect 66287 70005 66355 70051
rect 66401 70005 66469 70051
rect 66515 70005 66583 70051
rect 66629 70005 66697 70051
rect 66743 70005 66811 70051
rect 66857 70005 66925 70051
rect 66971 70005 67039 70051
rect 67085 70005 67153 70051
rect 67199 70005 67267 70051
rect 67313 70005 67381 70051
rect 67427 70005 67495 70051
rect 67541 70005 67609 70051
rect 67655 70005 67723 70051
rect 67769 70005 67837 70051
rect 67883 70005 67951 70051
rect 67997 70005 68065 70051
rect 68111 70005 68179 70051
rect 68225 70005 68293 70051
rect 68339 70005 68407 70051
rect 68453 70005 68521 70051
rect 68567 70005 68635 70051
rect 68681 70005 68749 70051
rect 68795 70005 68863 70051
rect 68909 70005 68977 70051
rect 69023 70005 69091 70051
rect 69137 70005 69205 70051
rect 69251 70005 69319 70051
rect 69365 70005 69433 70051
rect 69479 70005 69501 70051
rect 60177 69937 69501 70005
rect 60177 69891 60199 69937
rect 60245 69891 60313 69937
rect 60359 69891 60427 69937
rect 60473 69891 60541 69937
rect 60587 69891 60655 69937
rect 60701 69891 60769 69937
rect 60815 69891 60883 69937
rect 60929 69891 60997 69937
rect 61043 69891 61111 69937
rect 61157 69891 61225 69937
rect 61271 69891 61339 69937
rect 61385 69891 61453 69937
rect 61499 69891 61567 69937
rect 61613 69891 61681 69937
rect 61727 69891 61795 69937
rect 61841 69891 61909 69937
rect 61955 69891 62023 69937
rect 62069 69891 62137 69937
rect 62183 69891 62251 69937
rect 62297 69891 62365 69937
rect 62411 69891 62479 69937
rect 62525 69891 62593 69937
rect 62639 69891 62707 69937
rect 62753 69891 62821 69937
rect 62867 69891 62935 69937
rect 62981 69891 63049 69937
rect 63095 69891 63163 69937
rect 63209 69891 63277 69937
rect 63323 69891 63391 69937
rect 63437 69891 63505 69937
rect 63551 69891 63619 69937
rect 63665 69891 63733 69937
rect 63779 69891 63847 69937
rect 63893 69891 63961 69937
rect 64007 69891 64075 69937
rect 64121 69891 64189 69937
rect 64235 69891 64303 69937
rect 64349 69891 64417 69937
rect 64463 69891 64531 69937
rect 64577 69891 64645 69937
rect 64691 69891 64759 69937
rect 64805 69891 64873 69937
rect 64919 69891 64987 69937
rect 65033 69891 65101 69937
rect 65147 69891 65215 69937
rect 65261 69891 65329 69937
rect 65375 69891 65443 69937
rect 65489 69891 65557 69937
rect 65603 69891 65671 69937
rect 65717 69891 65785 69937
rect 65831 69891 65899 69937
rect 65945 69891 66013 69937
rect 66059 69891 66127 69937
rect 66173 69891 66241 69937
rect 66287 69891 66355 69937
rect 66401 69891 66469 69937
rect 66515 69891 66583 69937
rect 66629 69891 66697 69937
rect 66743 69891 66811 69937
rect 66857 69891 66925 69937
rect 66971 69891 67039 69937
rect 67085 69891 67153 69937
rect 67199 69891 67267 69937
rect 67313 69891 67381 69937
rect 67427 69891 67495 69937
rect 67541 69891 67609 69937
rect 67655 69891 67723 69937
rect 67769 69891 67837 69937
rect 67883 69891 67951 69937
rect 67997 69891 68065 69937
rect 68111 69891 68179 69937
rect 68225 69891 68293 69937
rect 68339 69891 68407 69937
rect 68453 69891 68521 69937
rect 68567 69891 68635 69937
rect 68681 69891 68749 69937
rect 68795 69891 68863 69937
rect 68909 69891 68977 69937
rect 69023 69891 69091 69937
rect 69137 69891 69205 69937
rect 69251 69891 69319 69937
rect 69365 69891 69433 69937
rect 69479 69891 69501 69937
rect 60177 69823 69501 69891
rect 60177 69777 60199 69823
rect 60245 69777 60313 69823
rect 60359 69777 60427 69823
rect 60473 69777 60541 69823
rect 60587 69777 60655 69823
rect 60701 69777 60769 69823
rect 60815 69777 60883 69823
rect 60929 69777 60997 69823
rect 61043 69777 61111 69823
rect 61157 69777 61225 69823
rect 61271 69777 61339 69823
rect 61385 69777 61453 69823
rect 61499 69777 61567 69823
rect 61613 69777 61681 69823
rect 61727 69777 61795 69823
rect 61841 69777 61909 69823
rect 61955 69777 62023 69823
rect 62069 69777 62137 69823
rect 62183 69777 62251 69823
rect 62297 69777 62365 69823
rect 62411 69777 62479 69823
rect 62525 69777 62593 69823
rect 62639 69777 62707 69823
rect 62753 69777 62821 69823
rect 62867 69777 62935 69823
rect 62981 69777 63049 69823
rect 63095 69777 63163 69823
rect 63209 69777 63277 69823
rect 63323 69777 63391 69823
rect 63437 69777 63505 69823
rect 63551 69777 63619 69823
rect 63665 69777 63733 69823
rect 63779 69777 63847 69823
rect 63893 69777 63961 69823
rect 64007 69777 64075 69823
rect 64121 69777 64189 69823
rect 64235 69777 64303 69823
rect 64349 69777 64417 69823
rect 64463 69777 64531 69823
rect 64577 69777 64645 69823
rect 64691 69777 64759 69823
rect 64805 69777 64873 69823
rect 64919 69777 64987 69823
rect 65033 69777 65101 69823
rect 65147 69777 65215 69823
rect 65261 69777 65329 69823
rect 65375 69777 65443 69823
rect 65489 69777 65557 69823
rect 65603 69777 65671 69823
rect 65717 69777 65785 69823
rect 65831 69777 65899 69823
rect 65945 69777 66013 69823
rect 66059 69777 66127 69823
rect 66173 69777 66241 69823
rect 66287 69777 66355 69823
rect 66401 69777 66469 69823
rect 66515 69777 66583 69823
rect 66629 69777 66697 69823
rect 66743 69777 66811 69823
rect 66857 69777 66925 69823
rect 66971 69777 67039 69823
rect 67085 69777 67153 69823
rect 67199 69777 67267 69823
rect 67313 69777 67381 69823
rect 67427 69777 67495 69823
rect 67541 69777 67609 69823
rect 67655 69777 67723 69823
rect 67769 69777 67837 69823
rect 67883 69777 67951 69823
rect 67997 69777 68065 69823
rect 68111 69777 68179 69823
rect 68225 69777 68293 69823
rect 68339 69777 68407 69823
rect 68453 69777 68521 69823
rect 68567 69777 68635 69823
rect 68681 69777 68749 69823
rect 68795 69777 68863 69823
rect 68909 69777 68977 69823
rect 69023 69777 69091 69823
rect 69137 69777 69205 69823
rect 69251 69777 69319 69823
rect 69365 69777 69433 69823
rect 69479 69777 69501 69823
rect 60177 69709 69501 69777
rect 60177 69663 60199 69709
rect 60245 69663 60313 69709
rect 60359 69663 60427 69709
rect 60473 69663 60541 69709
rect 60587 69663 60655 69709
rect 60701 69663 60769 69709
rect 60815 69663 60883 69709
rect 60929 69663 60997 69709
rect 61043 69663 61111 69709
rect 61157 69663 61225 69709
rect 61271 69663 61339 69709
rect 61385 69663 61453 69709
rect 61499 69663 61567 69709
rect 61613 69663 61681 69709
rect 61727 69663 61795 69709
rect 61841 69663 61909 69709
rect 61955 69663 62023 69709
rect 62069 69663 62137 69709
rect 62183 69663 62251 69709
rect 62297 69663 62365 69709
rect 62411 69663 62479 69709
rect 62525 69663 62593 69709
rect 62639 69663 62707 69709
rect 62753 69663 62821 69709
rect 62867 69663 62935 69709
rect 62981 69663 63049 69709
rect 63095 69663 63163 69709
rect 63209 69663 63277 69709
rect 63323 69663 63391 69709
rect 63437 69663 63505 69709
rect 63551 69663 63619 69709
rect 63665 69663 63733 69709
rect 63779 69663 63847 69709
rect 63893 69663 63961 69709
rect 64007 69663 64075 69709
rect 64121 69663 64189 69709
rect 64235 69663 64303 69709
rect 64349 69663 64417 69709
rect 64463 69663 64531 69709
rect 64577 69663 64645 69709
rect 64691 69663 64759 69709
rect 64805 69663 64873 69709
rect 64919 69663 64987 69709
rect 65033 69663 65101 69709
rect 65147 69663 65215 69709
rect 65261 69663 65329 69709
rect 65375 69663 65443 69709
rect 65489 69663 65557 69709
rect 65603 69663 65671 69709
rect 65717 69663 65785 69709
rect 65831 69663 65899 69709
rect 65945 69663 66013 69709
rect 66059 69663 66127 69709
rect 66173 69663 66241 69709
rect 66287 69663 66355 69709
rect 66401 69663 66469 69709
rect 66515 69663 66583 69709
rect 66629 69663 66697 69709
rect 66743 69663 66811 69709
rect 66857 69663 66925 69709
rect 66971 69663 67039 69709
rect 67085 69663 67153 69709
rect 67199 69663 67267 69709
rect 67313 69663 67381 69709
rect 67427 69663 67495 69709
rect 67541 69663 67609 69709
rect 67655 69663 67723 69709
rect 67769 69663 67837 69709
rect 67883 69663 67951 69709
rect 67997 69663 68065 69709
rect 68111 69663 68179 69709
rect 68225 69663 68293 69709
rect 68339 69663 68407 69709
rect 68453 69663 68521 69709
rect 68567 69663 68635 69709
rect 68681 69663 68749 69709
rect 68795 69663 68863 69709
rect 68909 69663 68977 69709
rect 69023 69663 69091 69709
rect 69137 69663 69205 69709
rect 69251 69663 69319 69709
rect 69365 69663 69433 69709
rect 69479 69663 69501 69709
rect 60177 69595 69501 69663
rect 60177 69549 60199 69595
rect 60245 69549 60313 69595
rect 60359 69549 60427 69595
rect 60473 69549 60541 69595
rect 60587 69549 60655 69595
rect 60701 69549 60769 69595
rect 60815 69549 60883 69595
rect 60929 69549 60997 69595
rect 61043 69549 61111 69595
rect 61157 69549 61225 69595
rect 61271 69549 61339 69595
rect 61385 69549 61453 69595
rect 61499 69549 61567 69595
rect 61613 69549 61681 69595
rect 61727 69549 61795 69595
rect 61841 69549 61909 69595
rect 61955 69549 62023 69595
rect 62069 69549 62137 69595
rect 62183 69549 62251 69595
rect 62297 69549 62365 69595
rect 62411 69549 62479 69595
rect 62525 69549 62593 69595
rect 62639 69549 62707 69595
rect 62753 69549 62821 69595
rect 62867 69549 62935 69595
rect 62981 69549 63049 69595
rect 63095 69549 63163 69595
rect 63209 69549 63277 69595
rect 63323 69549 63391 69595
rect 63437 69549 63505 69595
rect 63551 69549 63619 69595
rect 63665 69549 63733 69595
rect 63779 69549 63847 69595
rect 63893 69549 63961 69595
rect 64007 69549 64075 69595
rect 64121 69549 64189 69595
rect 64235 69549 64303 69595
rect 64349 69549 64417 69595
rect 64463 69549 64531 69595
rect 64577 69549 64645 69595
rect 64691 69549 64759 69595
rect 64805 69549 64873 69595
rect 64919 69549 64987 69595
rect 65033 69549 65101 69595
rect 65147 69549 65215 69595
rect 65261 69549 65329 69595
rect 65375 69549 65443 69595
rect 65489 69549 65557 69595
rect 65603 69549 65671 69595
rect 65717 69549 65785 69595
rect 65831 69549 65899 69595
rect 65945 69549 66013 69595
rect 66059 69549 66127 69595
rect 66173 69549 66241 69595
rect 66287 69549 66355 69595
rect 66401 69549 66469 69595
rect 66515 69549 66583 69595
rect 66629 69549 66697 69595
rect 66743 69549 66811 69595
rect 66857 69549 66925 69595
rect 66971 69549 67039 69595
rect 67085 69549 67153 69595
rect 67199 69549 67267 69595
rect 67313 69549 67381 69595
rect 67427 69549 67495 69595
rect 67541 69549 67609 69595
rect 67655 69549 67723 69595
rect 67769 69549 67837 69595
rect 67883 69549 67951 69595
rect 67997 69549 68065 69595
rect 68111 69549 68179 69595
rect 68225 69549 68293 69595
rect 68339 69549 68407 69595
rect 68453 69549 68521 69595
rect 68567 69549 68635 69595
rect 68681 69549 68749 69595
rect 68795 69549 68863 69595
rect 68909 69549 68977 69595
rect 69023 69549 69091 69595
rect 69137 69549 69205 69595
rect 69251 69549 69319 69595
rect 69365 69549 69433 69595
rect 69479 69549 69501 69595
rect 60177 69481 69501 69549
rect 60177 69435 60199 69481
rect 60245 69435 60313 69481
rect 60359 69435 60427 69481
rect 60473 69435 60541 69481
rect 60587 69435 60655 69481
rect 60701 69435 60769 69481
rect 60815 69435 60883 69481
rect 60929 69435 60997 69481
rect 61043 69435 61111 69481
rect 61157 69435 61225 69481
rect 61271 69435 61339 69481
rect 61385 69435 61453 69481
rect 61499 69435 61567 69481
rect 61613 69435 61681 69481
rect 61727 69435 61795 69481
rect 61841 69435 61909 69481
rect 61955 69435 62023 69481
rect 62069 69435 62137 69481
rect 62183 69435 62251 69481
rect 62297 69435 62365 69481
rect 62411 69435 62479 69481
rect 62525 69435 62593 69481
rect 62639 69435 62707 69481
rect 62753 69435 62821 69481
rect 62867 69435 62935 69481
rect 62981 69435 63049 69481
rect 63095 69435 63163 69481
rect 63209 69435 63277 69481
rect 63323 69435 63391 69481
rect 63437 69435 63505 69481
rect 63551 69435 63619 69481
rect 63665 69435 63733 69481
rect 63779 69435 63847 69481
rect 63893 69435 63961 69481
rect 64007 69435 64075 69481
rect 64121 69435 64189 69481
rect 64235 69435 64303 69481
rect 64349 69435 64417 69481
rect 64463 69435 64531 69481
rect 64577 69435 64645 69481
rect 64691 69435 64759 69481
rect 64805 69435 64873 69481
rect 64919 69435 64987 69481
rect 65033 69435 65101 69481
rect 65147 69435 65215 69481
rect 65261 69435 65329 69481
rect 65375 69435 65443 69481
rect 65489 69435 65557 69481
rect 65603 69435 65671 69481
rect 65717 69435 65785 69481
rect 65831 69435 65899 69481
rect 65945 69435 66013 69481
rect 66059 69435 66127 69481
rect 66173 69435 66241 69481
rect 66287 69435 66355 69481
rect 66401 69435 66469 69481
rect 66515 69435 66583 69481
rect 66629 69435 66697 69481
rect 66743 69435 66811 69481
rect 66857 69435 66925 69481
rect 66971 69435 67039 69481
rect 67085 69435 67153 69481
rect 67199 69435 67267 69481
rect 67313 69435 67381 69481
rect 67427 69435 67495 69481
rect 67541 69435 67609 69481
rect 67655 69435 67723 69481
rect 67769 69435 67837 69481
rect 67883 69435 67951 69481
rect 67997 69435 68065 69481
rect 68111 69435 68179 69481
rect 68225 69435 68293 69481
rect 68339 69435 68407 69481
rect 68453 69435 68521 69481
rect 68567 69435 68635 69481
rect 68681 69435 68749 69481
rect 68795 69435 68863 69481
rect 68909 69435 68977 69481
rect 69023 69435 69091 69481
rect 69137 69435 69205 69481
rect 69251 69435 69319 69481
rect 69365 69435 69433 69481
rect 69479 69435 69501 69481
rect 60177 69367 69501 69435
rect 60177 69321 60199 69367
rect 60245 69321 60313 69367
rect 60359 69321 60427 69367
rect 60473 69321 60541 69367
rect 60587 69321 60655 69367
rect 60701 69321 60769 69367
rect 60815 69321 60883 69367
rect 60929 69321 60997 69367
rect 61043 69321 61111 69367
rect 61157 69321 61225 69367
rect 61271 69321 61339 69367
rect 61385 69321 61453 69367
rect 61499 69321 61567 69367
rect 61613 69321 61681 69367
rect 61727 69321 61795 69367
rect 61841 69321 61909 69367
rect 61955 69321 62023 69367
rect 62069 69321 62137 69367
rect 62183 69321 62251 69367
rect 62297 69321 62365 69367
rect 62411 69321 62479 69367
rect 62525 69321 62593 69367
rect 62639 69321 62707 69367
rect 62753 69321 62821 69367
rect 62867 69321 62935 69367
rect 62981 69321 63049 69367
rect 63095 69321 63163 69367
rect 63209 69321 63277 69367
rect 63323 69321 63391 69367
rect 63437 69321 63505 69367
rect 63551 69321 63619 69367
rect 63665 69321 63733 69367
rect 63779 69321 63847 69367
rect 63893 69321 63961 69367
rect 64007 69321 64075 69367
rect 64121 69321 64189 69367
rect 64235 69321 64303 69367
rect 64349 69321 64417 69367
rect 64463 69321 64531 69367
rect 64577 69321 64645 69367
rect 64691 69321 64759 69367
rect 64805 69321 64873 69367
rect 64919 69321 64987 69367
rect 65033 69321 65101 69367
rect 65147 69321 65215 69367
rect 65261 69321 65329 69367
rect 65375 69321 65443 69367
rect 65489 69321 65557 69367
rect 65603 69321 65671 69367
rect 65717 69321 65785 69367
rect 65831 69321 65899 69367
rect 65945 69321 66013 69367
rect 66059 69321 66127 69367
rect 66173 69321 66241 69367
rect 66287 69321 66355 69367
rect 66401 69321 66469 69367
rect 66515 69321 66583 69367
rect 66629 69321 66697 69367
rect 66743 69321 66811 69367
rect 66857 69321 66925 69367
rect 66971 69321 67039 69367
rect 67085 69321 67153 69367
rect 67199 69321 67267 69367
rect 67313 69321 67381 69367
rect 67427 69321 67495 69367
rect 67541 69321 67609 69367
rect 67655 69321 67723 69367
rect 67769 69321 67837 69367
rect 67883 69321 67951 69367
rect 67997 69321 68065 69367
rect 68111 69321 68179 69367
rect 68225 69321 68293 69367
rect 68339 69321 68407 69367
rect 68453 69321 68521 69367
rect 68567 69321 68635 69367
rect 68681 69321 68749 69367
rect 68795 69321 68863 69367
rect 68909 69321 68977 69367
rect 69023 69321 69091 69367
rect 69137 69321 69205 69367
rect 69251 69321 69319 69367
rect 69365 69321 69433 69367
rect 69479 69321 69501 69367
rect 60177 69253 69501 69321
rect 60177 69207 60199 69253
rect 60245 69207 60313 69253
rect 60359 69207 60427 69253
rect 60473 69207 60541 69253
rect 60587 69207 60655 69253
rect 60701 69207 60769 69253
rect 60815 69207 60883 69253
rect 60929 69207 60997 69253
rect 61043 69207 61111 69253
rect 61157 69207 61225 69253
rect 61271 69207 61339 69253
rect 61385 69207 61453 69253
rect 61499 69207 61567 69253
rect 61613 69207 61681 69253
rect 61727 69207 61795 69253
rect 61841 69207 61909 69253
rect 61955 69207 62023 69253
rect 62069 69207 62137 69253
rect 62183 69207 62251 69253
rect 62297 69207 62365 69253
rect 62411 69207 62479 69253
rect 62525 69207 62593 69253
rect 62639 69207 62707 69253
rect 62753 69207 62821 69253
rect 62867 69207 62935 69253
rect 62981 69207 63049 69253
rect 63095 69207 63163 69253
rect 63209 69207 63277 69253
rect 63323 69207 63391 69253
rect 63437 69207 63505 69253
rect 63551 69207 63619 69253
rect 63665 69207 63733 69253
rect 63779 69207 63847 69253
rect 63893 69207 63961 69253
rect 64007 69207 64075 69253
rect 64121 69207 64189 69253
rect 64235 69207 64303 69253
rect 64349 69207 64417 69253
rect 64463 69207 64531 69253
rect 64577 69207 64645 69253
rect 64691 69207 64759 69253
rect 64805 69207 64873 69253
rect 64919 69207 64987 69253
rect 65033 69207 65101 69253
rect 65147 69207 65215 69253
rect 65261 69207 65329 69253
rect 65375 69207 65443 69253
rect 65489 69207 65557 69253
rect 65603 69207 65671 69253
rect 65717 69207 65785 69253
rect 65831 69207 65899 69253
rect 65945 69207 66013 69253
rect 66059 69207 66127 69253
rect 66173 69207 66241 69253
rect 66287 69207 66355 69253
rect 66401 69207 66469 69253
rect 66515 69207 66583 69253
rect 66629 69207 66697 69253
rect 66743 69207 66811 69253
rect 66857 69207 66925 69253
rect 66971 69207 67039 69253
rect 67085 69207 67153 69253
rect 67199 69207 67267 69253
rect 67313 69207 67381 69253
rect 67427 69207 67495 69253
rect 67541 69207 67609 69253
rect 67655 69207 67723 69253
rect 67769 69207 67837 69253
rect 67883 69207 67951 69253
rect 67997 69207 68065 69253
rect 68111 69207 68179 69253
rect 68225 69207 68293 69253
rect 68339 69207 68407 69253
rect 68453 69207 68521 69253
rect 68567 69207 68635 69253
rect 68681 69207 68749 69253
rect 68795 69207 68863 69253
rect 68909 69207 68977 69253
rect 69023 69207 69091 69253
rect 69137 69207 69205 69253
rect 69251 69207 69319 69253
rect 69365 69207 69433 69253
rect 69479 69207 69501 69253
rect 60177 69139 69501 69207
rect 60177 69093 60199 69139
rect 60245 69093 60313 69139
rect 60359 69093 60427 69139
rect 60473 69093 60541 69139
rect 60587 69093 60655 69139
rect 60701 69093 60769 69139
rect 60815 69093 60883 69139
rect 60929 69093 60997 69139
rect 61043 69093 61111 69139
rect 61157 69093 61225 69139
rect 61271 69093 61339 69139
rect 61385 69093 61453 69139
rect 61499 69093 61567 69139
rect 61613 69093 61681 69139
rect 61727 69093 61795 69139
rect 61841 69093 61909 69139
rect 61955 69093 62023 69139
rect 62069 69093 62137 69139
rect 62183 69093 62251 69139
rect 62297 69093 62365 69139
rect 62411 69093 62479 69139
rect 62525 69093 62593 69139
rect 62639 69093 62707 69139
rect 62753 69093 62821 69139
rect 62867 69093 62935 69139
rect 62981 69093 63049 69139
rect 63095 69093 63163 69139
rect 63209 69093 63277 69139
rect 63323 69093 63391 69139
rect 63437 69093 63505 69139
rect 63551 69093 63619 69139
rect 63665 69093 63733 69139
rect 63779 69093 63847 69139
rect 63893 69093 63961 69139
rect 64007 69093 64075 69139
rect 64121 69093 64189 69139
rect 64235 69093 64303 69139
rect 64349 69093 64417 69139
rect 64463 69093 64531 69139
rect 64577 69093 64645 69139
rect 64691 69093 64759 69139
rect 64805 69093 64873 69139
rect 64919 69093 64987 69139
rect 65033 69093 65101 69139
rect 65147 69093 65215 69139
rect 65261 69093 65329 69139
rect 65375 69093 65443 69139
rect 65489 69093 65557 69139
rect 65603 69093 65671 69139
rect 65717 69093 65785 69139
rect 65831 69093 65899 69139
rect 65945 69093 66013 69139
rect 66059 69093 66127 69139
rect 66173 69093 66241 69139
rect 66287 69093 66355 69139
rect 66401 69093 66469 69139
rect 66515 69093 66583 69139
rect 66629 69093 66697 69139
rect 66743 69093 66811 69139
rect 66857 69093 66925 69139
rect 66971 69093 67039 69139
rect 67085 69093 67153 69139
rect 67199 69093 67267 69139
rect 67313 69093 67381 69139
rect 67427 69093 67495 69139
rect 67541 69093 67609 69139
rect 67655 69093 67723 69139
rect 67769 69093 67837 69139
rect 67883 69093 67951 69139
rect 67997 69093 68065 69139
rect 68111 69093 68179 69139
rect 68225 69093 68293 69139
rect 68339 69093 68407 69139
rect 68453 69093 68521 69139
rect 68567 69093 68635 69139
rect 68681 69093 68749 69139
rect 68795 69093 68863 69139
rect 68909 69093 68977 69139
rect 69023 69093 69091 69139
rect 69137 69093 69205 69139
rect 69251 69093 69319 69139
rect 69365 69093 69433 69139
rect 69479 69093 69501 69139
rect 60177 69025 69501 69093
rect 60177 68979 60199 69025
rect 60245 68979 60313 69025
rect 60359 68979 60427 69025
rect 60473 68979 60541 69025
rect 60587 68979 60655 69025
rect 60701 68979 60769 69025
rect 60815 68979 60883 69025
rect 60929 68979 60997 69025
rect 61043 68979 61111 69025
rect 61157 68979 61225 69025
rect 61271 68979 61339 69025
rect 61385 68979 61453 69025
rect 61499 68979 61567 69025
rect 61613 68979 61681 69025
rect 61727 68979 61795 69025
rect 61841 68979 61909 69025
rect 61955 68979 62023 69025
rect 62069 68979 62137 69025
rect 62183 68979 62251 69025
rect 62297 68979 62365 69025
rect 62411 68979 62479 69025
rect 62525 68979 62593 69025
rect 62639 68979 62707 69025
rect 62753 68979 62821 69025
rect 62867 68979 62935 69025
rect 62981 68979 63049 69025
rect 63095 68979 63163 69025
rect 63209 68979 63277 69025
rect 63323 68979 63391 69025
rect 63437 68979 63505 69025
rect 63551 68979 63619 69025
rect 63665 68979 63733 69025
rect 63779 68979 63847 69025
rect 63893 68979 63961 69025
rect 64007 68979 64075 69025
rect 64121 68979 64189 69025
rect 64235 68979 64303 69025
rect 64349 68979 64417 69025
rect 64463 68979 64531 69025
rect 64577 68979 64645 69025
rect 64691 68979 64759 69025
rect 64805 68979 64873 69025
rect 64919 68979 64987 69025
rect 65033 68979 65101 69025
rect 65147 68979 65215 69025
rect 65261 68979 65329 69025
rect 65375 68979 65443 69025
rect 65489 68979 65557 69025
rect 65603 68979 65671 69025
rect 65717 68979 65785 69025
rect 65831 68979 65899 69025
rect 65945 68979 66013 69025
rect 66059 68979 66127 69025
rect 66173 68979 66241 69025
rect 66287 68979 66355 69025
rect 66401 68979 66469 69025
rect 66515 68979 66583 69025
rect 66629 68979 66697 69025
rect 66743 68979 66811 69025
rect 66857 68979 66925 69025
rect 66971 68979 67039 69025
rect 67085 68979 67153 69025
rect 67199 68979 67267 69025
rect 67313 68979 67381 69025
rect 67427 68979 67495 69025
rect 67541 68979 67609 69025
rect 67655 68979 67723 69025
rect 67769 68979 67837 69025
rect 67883 68979 67951 69025
rect 67997 68979 68065 69025
rect 68111 68979 68179 69025
rect 68225 68979 68293 69025
rect 68339 68979 68407 69025
rect 68453 68979 68521 69025
rect 68567 68979 68635 69025
rect 68681 68979 68749 69025
rect 68795 68979 68863 69025
rect 68909 68979 68977 69025
rect 69023 68979 69091 69025
rect 69137 68979 69205 69025
rect 69251 68979 69319 69025
rect 69365 68979 69433 69025
rect 69479 68979 69501 69025
rect 60177 68957 69501 68979
<< psubdiffcont >>
rect 60199 70461 60245 70507
rect 60313 70461 60359 70507
rect 60427 70461 60473 70507
rect 60541 70461 60587 70507
rect 60655 70461 60701 70507
rect 60769 70461 60815 70507
rect 60883 70461 60929 70507
rect 60997 70461 61043 70507
rect 61111 70461 61157 70507
rect 61225 70461 61271 70507
rect 61339 70461 61385 70507
rect 61453 70461 61499 70507
rect 61567 70461 61613 70507
rect 61681 70461 61727 70507
rect 61795 70461 61841 70507
rect 61909 70461 61955 70507
rect 62023 70461 62069 70507
rect 62137 70461 62183 70507
rect 62251 70461 62297 70507
rect 62365 70461 62411 70507
rect 62479 70461 62525 70507
rect 62593 70461 62639 70507
rect 62707 70461 62753 70507
rect 62821 70461 62867 70507
rect 62935 70461 62981 70507
rect 63049 70461 63095 70507
rect 63163 70461 63209 70507
rect 63277 70461 63323 70507
rect 63391 70461 63437 70507
rect 63505 70461 63551 70507
rect 63619 70461 63665 70507
rect 63733 70461 63779 70507
rect 63847 70461 63893 70507
rect 63961 70461 64007 70507
rect 64075 70461 64121 70507
rect 64189 70461 64235 70507
rect 64303 70461 64349 70507
rect 64417 70461 64463 70507
rect 64531 70461 64577 70507
rect 64645 70461 64691 70507
rect 64759 70461 64805 70507
rect 64873 70461 64919 70507
rect 64987 70461 65033 70507
rect 65101 70461 65147 70507
rect 65215 70461 65261 70507
rect 65329 70461 65375 70507
rect 65443 70461 65489 70507
rect 65557 70461 65603 70507
rect 65671 70461 65717 70507
rect 65785 70461 65831 70507
rect 65899 70461 65945 70507
rect 66013 70461 66059 70507
rect 66127 70461 66173 70507
rect 66241 70461 66287 70507
rect 66355 70461 66401 70507
rect 66469 70461 66515 70507
rect 66583 70461 66629 70507
rect 66697 70461 66743 70507
rect 66811 70461 66857 70507
rect 66925 70461 66971 70507
rect 67039 70461 67085 70507
rect 67153 70461 67199 70507
rect 67267 70461 67313 70507
rect 67381 70461 67427 70507
rect 67495 70461 67541 70507
rect 67609 70461 67655 70507
rect 67723 70461 67769 70507
rect 67837 70461 67883 70507
rect 67951 70461 67997 70507
rect 68065 70461 68111 70507
rect 68179 70461 68225 70507
rect 68293 70461 68339 70507
rect 68407 70461 68453 70507
rect 68521 70461 68567 70507
rect 68635 70461 68681 70507
rect 68749 70461 68795 70507
rect 68863 70461 68909 70507
rect 68977 70461 69023 70507
rect 69091 70461 69137 70507
rect 69205 70461 69251 70507
rect 69319 70461 69365 70507
rect 69433 70461 69479 70507
rect 60199 70347 60245 70393
rect 60313 70347 60359 70393
rect 60427 70347 60473 70393
rect 60541 70347 60587 70393
rect 60655 70347 60701 70393
rect 60769 70347 60815 70393
rect 60883 70347 60929 70393
rect 60997 70347 61043 70393
rect 61111 70347 61157 70393
rect 61225 70347 61271 70393
rect 61339 70347 61385 70393
rect 61453 70347 61499 70393
rect 61567 70347 61613 70393
rect 61681 70347 61727 70393
rect 61795 70347 61841 70393
rect 61909 70347 61955 70393
rect 62023 70347 62069 70393
rect 62137 70347 62183 70393
rect 62251 70347 62297 70393
rect 62365 70347 62411 70393
rect 62479 70347 62525 70393
rect 62593 70347 62639 70393
rect 62707 70347 62753 70393
rect 62821 70347 62867 70393
rect 62935 70347 62981 70393
rect 63049 70347 63095 70393
rect 63163 70347 63209 70393
rect 63277 70347 63323 70393
rect 63391 70347 63437 70393
rect 63505 70347 63551 70393
rect 63619 70347 63665 70393
rect 63733 70347 63779 70393
rect 63847 70347 63893 70393
rect 63961 70347 64007 70393
rect 64075 70347 64121 70393
rect 64189 70347 64235 70393
rect 64303 70347 64349 70393
rect 64417 70347 64463 70393
rect 64531 70347 64577 70393
rect 64645 70347 64691 70393
rect 64759 70347 64805 70393
rect 64873 70347 64919 70393
rect 64987 70347 65033 70393
rect 65101 70347 65147 70393
rect 65215 70347 65261 70393
rect 65329 70347 65375 70393
rect 65443 70347 65489 70393
rect 65557 70347 65603 70393
rect 65671 70347 65717 70393
rect 65785 70347 65831 70393
rect 65899 70347 65945 70393
rect 66013 70347 66059 70393
rect 66127 70347 66173 70393
rect 66241 70347 66287 70393
rect 66355 70347 66401 70393
rect 66469 70347 66515 70393
rect 66583 70347 66629 70393
rect 66697 70347 66743 70393
rect 66811 70347 66857 70393
rect 66925 70347 66971 70393
rect 67039 70347 67085 70393
rect 67153 70347 67199 70393
rect 67267 70347 67313 70393
rect 67381 70347 67427 70393
rect 67495 70347 67541 70393
rect 67609 70347 67655 70393
rect 67723 70347 67769 70393
rect 67837 70347 67883 70393
rect 67951 70347 67997 70393
rect 68065 70347 68111 70393
rect 68179 70347 68225 70393
rect 68293 70347 68339 70393
rect 68407 70347 68453 70393
rect 68521 70347 68567 70393
rect 68635 70347 68681 70393
rect 68749 70347 68795 70393
rect 68863 70347 68909 70393
rect 68977 70347 69023 70393
rect 69091 70347 69137 70393
rect 69205 70347 69251 70393
rect 69319 70347 69365 70393
rect 69433 70347 69479 70393
rect 60199 70233 60245 70279
rect 60313 70233 60359 70279
rect 60427 70233 60473 70279
rect 60541 70233 60587 70279
rect 60655 70233 60701 70279
rect 60769 70233 60815 70279
rect 60883 70233 60929 70279
rect 60997 70233 61043 70279
rect 61111 70233 61157 70279
rect 61225 70233 61271 70279
rect 61339 70233 61385 70279
rect 61453 70233 61499 70279
rect 61567 70233 61613 70279
rect 61681 70233 61727 70279
rect 61795 70233 61841 70279
rect 61909 70233 61955 70279
rect 62023 70233 62069 70279
rect 62137 70233 62183 70279
rect 62251 70233 62297 70279
rect 62365 70233 62411 70279
rect 62479 70233 62525 70279
rect 62593 70233 62639 70279
rect 62707 70233 62753 70279
rect 62821 70233 62867 70279
rect 62935 70233 62981 70279
rect 63049 70233 63095 70279
rect 63163 70233 63209 70279
rect 63277 70233 63323 70279
rect 63391 70233 63437 70279
rect 63505 70233 63551 70279
rect 63619 70233 63665 70279
rect 63733 70233 63779 70279
rect 63847 70233 63893 70279
rect 63961 70233 64007 70279
rect 64075 70233 64121 70279
rect 64189 70233 64235 70279
rect 64303 70233 64349 70279
rect 64417 70233 64463 70279
rect 64531 70233 64577 70279
rect 64645 70233 64691 70279
rect 64759 70233 64805 70279
rect 64873 70233 64919 70279
rect 64987 70233 65033 70279
rect 65101 70233 65147 70279
rect 65215 70233 65261 70279
rect 65329 70233 65375 70279
rect 65443 70233 65489 70279
rect 65557 70233 65603 70279
rect 65671 70233 65717 70279
rect 65785 70233 65831 70279
rect 65899 70233 65945 70279
rect 66013 70233 66059 70279
rect 66127 70233 66173 70279
rect 66241 70233 66287 70279
rect 66355 70233 66401 70279
rect 66469 70233 66515 70279
rect 66583 70233 66629 70279
rect 66697 70233 66743 70279
rect 66811 70233 66857 70279
rect 66925 70233 66971 70279
rect 67039 70233 67085 70279
rect 67153 70233 67199 70279
rect 67267 70233 67313 70279
rect 67381 70233 67427 70279
rect 67495 70233 67541 70279
rect 67609 70233 67655 70279
rect 67723 70233 67769 70279
rect 67837 70233 67883 70279
rect 67951 70233 67997 70279
rect 68065 70233 68111 70279
rect 68179 70233 68225 70279
rect 68293 70233 68339 70279
rect 68407 70233 68453 70279
rect 68521 70233 68567 70279
rect 68635 70233 68681 70279
rect 68749 70233 68795 70279
rect 68863 70233 68909 70279
rect 68977 70233 69023 70279
rect 69091 70233 69137 70279
rect 69205 70233 69251 70279
rect 69319 70233 69365 70279
rect 69433 70233 69479 70279
rect 60199 70119 60245 70165
rect 60313 70119 60359 70165
rect 60427 70119 60473 70165
rect 60541 70119 60587 70165
rect 60655 70119 60701 70165
rect 60769 70119 60815 70165
rect 60883 70119 60929 70165
rect 60997 70119 61043 70165
rect 61111 70119 61157 70165
rect 61225 70119 61271 70165
rect 61339 70119 61385 70165
rect 61453 70119 61499 70165
rect 61567 70119 61613 70165
rect 61681 70119 61727 70165
rect 61795 70119 61841 70165
rect 61909 70119 61955 70165
rect 62023 70119 62069 70165
rect 62137 70119 62183 70165
rect 62251 70119 62297 70165
rect 62365 70119 62411 70165
rect 62479 70119 62525 70165
rect 62593 70119 62639 70165
rect 62707 70119 62753 70165
rect 62821 70119 62867 70165
rect 62935 70119 62981 70165
rect 63049 70119 63095 70165
rect 63163 70119 63209 70165
rect 63277 70119 63323 70165
rect 63391 70119 63437 70165
rect 63505 70119 63551 70165
rect 63619 70119 63665 70165
rect 63733 70119 63779 70165
rect 63847 70119 63893 70165
rect 63961 70119 64007 70165
rect 64075 70119 64121 70165
rect 64189 70119 64235 70165
rect 64303 70119 64349 70165
rect 64417 70119 64463 70165
rect 64531 70119 64577 70165
rect 64645 70119 64691 70165
rect 64759 70119 64805 70165
rect 64873 70119 64919 70165
rect 64987 70119 65033 70165
rect 65101 70119 65147 70165
rect 65215 70119 65261 70165
rect 65329 70119 65375 70165
rect 65443 70119 65489 70165
rect 65557 70119 65603 70165
rect 65671 70119 65717 70165
rect 65785 70119 65831 70165
rect 65899 70119 65945 70165
rect 66013 70119 66059 70165
rect 66127 70119 66173 70165
rect 66241 70119 66287 70165
rect 66355 70119 66401 70165
rect 66469 70119 66515 70165
rect 66583 70119 66629 70165
rect 66697 70119 66743 70165
rect 66811 70119 66857 70165
rect 66925 70119 66971 70165
rect 67039 70119 67085 70165
rect 67153 70119 67199 70165
rect 67267 70119 67313 70165
rect 67381 70119 67427 70165
rect 67495 70119 67541 70165
rect 67609 70119 67655 70165
rect 67723 70119 67769 70165
rect 67837 70119 67883 70165
rect 67951 70119 67997 70165
rect 68065 70119 68111 70165
rect 68179 70119 68225 70165
rect 68293 70119 68339 70165
rect 68407 70119 68453 70165
rect 68521 70119 68567 70165
rect 68635 70119 68681 70165
rect 68749 70119 68795 70165
rect 68863 70119 68909 70165
rect 68977 70119 69023 70165
rect 69091 70119 69137 70165
rect 69205 70119 69251 70165
rect 69319 70119 69365 70165
rect 69433 70119 69479 70165
rect 60199 70005 60245 70051
rect 60313 70005 60359 70051
rect 60427 70005 60473 70051
rect 60541 70005 60587 70051
rect 60655 70005 60701 70051
rect 60769 70005 60815 70051
rect 60883 70005 60929 70051
rect 60997 70005 61043 70051
rect 61111 70005 61157 70051
rect 61225 70005 61271 70051
rect 61339 70005 61385 70051
rect 61453 70005 61499 70051
rect 61567 70005 61613 70051
rect 61681 70005 61727 70051
rect 61795 70005 61841 70051
rect 61909 70005 61955 70051
rect 62023 70005 62069 70051
rect 62137 70005 62183 70051
rect 62251 70005 62297 70051
rect 62365 70005 62411 70051
rect 62479 70005 62525 70051
rect 62593 70005 62639 70051
rect 62707 70005 62753 70051
rect 62821 70005 62867 70051
rect 62935 70005 62981 70051
rect 63049 70005 63095 70051
rect 63163 70005 63209 70051
rect 63277 70005 63323 70051
rect 63391 70005 63437 70051
rect 63505 70005 63551 70051
rect 63619 70005 63665 70051
rect 63733 70005 63779 70051
rect 63847 70005 63893 70051
rect 63961 70005 64007 70051
rect 64075 70005 64121 70051
rect 64189 70005 64235 70051
rect 64303 70005 64349 70051
rect 64417 70005 64463 70051
rect 64531 70005 64577 70051
rect 64645 70005 64691 70051
rect 64759 70005 64805 70051
rect 64873 70005 64919 70051
rect 64987 70005 65033 70051
rect 65101 70005 65147 70051
rect 65215 70005 65261 70051
rect 65329 70005 65375 70051
rect 65443 70005 65489 70051
rect 65557 70005 65603 70051
rect 65671 70005 65717 70051
rect 65785 70005 65831 70051
rect 65899 70005 65945 70051
rect 66013 70005 66059 70051
rect 66127 70005 66173 70051
rect 66241 70005 66287 70051
rect 66355 70005 66401 70051
rect 66469 70005 66515 70051
rect 66583 70005 66629 70051
rect 66697 70005 66743 70051
rect 66811 70005 66857 70051
rect 66925 70005 66971 70051
rect 67039 70005 67085 70051
rect 67153 70005 67199 70051
rect 67267 70005 67313 70051
rect 67381 70005 67427 70051
rect 67495 70005 67541 70051
rect 67609 70005 67655 70051
rect 67723 70005 67769 70051
rect 67837 70005 67883 70051
rect 67951 70005 67997 70051
rect 68065 70005 68111 70051
rect 68179 70005 68225 70051
rect 68293 70005 68339 70051
rect 68407 70005 68453 70051
rect 68521 70005 68567 70051
rect 68635 70005 68681 70051
rect 68749 70005 68795 70051
rect 68863 70005 68909 70051
rect 68977 70005 69023 70051
rect 69091 70005 69137 70051
rect 69205 70005 69251 70051
rect 69319 70005 69365 70051
rect 69433 70005 69479 70051
rect 60199 69891 60245 69937
rect 60313 69891 60359 69937
rect 60427 69891 60473 69937
rect 60541 69891 60587 69937
rect 60655 69891 60701 69937
rect 60769 69891 60815 69937
rect 60883 69891 60929 69937
rect 60997 69891 61043 69937
rect 61111 69891 61157 69937
rect 61225 69891 61271 69937
rect 61339 69891 61385 69937
rect 61453 69891 61499 69937
rect 61567 69891 61613 69937
rect 61681 69891 61727 69937
rect 61795 69891 61841 69937
rect 61909 69891 61955 69937
rect 62023 69891 62069 69937
rect 62137 69891 62183 69937
rect 62251 69891 62297 69937
rect 62365 69891 62411 69937
rect 62479 69891 62525 69937
rect 62593 69891 62639 69937
rect 62707 69891 62753 69937
rect 62821 69891 62867 69937
rect 62935 69891 62981 69937
rect 63049 69891 63095 69937
rect 63163 69891 63209 69937
rect 63277 69891 63323 69937
rect 63391 69891 63437 69937
rect 63505 69891 63551 69937
rect 63619 69891 63665 69937
rect 63733 69891 63779 69937
rect 63847 69891 63893 69937
rect 63961 69891 64007 69937
rect 64075 69891 64121 69937
rect 64189 69891 64235 69937
rect 64303 69891 64349 69937
rect 64417 69891 64463 69937
rect 64531 69891 64577 69937
rect 64645 69891 64691 69937
rect 64759 69891 64805 69937
rect 64873 69891 64919 69937
rect 64987 69891 65033 69937
rect 65101 69891 65147 69937
rect 65215 69891 65261 69937
rect 65329 69891 65375 69937
rect 65443 69891 65489 69937
rect 65557 69891 65603 69937
rect 65671 69891 65717 69937
rect 65785 69891 65831 69937
rect 65899 69891 65945 69937
rect 66013 69891 66059 69937
rect 66127 69891 66173 69937
rect 66241 69891 66287 69937
rect 66355 69891 66401 69937
rect 66469 69891 66515 69937
rect 66583 69891 66629 69937
rect 66697 69891 66743 69937
rect 66811 69891 66857 69937
rect 66925 69891 66971 69937
rect 67039 69891 67085 69937
rect 67153 69891 67199 69937
rect 67267 69891 67313 69937
rect 67381 69891 67427 69937
rect 67495 69891 67541 69937
rect 67609 69891 67655 69937
rect 67723 69891 67769 69937
rect 67837 69891 67883 69937
rect 67951 69891 67997 69937
rect 68065 69891 68111 69937
rect 68179 69891 68225 69937
rect 68293 69891 68339 69937
rect 68407 69891 68453 69937
rect 68521 69891 68567 69937
rect 68635 69891 68681 69937
rect 68749 69891 68795 69937
rect 68863 69891 68909 69937
rect 68977 69891 69023 69937
rect 69091 69891 69137 69937
rect 69205 69891 69251 69937
rect 69319 69891 69365 69937
rect 69433 69891 69479 69937
rect 60199 69777 60245 69823
rect 60313 69777 60359 69823
rect 60427 69777 60473 69823
rect 60541 69777 60587 69823
rect 60655 69777 60701 69823
rect 60769 69777 60815 69823
rect 60883 69777 60929 69823
rect 60997 69777 61043 69823
rect 61111 69777 61157 69823
rect 61225 69777 61271 69823
rect 61339 69777 61385 69823
rect 61453 69777 61499 69823
rect 61567 69777 61613 69823
rect 61681 69777 61727 69823
rect 61795 69777 61841 69823
rect 61909 69777 61955 69823
rect 62023 69777 62069 69823
rect 62137 69777 62183 69823
rect 62251 69777 62297 69823
rect 62365 69777 62411 69823
rect 62479 69777 62525 69823
rect 62593 69777 62639 69823
rect 62707 69777 62753 69823
rect 62821 69777 62867 69823
rect 62935 69777 62981 69823
rect 63049 69777 63095 69823
rect 63163 69777 63209 69823
rect 63277 69777 63323 69823
rect 63391 69777 63437 69823
rect 63505 69777 63551 69823
rect 63619 69777 63665 69823
rect 63733 69777 63779 69823
rect 63847 69777 63893 69823
rect 63961 69777 64007 69823
rect 64075 69777 64121 69823
rect 64189 69777 64235 69823
rect 64303 69777 64349 69823
rect 64417 69777 64463 69823
rect 64531 69777 64577 69823
rect 64645 69777 64691 69823
rect 64759 69777 64805 69823
rect 64873 69777 64919 69823
rect 64987 69777 65033 69823
rect 65101 69777 65147 69823
rect 65215 69777 65261 69823
rect 65329 69777 65375 69823
rect 65443 69777 65489 69823
rect 65557 69777 65603 69823
rect 65671 69777 65717 69823
rect 65785 69777 65831 69823
rect 65899 69777 65945 69823
rect 66013 69777 66059 69823
rect 66127 69777 66173 69823
rect 66241 69777 66287 69823
rect 66355 69777 66401 69823
rect 66469 69777 66515 69823
rect 66583 69777 66629 69823
rect 66697 69777 66743 69823
rect 66811 69777 66857 69823
rect 66925 69777 66971 69823
rect 67039 69777 67085 69823
rect 67153 69777 67199 69823
rect 67267 69777 67313 69823
rect 67381 69777 67427 69823
rect 67495 69777 67541 69823
rect 67609 69777 67655 69823
rect 67723 69777 67769 69823
rect 67837 69777 67883 69823
rect 67951 69777 67997 69823
rect 68065 69777 68111 69823
rect 68179 69777 68225 69823
rect 68293 69777 68339 69823
rect 68407 69777 68453 69823
rect 68521 69777 68567 69823
rect 68635 69777 68681 69823
rect 68749 69777 68795 69823
rect 68863 69777 68909 69823
rect 68977 69777 69023 69823
rect 69091 69777 69137 69823
rect 69205 69777 69251 69823
rect 69319 69777 69365 69823
rect 69433 69777 69479 69823
rect 60199 69663 60245 69709
rect 60313 69663 60359 69709
rect 60427 69663 60473 69709
rect 60541 69663 60587 69709
rect 60655 69663 60701 69709
rect 60769 69663 60815 69709
rect 60883 69663 60929 69709
rect 60997 69663 61043 69709
rect 61111 69663 61157 69709
rect 61225 69663 61271 69709
rect 61339 69663 61385 69709
rect 61453 69663 61499 69709
rect 61567 69663 61613 69709
rect 61681 69663 61727 69709
rect 61795 69663 61841 69709
rect 61909 69663 61955 69709
rect 62023 69663 62069 69709
rect 62137 69663 62183 69709
rect 62251 69663 62297 69709
rect 62365 69663 62411 69709
rect 62479 69663 62525 69709
rect 62593 69663 62639 69709
rect 62707 69663 62753 69709
rect 62821 69663 62867 69709
rect 62935 69663 62981 69709
rect 63049 69663 63095 69709
rect 63163 69663 63209 69709
rect 63277 69663 63323 69709
rect 63391 69663 63437 69709
rect 63505 69663 63551 69709
rect 63619 69663 63665 69709
rect 63733 69663 63779 69709
rect 63847 69663 63893 69709
rect 63961 69663 64007 69709
rect 64075 69663 64121 69709
rect 64189 69663 64235 69709
rect 64303 69663 64349 69709
rect 64417 69663 64463 69709
rect 64531 69663 64577 69709
rect 64645 69663 64691 69709
rect 64759 69663 64805 69709
rect 64873 69663 64919 69709
rect 64987 69663 65033 69709
rect 65101 69663 65147 69709
rect 65215 69663 65261 69709
rect 65329 69663 65375 69709
rect 65443 69663 65489 69709
rect 65557 69663 65603 69709
rect 65671 69663 65717 69709
rect 65785 69663 65831 69709
rect 65899 69663 65945 69709
rect 66013 69663 66059 69709
rect 66127 69663 66173 69709
rect 66241 69663 66287 69709
rect 66355 69663 66401 69709
rect 66469 69663 66515 69709
rect 66583 69663 66629 69709
rect 66697 69663 66743 69709
rect 66811 69663 66857 69709
rect 66925 69663 66971 69709
rect 67039 69663 67085 69709
rect 67153 69663 67199 69709
rect 67267 69663 67313 69709
rect 67381 69663 67427 69709
rect 67495 69663 67541 69709
rect 67609 69663 67655 69709
rect 67723 69663 67769 69709
rect 67837 69663 67883 69709
rect 67951 69663 67997 69709
rect 68065 69663 68111 69709
rect 68179 69663 68225 69709
rect 68293 69663 68339 69709
rect 68407 69663 68453 69709
rect 68521 69663 68567 69709
rect 68635 69663 68681 69709
rect 68749 69663 68795 69709
rect 68863 69663 68909 69709
rect 68977 69663 69023 69709
rect 69091 69663 69137 69709
rect 69205 69663 69251 69709
rect 69319 69663 69365 69709
rect 69433 69663 69479 69709
rect 60199 69549 60245 69595
rect 60313 69549 60359 69595
rect 60427 69549 60473 69595
rect 60541 69549 60587 69595
rect 60655 69549 60701 69595
rect 60769 69549 60815 69595
rect 60883 69549 60929 69595
rect 60997 69549 61043 69595
rect 61111 69549 61157 69595
rect 61225 69549 61271 69595
rect 61339 69549 61385 69595
rect 61453 69549 61499 69595
rect 61567 69549 61613 69595
rect 61681 69549 61727 69595
rect 61795 69549 61841 69595
rect 61909 69549 61955 69595
rect 62023 69549 62069 69595
rect 62137 69549 62183 69595
rect 62251 69549 62297 69595
rect 62365 69549 62411 69595
rect 62479 69549 62525 69595
rect 62593 69549 62639 69595
rect 62707 69549 62753 69595
rect 62821 69549 62867 69595
rect 62935 69549 62981 69595
rect 63049 69549 63095 69595
rect 63163 69549 63209 69595
rect 63277 69549 63323 69595
rect 63391 69549 63437 69595
rect 63505 69549 63551 69595
rect 63619 69549 63665 69595
rect 63733 69549 63779 69595
rect 63847 69549 63893 69595
rect 63961 69549 64007 69595
rect 64075 69549 64121 69595
rect 64189 69549 64235 69595
rect 64303 69549 64349 69595
rect 64417 69549 64463 69595
rect 64531 69549 64577 69595
rect 64645 69549 64691 69595
rect 64759 69549 64805 69595
rect 64873 69549 64919 69595
rect 64987 69549 65033 69595
rect 65101 69549 65147 69595
rect 65215 69549 65261 69595
rect 65329 69549 65375 69595
rect 65443 69549 65489 69595
rect 65557 69549 65603 69595
rect 65671 69549 65717 69595
rect 65785 69549 65831 69595
rect 65899 69549 65945 69595
rect 66013 69549 66059 69595
rect 66127 69549 66173 69595
rect 66241 69549 66287 69595
rect 66355 69549 66401 69595
rect 66469 69549 66515 69595
rect 66583 69549 66629 69595
rect 66697 69549 66743 69595
rect 66811 69549 66857 69595
rect 66925 69549 66971 69595
rect 67039 69549 67085 69595
rect 67153 69549 67199 69595
rect 67267 69549 67313 69595
rect 67381 69549 67427 69595
rect 67495 69549 67541 69595
rect 67609 69549 67655 69595
rect 67723 69549 67769 69595
rect 67837 69549 67883 69595
rect 67951 69549 67997 69595
rect 68065 69549 68111 69595
rect 68179 69549 68225 69595
rect 68293 69549 68339 69595
rect 68407 69549 68453 69595
rect 68521 69549 68567 69595
rect 68635 69549 68681 69595
rect 68749 69549 68795 69595
rect 68863 69549 68909 69595
rect 68977 69549 69023 69595
rect 69091 69549 69137 69595
rect 69205 69549 69251 69595
rect 69319 69549 69365 69595
rect 69433 69549 69479 69595
rect 60199 69435 60245 69481
rect 60313 69435 60359 69481
rect 60427 69435 60473 69481
rect 60541 69435 60587 69481
rect 60655 69435 60701 69481
rect 60769 69435 60815 69481
rect 60883 69435 60929 69481
rect 60997 69435 61043 69481
rect 61111 69435 61157 69481
rect 61225 69435 61271 69481
rect 61339 69435 61385 69481
rect 61453 69435 61499 69481
rect 61567 69435 61613 69481
rect 61681 69435 61727 69481
rect 61795 69435 61841 69481
rect 61909 69435 61955 69481
rect 62023 69435 62069 69481
rect 62137 69435 62183 69481
rect 62251 69435 62297 69481
rect 62365 69435 62411 69481
rect 62479 69435 62525 69481
rect 62593 69435 62639 69481
rect 62707 69435 62753 69481
rect 62821 69435 62867 69481
rect 62935 69435 62981 69481
rect 63049 69435 63095 69481
rect 63163 69435 63209 69481
rect 63277 69435 63323 69481
rect 63391 69435 63437 69481
rect 63505 69435 63551 69481
rect 63619 69435 63665 69481
rect 63733 69435 63779 69481
rect 63847 69435 63893 69481
rect 63961 69435 64007 69481
rect 64075 69435 64121 69481
rect 64189 69435 64235 69481
rect 64303 69435 64349 69481
rect 64417 69435 64463 69481
rect 64531 69435 64577 69481
rect 64645 69435 64691 69481
rect 64759 69435 64805 69481
rect 64873 69435 64919 69481
rect 64987 69435 65033 69481
rect 65101 69435 65147 69481
rect 65215 69435 65261 69481
rect 65329 69435 65375 69481
rect 65443 69435 65489 69481
rect 65557 69435 65603 69481
rect 65671 69435 65717 69481
rect 65785 69435 65831 69481
rect 65899 69435 65945 69481
rect 66013 69435 66059 69481
rect 66127 69435 66173 69481
rect 66241 69435 66287 69481
rect 66355 69435 66401 69481
rect 66469 69435 66515 69481
rect 66583 69435 66629 69481
rect 66697 69435 66743 69481
rect 66811 69435 66857 69481
rect 66925 69435 66971 69481
rect 67039 69435 67085 69481
rect 67153 69435 67199 69481
rect 67267 69435 67313 69481
rect 67381 69435 67427 69481
rect 67495 69435 67541 69481
rect 67609 69435 67655 69481
rect 67723 69435 67769 69481
rect 67837 69435 67883 69481
rect 67951 69435 67997 69481
rect 68065 69435 68111 69481
rect 68179 69435 68225 69481
rect 68293 69435 68339 69481
rect 68407 69435 68453 69481
rect 68521 69435 68567 69481
rect 68635 69435 68681 69481
rect 68749 69435 68795 69481
rect 68863 69435 68909 69481
rect 68977 69435 69023 69481
rect 69091 69435 69137 69481
rect 69205 69435 69251 69481
rect 69319 69435 69365 69481
rect 69433 69435 69479 69481
rect 60199 69321 60245 69367
rect 60313 69321 60359 69367
rect 60427 69321 60473 69367
rect 60541 69321 60587 69367
rect 60655 69321 60701 69367
rect 60769 69321 60815 69367
rect 60883 69321 60929 69367
rect 60997 69321 61043 69367
rect 61111 69321 61157 69367
rect 61225 69321 61271 69367
rect 61339 69321 61385 69367
rect 61453 69321 61499 69367
rect 61567 69321 61613 69367
rect 61681 69321 61727 69367
rect 61795 69321 61841 69367
rect 61909 69321 61955 69367
rect 62023 69321 62069 69367
rect 62137 69321 62183 69367
rect 62251 69321 62297 69367
rect 62365 69321 62411 69367
rect 62479 69321 62525 69367
rect 62593 69321 62639 69367
rect 62707 69321 62753 69367
rect 62821 69321 62867 69367
rect 62935 69321 62981 69367
rect 63049 69321 63095 69367
rect 63163 69321 63209 69367
rect 63277 69321 63323 69367
rect 63391 69321 63437 69367
rect 63505 69321 63551 69367
rect 63619 69321 63665 69367
rect 63733 69321 63779 69367
rect 63847 69321 63893 69367
rect 63961 69321 64007 69367
rect 64075 69321 64121 69367
rect 64189 69321 64235 69367
rect 64303 69321 64349 69367
rect 64417 69321 64463 69367
rect 64531 69321 64577 69367
rect 64645 69321 64691 69367
rect 64759 69321 64805 69367
rect 64873 69321 64919 69367
rect 64987 69321 65033 69367
rect 65101 69321 65147 69367
rect 65215 69321 65261 69367
rect 65329 69321 65375 69367
rect 65443 69321 65489 69367
rect 65557 69321 65603 69367
rect 65671 69321 65717 69367
rect 65785 69321 65831 69367
rect 65899 69321 65945 69367
rect 66013 69321 66059 69367
rect 66127 69321 66173 69367
rect 66241 69321 66287 69367
rect 66355 69321 66401 69367
rect 66469 69321 66515 69367
rect 66583 69321 66629 69367
rect 66697 69321 66743 69367
rect 66811 69321 66857 69367
rect 66925 69321 66971 69367
rect 67039 69321 67085 69367
rect 67153 69321 67199 69367
rect 67267 69321 67313 69367
rect 67381 69321 67427 69367
rect 67495 69321 67541 69367
rect 67609 69321 67655 69367
rect 67723 69321 67769 69367
rect 67837 69321 67883 69367
rect 67951 69321 67997 69367
rect 68065 69321 68111 69367
rect 68179 69321 68225 69367
rect 68293 69321 68339 69367
rect 68407 69321 68453 69367
rect 68521 69321 68567 69367
rect 68635 69321 68681 69367
rect 68749 69321 68795 69367
rect 68863 69321 68909 69367
rect 68977 69321 69023 69367
rect 69091 69321 69137 69367
rect 69205 69321 69251 69367
rect 69319 69321 69365 69367
rect 69433 69321 69479 69367
rect 60199 69207 60245 69253
rect 60313 69207 60359 69253
rect 60427 69207 60473 69253
rect 60541 69207 60587 69253
rect 60655 69207 60701 69253
rect 60769 69207 60815 69253
rect 60883 69207 60929 69253
rect 60997 69207 61043 69253
rect 61111 69207 61157 69253
rect 61225 69207 61271 69253
rect 61339 69207 61385 69253
rect 61453 69207 61499 69253
rect 61567 69207 61613 69253
rect 61681 69207 61727 69253
rect 61795 69207 61841 69253
rect 61909 69207 61955 69253
rect 62023 69207 62069 69253
rect 62137 69207 62183 69253
rect 62251 69207 62297 69253
rect 62365 69207 62411 69253
rect 62479 69207 62525 69253
rect 62593 69207 62639 69253
rect 62707 69207 62753 69253
rect 62821 69207 62867 69253
rect 62935 69207 62981 69253
rect 63049 69207 63095 69253
rect 63163 69207 63209 69253
rect 63277 69207 63323 69253
rect 63391 69207 63437 69253
rect 63505 69207 63551 69253
rect 63619 69207 63665 69253
rect 63733 69207 63779 69253
rect 63847 69207 63893 69253
rect 63961 69207 64007 69253
rect 64075 69207 64121 69253
rect 64189 69207 64235 69253
rect 64303 69207 64349 69253
rect 64417 69207 64463 69253
rect 64531 69207 64577 69253
rect 64645 69207 64691 69253
rect 64759 69207 64805 69253
rect 64873 69207 64919 69253
rect 64987 69207 65033 69253
rect 65101 69207 65147 69253
rect 65215 69207 65261 69253
rect 65329 69207 65375 69253
rect 65443 69207 65489 69253
rect 65557 69207 65603 69253
rect 65671 69207 65717 69253
rect 65785 69207 65831 69253
rect 65899 69207 65945 69253
rect 66013 69207 66059 69253
rect 66127 69207 66173 69253
rect 66241 69207 66287 69253
rect 66355 69207 66401 69253
rect 66469 69207 66515 69253
rect 66583 69207 66629 69253
rect 66697 69207 66743 69253
rect 66811 69207 66857 69253
rect 66925 69207 66971 69253
rect 67039 69207 67085 69253
rect 67153 69207 67199 69253
rect 67267 69207 67313 69253
rect 67381 69207 67427 69253
rect 67495 69207 67541 69253
rect 67609 69207 67655 69253
rect 67723 69207 67769 69253
rect 67837 69207 67883 69253
rect 67951 69207 67997 69253
rect 68065 69207 68111 69253
rect 68179 69207 68225 69253
rect 68293 69207 68339 69253
rect 68407 69207 68453 69253
rect 68521 69207 68567 69253
rect 68635 69207 68681 69253
rect 68749 69207 68795 69253
rect 68863 69207 68909 69253
rect 68977 69207 69023 69253
rect 69091 69207 69137 69253
rect 69205 69207 69251 69253
rect 69319 69207 69365 69253
rect 69433 69207 69479 69253
rect 60199 69093 60245 69139
rect 60313 69093 60359 69139
rect 60427 69093 60473 69139
rect 60541 69093 60587 69139
rect 60655 69093 60701 69139
rect 60769 69093 60815 69139
rect 60883 69093 60929 69139
rect 60997 69093 61043 69139
rect 61111 69093 61157 69139
rect 61225 69093 61271 69139
rect 61339 69093 61385 69139
rect 61453 69093 61499 69139
rect 61567 69093 61613 69139
rect 61681 69093 61727 69139
rect 61795 69093 61841 69139
rect 61909 69093 61955 69139
rect 62023 69093 62069 69139
rect 62137 69093 62183 69139
rect 62251 69093 62297 69139
rect 62365 69093 62411 69139
rect 62479 69093 62525 69139
rect 62593 69093 62639 69139
rect 62707 69093 62753 69139
rect 62821 69093 62867 69139
rect 62935 69093 62981 69139
rect 63049 69093 63095 69139
rect 63163 69093 63209 69139
rect 63277 69093 63323 69139
rect 63391 69093 63437 69139
rect 63505 69093 63551 69139
rect 63619 69093 63665 69139
rect 63733 69093 63779 69139
rect 63847 69093 63893 69139
rect 63961 69093 64007 69139
rect 64075 69093 64121 69139
rect 64189 69093 64235 69139
rect 64303 69093 64349 69139
rect 64417 69093 64463 69139
rect 64531 69093 64577 69139
rect 64645 69093 64691 69139
rect 64759 69093 64805 69139
rect 64873 69093 64919 69139
rect 64987 69093 65033 69139
rect 65101 69093 65147 69139
rect 65215 69093 65261 69139
rect 65329 69093 65375 69139
rect 65443 69093 65489 69139
rect 65557 69093 65603 69139
rect 65671 69093 65717 69139
rect 65785 69093 65831 69139
rect 65899 69093 65945 69139
rect 66013 69093 66059 69139
rect 66127 69093 66173 69139
rect 66241 69093 66287 69139
rect 66355 69093 66401 69139
rect 66469 69093 66515 69139
rect 66583 69093 66629 69139
rect 66697 69093 66743 69139
rect 66811 69093 66857 69139
rect 66925 69093 66971 69139
rect 67039 69093 67085 69139
rect 67153 69093 67199 69139
rect 67267 69093 67313 69139
rect 67381 69093 67427 69139
rect 67495 69093 67541 69139
rect 67609 69093 67655 69139
rect 67723 69093 67769 69139
rect 67837 69093 67883 69139
rect 67951 69093 67997 69139
rect 68065 69093 68111 69139
rect 68179 69093 68225 69139
rect 68293 69093 68339 69139
rect 68407 69093 68453 69139
rect 68521 69093 68567 69139
rect 68635 69093 68681 69139
rect 68749 69093 68795 69139
rect 68863 69093 68909 69139
rect 68977 69093 69023 69139
rect 69091 69093 69137 69139
rect 69205 69093 69251 69139
rect 69319 69093 69365 69139
rect 69433 69093 69479 69139
rect 60199 68979 60245 69025
rect 60313 68979 60359 69025
rect 60427 68979 60473 69025
rect 60541 68979 60587 69025
rect 60655 68979 60701 69025
rect 60769 68979 60815 69025
rect 60883 68979 60929 69025
rect 60997 68979 61043 69025
rect 61111 68979 61157 69025
rect 61225 68979 61271 69025
rect 61339 68979 61385 69025
rect 61453 68979 61499 69025
rect 61567 68979 61613 69025
rect 61681 68979 61727 69025
rect 61795 68979 61841 69025
rect 61909 68979 61955 69025
rect 62023 68979 62069 69025
rect 62137 68979 62183 69025
rect 62251 68979 62297 69025
rect 62365 68979 62411 69025
rect 62479 68979 62525 69025
rect 62593 68979 62639 69025
rect 62707 68979 62753 69025
rect 62821 68979 62867 69025
rect 62935 68979 62981 69025
rect 63049 68979 63095 69025
rect 63163 68979 63209 69025
rect 63277 68979 63323 69025
rect 63391 68979 63437 69025
rect 63505 68979 63551 69025
rect 63619 68979 63665 69025
rect 63733 68979 63779 69025
rect 63847 68979 63893 69025
rect 63961 68979 64007 69025
rect 64075 68979 64121 69025
rect 64189 68979 64235 69025
rect 64303 68979 64349 69025
rect 64417 68979 64463 69025
rect 64531 68979 64577 69025
rect 64645 68979 64691 69025
rect 64759 68979 64805 69025
rect 64873 68979 64919 69025
rect 64987 68979 65033 69025
rect 65101 68979 65147 69025
rect 65215 68979 65261 69025
rect 65329 68979 65375 69025
rect 65443 68979 65489 69025
rect 65557 68979 65603 69025
rect 65671 68979 65717 69025
rect 65785 68979 65831 69025
rect 65899 68979 65945 69025
rect 66013 68979 66059 69025
rect 66127 68979 66173 69025
rect 66241 68979 66287 69025
rect 66355 68979 66401 69025
rect 66469 68979 66515 69025
rect 66583 68979 66629 69025
rect 66697 68979 66743 69025
rect 66811 68979 66857 69025
rect 66925 68979 66971 69025
rect 67039 68979 67085 69025
rect 67153 68979 67199 69025
rect 67267 68979 67313 69025
rect 67381 68979 67427 69025
rect 67495 68979 67541 69025
rect 67609 68979 67655 69025
rect 67723 68979 67769 69025
rect 67837 68979 67883 69025
rect 67951 68979 67997 69025
rect 68065 68979 68111 69025
rect 68179 68979 68225 69025
rect 68293 68979 68339 69025
rect 68407 68979 68453 69025
rect 68521 68979 68567 69025
rect 68635 68979 68681 69025
rect 68749 68979 68795 69025
rect 68863 68979 68909 69025
rect 68977 68979 69023 69025
rect 69091 68979 69137 69025
rect 69205 68979 69251 69025
rect 69319 68979 69365 69025
rect 69433 68979 69479 69025
<< metal1 >>
rect 60188 70507 69490 70518
rect 60188 70461 60199 70507
rect 60245 70461 60313 70507
rect 60359 70461 60427 70507
rect 60473 70461 60541 70507
rect 60587 70461 60655 70507
rect 60701 70461 60769 70507
rect 60815 70461 60883 70507
rect 60929 70461 60997 70507
rect 61043 70461 61111 70507
rect 61157 70461 61225 70507
rect 61271 70461 61339 70507
rect 61385 70461 61453 70507
rect 61499 70461 61567 70507
rect 61613 70461 61681 70507
rect 61727 70461 61795 70507
rect 61841 70461 61909 70507
rect 61955 70461 62023 70507
rect 62069 70461 62137 70507
rect 62183 70461 62251 70507
rect 62297 70461 62365 70507
rect 62411 70461 62479 70507
rect 62525 70461 62593 70507
rect 62639 70461 62707 70507
rect 62753 70461 62821 70507
rect 62867 70461 62935 70507
rect 62981 70461 63049 70507
rect 63095 70461 63163 70507
rect 63209 70461 63277 70507
rect 63323 70461 63391 70507
rect 63437 70461 63505 70507
rect 63551 70461 63619 70507
rect 63665 70461 63733 70507
rect 63779 70461 63847 70507
rect 63893 70461 63961 70507
rect 64007 70461 64075 70507
rect 64121 70461 64189 70507
rect 64235 70461 64303 70507
rect 64349 70461 64417 70507
rect 64463 70461 64531 70507
rect 64577 70461 64645 70507
rect 64691 70461 64759 70507
rect 64805 70461 64873 70507
rect 64919 70461 64987 70507
rect 65033 70461 65101 70507
rect 65147 70461 65215 70507
rect 65261 70461 65329 70507
rect 65375 70461 65443 70507
rect 65489 70461 65557 70507
rect 65603 70461 65671 70507
rect 65717 70461 65785 70507
rect 65831 70461 65899 70507
rect 65945 70461 66013 70507
rect 66059 70461 66127 70507
rect 66173 70461 66241 70507
rect 66287 70461 66355 70507
rect 66401 70461 66469 70507
rect 66515 70461 66583 70507
rect 66629 70461 66697 70507
rect 66743 70461 66811 70507
rect 66857 70461 66925 70507
rect 66971 70461 67039 70507
rect 67085 70461 67153 70507
rect 67199 70461 67267 70507
rect 67313 70461 67381 70507
rect 67427 70461 67495 70507
rect 67541 70461 67609 70507
rect 67655 70461 67723 70507
rect 67769 70461 67837 70507
rect 67883 70461 67951 70507
rect 67997 70461 68065 70507
rect 68111 70461 68179 70507
rect 68225 70461 68293 70507
rect 68339 70461 68407 70507
rect 68453 70461 68521 70507
rect 68567 70461 68635 70507
rect 68681 70461 68749 70507
rect 68795 70461 68863 70507
rect 68909 70461 68977 70507
rect 69023 70461 69091 70507
rect 69137 70461 69205 70507
rect 69251 70461 69319 70507
rect 69365 70461 69433 70507
rect 69479 70461 69490 70507
rect 60188 70393 69490 70461
rect 60188 70347 60199 70393
rect 60245 70347 60313 70393
rect 60359 70347 60427 70393
rect 60473 70347 60541 70393
rect 60587 70347 60655 70393
rect 60701 70347 60769 70393
rect 60815 70347 60883 70393
rect 60929 70347 60997 70393
rect 61043 70347 61111 70393
rect 61157 70347 61225 70393
rect 61271 70347 61339 70393
rect 61385 70347 61453 70393
rect 61499 70347 61567 70393
rect 61613 70347 61681 70393
rect 61727 70347 61795 70393
rect 61841 70347 61909 70393
rect 61955 70347 62023 70393
rect 62069 70347 62137 70393
rect 62183 70347 62251 70393
rect 62297 70347 62365 70393
rect 62411 70347 62479 70393
rect 62525 70347 62593 70393
rect 62639 70347 62707 70393
rect 62753 70347 62821 70393
rect 62867 70347 62935 70393
rect 62981 70347 63049 70393
rect 63095 70347 63163 70393
rect 63209 70347 63277 70393
rect 63323 70347 63391 70393
rect 63437 70347 63505 70393
rect 63551 70347 63619 70393
rect 63665 70347 63733 70393
rect 63779 70347 63847 70393
rect 63893 70347 63961 70393
rect 64007 70347 64075 70393
rect 64121 70347 64189 70393
rect 64235 70347 64303 70393
rect 64349 70347 64417 70393
rect 64463 70347 64531 70393
rect 64577 70347 64645 70393
rect 64691 70347 64759 70393
rect 64805 70347 64873 70393
rect 64919 70347 64987 70393
rect 65033 70347 65101 70393
rect 65147 70347 65215 70393
rect 65261 70347 65329 70393
rect 65375 70347 65443 70393
rect 65489 70347 65557 70393
rect 65603 70347 65671 70393
rect 65717 70347 65785 70393
rect 65831 70347 65899 70393
rect 65945 70347 66013 70393
rect 66059 70347 66127 70393
rect 66173 70347 66241 70393
rect 66287 70347 66355 70393
rect 66401 70347 66469 70393
rect 66515 70347 66583 70393
rect 66629 70347 66697 70393
rect 66743 70347 66811 70393
rect 66857 70347 66925 70393
rect 66971 70347 67039 70393
rect 67085 70347 67153 70393
rect 67199 70347 67267 70393
rect 67313 70347 67381 70393
rect 67427 70347 67495 70393
rect 67541 70347 67609 70393
rect 67655 70347 67723 70393
rect 67769 70347 67837 70393
rect 67883 70347 67951 70393
rect 67997 70347 68065 70393
rect 68111 70347 68179 70393
rect 68225 70347 68293 70393
rect 68339 70347 68407 70393
rect 68453 70347 68521 70393
rect 68567 70347 68635 70393
rect 68681 70347 68749 70393
rect 68795 70347 68863 70393
rect 68909 70347 68977 70393
rect 69023 70347 69091 70393
rect 69137 70347 69205 70393
rect 69251 70347 69319 70393
rect 69365 70347 69433 70393
rect 69479 70347 69490 70393
rect 60188 70279 69490 70347
rect 60188 70233 60199 70279
rect 60245 70233 60313 70279
rect 60359 70233 60427 70279
rect 60473 70233 60541 70279
rect 60587 70233 60655 70279
rect 60701 70233 60769 70279
rect 60815 70233 60883 70279
rect 60929 70233 60997 70279
rect 61043 70233 61111 70279
rect 61157 70233 61225 70279
rect 61271 70233 61339 70279
rect 61385 70233 61453 70279
rect 61499 70233 61567 70279
rect 61613 70233 61681 70279
rect 61727 70233 61795 70279
rect 61841 70233 61909 70279
rect 61955 70233 62023 70279
rect 62069 70233 62137 70279
rect 62183 70233 62251 70279
rect 62297 70233 62365 70279
rect 62411 70233 62479 70279
rect 62525 70233 62593 70279
rect 62639 70233 62707 70279
rect 62753 70233 62821 70279
rect 62867 70233 62935 70279
rect 62981 70233 63049 70279
rect 63095 70233 63163 70279
rect 63209 70233 63277 70279
rect 63323 70233 63391 70279
rect 63437 70233 63505 70279
rect 63551 70233 63619 70279
rect 63665 70233 63733 70279
rect 63779 70233 63847 70279
rect 63893 70233 63961 70279
rect 64007 70233 64075 70279
rect 64121 70233 64189 70279
rect 64235 70233 64303 70279
rect 64349 70233 64417 70279
rect 64463 70233 64531 70279
rect 64577 70233 64645 70279
rect 64691 70233 64759 70279
rect 64805 70233 64873 70279
rect 64919 70233 64987 70279
rect 65033 70233 65101 70279
rect 65147 70233 65215 70279
rect 65261 70233 65329 70279
rect 65375 70233 65443 70279
rect 65489 70233 65557 70279
rect 65603 70233 65671 70279
rect 65717 70233 65785 70279
rect 65831 70233 65899 70279
rect 65945 70233 66013 70279
rect 66059 70233 66127 70279
rect 66173 70233 66241 70279
rect 66287 70233 66355 70279
rect 66401 70233 66469 70279
rect 66515 70233 66583 70279
rect 66629 70233 66697 70279
rect 66743 70233 66811 70279
rect 66857 70233 66925 70279
rect 66971 70233 67039 70279
rect 67085 70233 67153 70279
rect 67199 70233 67267 70279
rect 67313 70233 67381 70279
rect 67427 70233 67495 70279
rect 67541 70233 67609 70279
rect 67655 70233 67723 70279
rect 67769 70233 67837 70279
rect 67883 70233 67951 70279
rect 67997 70233 68065 70279
rect 68111 70233 68179 70279
rect 68225 70233 68293 70279
rect 68339 70233 68407 70279
rect 68453 70233 68521 70279
rect 68567 70233 68635 70279
rect 68681 70233 68749 70279
rect 68795 70233 68863 70279
rect 68909 70233 68977 70279
rect 69023 70233 69091 70279
rect 69137 70233 69205 70279
rect 69251 70233 69319 70279
rect 69365 70233 69433 70279
rect 69479 70233 69490 70279
rect 60188 70165 69490 70233
rect 60188 70119 60199 70165
rect 60245 70119 60313 70165
rect 60359 70119 60427 70165
rect 60473 70119 60541 70165
rect 60587 70119 60655 70165
rect 60701 70119 60769 70165
rect 60815 70119 60883 70165
rect 60929 70119 60997 70165
rect 61043 70119 61111 70165
rect 61157 70119 61225 70165
rect 61271 70119 61339 70165
rect 61385 70119 61453 70165
rect 61499 70119 61567 70165
rect 61613 70119 61681 70165
rect 61727 70119 61795 70165
rect 61841 70119 61909 70165
rect 61955 70119 62023 70165
rect 62069 70119 62137 70165
rect 62183 70119 62251 70165
rect 62297 70119 62365 70165
rect 62411 70119 62479 70165
rect 62525 70119 62593 70165
rect 62639 70119 62707 70165
rect 62753 70119 62821 70165
rect 62867 70119 62935 70165
rect 62981 70119 63049 70165
rect 63095 70119 63163 70165
rect 63209 70119 63277 70165
rect 63323 70119 63391 70165
rect 63437 70119 63505 70165
rect 63551 70119 63619 70165
rect 63665 70119 63733 70165
rect 63779 70119 63847 70165
rect 63893 70119 63961 70165
rect 64007 70119 64075 70165
rect 64121 70119 64189 70165
rect 64235 70119 64303 70165
rect 64349 70119 64417 70165
rect 64463 70119 64531 70165
rect 64577 70119 64645 70165
rect 64691 70119 64759 70165
rect 64805 70119 64873 70165
rect 64919 70119 64987 70165
rect 65033 70119 65101 70165
rect 65147 70119 65215 70165
rect 65261 70119 65329 70165
rect 65375 70119 65443 70165
rect 65489 70119 65557 70165
rect 65603 70119 65671 70165
rect 65717 70119 65785 70165
rect 65831 70119 65899 70165
rect 65945 70119 66013 70165
rect 66059 70119 66127 70165
rect 66173 70119 66241 70165
rect 66287 70119 66355 70165
rect 66401 70119 66469 70165
rect 66515 70119 66583 70165
rect 66629 70119 66697 70165
rect 66743 70119 66811 70165
rect 66857 70119 66925 70165
rect 66971 70119 67039 70165
rect 67085 70119 67153 70165
rect 67199 70119 67267 70165
rect 67313 70119 67381 70165
rect 67427 70119 67495 70165
rect 67541 70119 67609 70165
rect 67655 70119 67723 70165
rect 67769 70119 67837 70165
rect 67883 70119 67951 70165
rect 67997 70119 68065 70165
rect 68111 70119 68179 70165
rect 68225 70119 68293 70165
rect 68339 70119 68407 70165
rect 68453 70119 68521 70165
rect 68567 70119 68635 70165
rect 68681 70119 68749 70165
rect 68795 70119 68863 70165
rect 68909 70119 68977 70165
rect 69023 70119 69091 70165
rect 69137 70119 69205 70165
rect 69251 70119 69319 70165
rect 69365 70119 69433 70165
rect 69479 70119 69490 70165
rect 60188 70051 69490 70119
rect 60188 70005 60199 70051
rect 60245 70005 60313 70051
rect 60359 70005 60427 70051
rect 60473 70005 60541 70051
rect 60587 70005 60655 70051
rect 60701 70005 60769 70051
rect 60815 70005 60883 70051
rect 60929 70005 60997 70051
rect 61043 70005 61111 70051
rect 61157 70005 61225 70051
rect 61271 70005 61339 70051
rect 61385 70005 61453 70051
rect 61499 70005 61567 70051
rect 61613 70005 61681 70051
rect 61727 70005 61795 70051
rect 61841 70005 61909 70051
rect 61955 70005 62023 70051
rect 62069 70005 62137 70051
rect 62183 70005 62251 70051
rect 62297 70005 62365 70051
rect 62411 70005 62479 70051
rect 62525 70005 62593 70051
rect 62639 70005 62707 70051
rect 62753 70005 62821 70051
rect 62867 70005 62935 70051
rect 62981 70005 63049 70051
rect 63095 70005 63163 70051
rect 63209 70005 63277 70051
rect 63323 70005 63391 70051
rect 63437 70005 63505 70051
rect 63551 70005 63619 70051
rect 63665 70005 63733 70051
rect 63779 70005 63847 70051
rect 63893 70005 63961 70051
rect 64007 70005 64075 70051
rect 64121 70005 64189 70051
rect 64235 70005 64303 70051
rect 64349 70005 64417 70051
rect 64463 70005 64531 70051
rect 64577 70005 64645 70051
rect 64691 70005 64759 70051
rect 64805 70005 64873 70051
rect 64919 70005 64987 70051
rect 65033 70005 65101 70051
rect 65147 70005 65215 70051
rect 65261 70005 65329 70051
rect 65375 70005 65443 70051
rect 65489 70005 65557 70051
rect 65603 70005 65671 70051
rect 65717 70005 65785 70051
rect 65831 70005 65899 70051
rect 65945 70005 66013 70051
rect 66059 70005 66127 70051
rect 66173 70005 66241 70051
rect 66287 70005 66355 70051
rect 66401 70005 66469 70051
rect 66515 70005 66583 70051
rect 66629 70005 66697 70051
rect 66743 70005 66811 70051
rect 66857 70005 66925 70051
rect 66971 70005 67039 70051
rect 67085 70005 67153 70051
rect 67199 70005 67267 70051
rect 67313 70005 67381 70051
rect 67427 70005 67495 70051
rect 67541 70005 67609 70051
rect 67655 70005 67723 70051
rect 67769 70005 67837 70051
rect 67883 70005 67951 70051
rect 67997 70005 68065 70051
rect 68111 70005 68179 70051
rect 68225 70005 68293 70051
rect 68339 70005 68407 70051
rect 68453 70005 68521 70051
rect 68567 70005 68635 70051
rect 68681 70005 68749 70051
rect 68795 70005 68863 70051
rect 68909 70005 68977 70051
rect 69023 70005 69091 70051
rect 69137 70005 69205 70051
rect 69251 70005 69319 70051
rect 69365 70005 69433 70051
rect 69479 70005 69490 70051
rect 60188 69937 69490 70005
rect 60188 69891 60199 69937
rect 60245 69891 60313 69937
rect 60359 69891 60427 69937
rect 60473 69891 60541 69937
rect 60587 69891 60655 69937
rect 60701 69891 60769 69937
rect 60815 69891 60883 69937
rect 60929 69891 60997 69937
rect 61043 69891 61111 69937
rect 61157 69891 61225 69937
rect 61271 69891 61339 69937
rect 61385 69891 61453 69937
rect 61499 69891 61567 69937
rect 61613 69891 61681 69937
rect 61727 69891 61795 69937
rect 61841 69891 61909 69937
rect 61955 69891 62023 69937
rect 62069 69891 62137 69937
rect 62183 69891 62251 69937
rect 62297 69891 62365 69937
rect 62411 69891 62479 69937
rect 62525 69891 62593 69937
rect 62639 69891 62707 69937
rect 62753 69891 62821 69937
rect 62867 69891 62935 69937
rect 62981 69891 63049 69937
rect 63095 69891 63163 69937
rect 63209 69891 63277 69937
rect 63323 69891 63391 69937
rect 63437 69891 63505 69937
rect 63551 69891 63619 69937
rect 63665 69891 63733 69937
rect 63779 69891 63847 69937
rect 63893 69891 63961 69937
rect 64007 69891 64075 69937
rect 64121 69891 64189 69937
rect 64235 69891 64303 69937
rect 64349 69891 64417 69937
rect 64463 69891 64531 69937
rect 64577 69891 64645 69937
rect 64691 69891 64759 69937
rect 64805 69891 64873 69937
rect 64919 69891 64987 69937
rect 65033 69891 65101 69937
rect 65147 69891 65215 69937
rect 65261 69891 65329 69937
rect 65375 69891 65443 69937
rect 65489 69891 65557 69937
rect 65603 69891 65671 69937
rect 65717 69891 65785 69937
rect 65831 69891 65899 69937
rect 65945 69891 66013 69937
rect 66059 69891 66127 69937
rect 66173 69891 66241 69937
rect 66287 69891 66355 69937
rect 66401 69891 66469 69937
rect 66515 69891 66583 69937
rect 66629 69891 66697 69937
rect 66743 69891 66811 69937
rect 66857 69891 66925 69937
rect 66971 69891 67039 69937
rect 67085 69891 67153 69937
rect 67199 69891 67267 69937
rect 67313 69891 67381 69937
rect 67427 69891 67495 69937
rect 67541 69891 67609 69937
rect 67655 69891 67723 69937
rect 67769 69891 67837 69937
rect 67883 69891 67951 69937
rect 67997 69891 68065 69937
rect 68111 69891 68179 69937
rect 68225 69891 68293 69937
rect 68339 69891 68407 69937
rect 68453 69891 68521 69937
rect 68567 69891 68635 69937
rect 68681 69891 68749 69937
rect 68795 69891 68863 69937
rect 68909 69891 68977 69937
rect 69023 69891 69091 69937
rect 69137 69891 69205 69937
rect 69251 69891 69319 69937
rect 69365 69891 69433 69937
rect 69479 69891 69490 69937
rect 60188 69823 69490 69891
rect 60188 69777 60199 69823
rect 60245 69777 60313 69823
rect 60359 69777 60427 69823
rect 60473 69777 60541 69823
rect 60587 69777 60655 69823
rect 60701 69777 60769 69823
rect 60815 69777 60883 69823
rect 60929 69777 60997 69823
rect 61043 69777 61111 69823
rect 61157 69777 61225 69823
rect 61271 69777 61339 69823
rect 61385 69777 61453 69823
rect 61499 69777 61567 69823
rect 61613 69777 61681 69823
rect 61727 69777 61795 69823
rect 61841 69777 61909 69823
rect 61955 69777 62023 69823
rect 62069 69777 62137 69823
rect 62183 69777 62251 69823
rect 62297 69777 62365 69823
rect 62411 69777 62479 69823
rect 62525 69777 62593 69823
rect 62639 69777 62707 69823
rect 62753 69777 62821 69823
rect 62867 69777 62935 69823
rect 62981 69777 63049 69823
rect 63095 69777 63163 69823
rect 63209 69777 63277 69823
rect 63323 69777 63391 69823
rect 63437 69777 63505 69823
rect 63551 69777 63619 69823
rect 63665 69777 63733 69823
rect 63779 69777 63847 69823
rect 63893 69777 63961 69823
rect 64007 69777 64075 69823
rect 64121 69777 64189 69823
rect 64235 69777 64303 69823
rect 64349 69777 64417 69823
rect 64463 69777 64531 69823
rect 64577 69777 64645 69823
rect 64691 69777 64759 69823
rect 64805 69777 64873 69823
rect 64919 69777 64987 69823
rect 65033 69777 65101 69823
rect 65147 69777 65215 69823
rect 65261 69777 65329 69823
rect 65375 69777 65443 69823
rect 65489 69777 65557 69823
rect 65603 69777 65671 69823
rect 65717 69777 65785 69823
rect 65831 69777 65899 69823
rect 65945 69777 66013 69823
rect 66059 69777 66127 69823
rect 66173 69777 66241 69823
rect 66287 69777 66355 69823
rect 66401 69777 66469 69823
rect 66515 69777 66583 69823
rect 66629 69777 66697 69823
rect 66743 69777 66811 69823
rect 66857 69777 66925 69823
rect 66971 69777 67039 69823
rect 67085 69777 67153 69823
rect 67199 69777 67267 69823
rect 67313 69777 67381 69823
rect 67427 69777 67495 69823
rect 67541 69777 67609 69823
rect 67655 69777 67723 69823
rect 67769 69777 67837 69823
rect 67883 69777 67951 69823
rect 67997 69777 68065 69823
rect 68111 69777 68179 69823
rect 68225 69777 68293 69823
rect 68339 69777 68407 69823
rect 68453 69777 68521 69823
rect 68567 69777 68635 69823
rect 68681 69777 68749 69823
rect 68795 69777 68863 69823
rect 68909 69777 68977 69823
rect 69023 69777 69091 69823
rect 69137 69777 69205 69823
rect 69251 69777 69319 69823
rect 69365 69777 69433 69823
rect 69479 69777 69490 69823
rect 60188 69709 69490 69777
rect 60188 69663 60199 69709
rect 60245 69663 60313 69709
rect 60359 69663 60427 69709
rect 60473 69663 60541 69709
rect 60587 69663 60655 69709
rect 60701 69663 60769 69709
rect 60815 69663 60883 69709
rect 60929 69663 60997 69709
rect 61043 69663 61111 69709
rect 61157 69663 61225 69709
rect 61271 69663 61339 69709
rect 61385 69663 61453 69709
rect 61499 69663 61567 69709
rect 61613 69663 61681 69709
rect 61727 69663 61795 69709
rect 61841 69663 61909 69709
rect 61955 69663 62023 69709
rect 62069 69663 62137 69709
rect 62183 69663 62251 69709
rect 62297 69663 62365 69709
rect 62411 69663 62479 69709
rect 62525 69663 62593 69709
rect 62639 69663 62707 69709
rect 62753 69663 62821 69709
rect 62867 69663 62935 69709
rect 62981 69663 63049 69709
rect 63095 69663 63163 69709
rect 63209 69663 63277 69709
rect 63323 69663 63391 69709
rect 63437 69663 63505 69709
rect 63551 69663 63619 69709
rect 63665 69663 63733 69709
rect 63779 69663 63847 69709
rect 63893 69663 63961 69709
rect 64007 69663 64075 69709
rect 64121 69663 64189 69709
rect 64235 69663 64303 69709
rect 64349 69663 64417 69709
rect 64463 69663 64531 69709
rect 64577 69663 64645 69709
rect 64691 69663 64759 69709
rect 64805 69663 64873 69709
rect 64919 69663 64987 69709
rect 65033 69663 65101 69709
rect 65147 69663 65215 69709
rect 65261 69663 65329 69709
rect 65375 69663 65443 69709
rect 65489 69663 65557 69709
rect 65603 69663 65671 69709
rect 65717 69663 65785 69709
rect 65831 69663 65899 69709
rect 65945 69663 66013 69709
rect 66059 69663 66127 69709
rect 66173 69663 66241 69709
rect 66287 69663 66355 69709
rect 66401 69663 66469 69709
rect 66515 69663 66583 69709
rect 66629 69663 66697 69709
rect 66743 69663 66811 69709
rect 66857 69663 66925 69709
rect 66971 69663 67039 69709
rect 67085 69663 67153 69709
rect 67199 69663 67267 69709
rect 67313 69663 67381 69709
rect 67427 69663 67495 69709
rect 67541 69663 67609 69709
rect 67655 69663 67723 69709
rect 67769 69663 67837 69709
rect 67883 69663 67951 69709
rect 67997 69663 68065 69709
rect 68111 69663 68179 69709
rect 68225 69663 68293 69709
rect 68339 69663 68407 69709
rect 68453 69663 68521 69709
rect 68567 69663 68635 69709
rect 68681 69663 68749 69709
rect 68795 69663 68863 69709
rect 68909 69663 68977 69709
rect 69023 69663 69091 69709
rect 69137 69663 69205 69709
rect 69251 69663 69319 69709
rect 69365 69663 69433 69709
rect 69479 69663 69490 69709
rect 60188 69595 69490 69663
rect 60188 69549 60199 69595
rect 60245 69549 60313 69595
rect 60359 69549 60427 69595
rect 60473 69549 60541 69595
rect 60587 69549 60655 69595
rect 60701 69549 60769 69595
rect 60815 69549 60883 69595
rect 60929 69549 60997 69595
rect 61043 69549 61111 69595
rect 61157 69549 61225 69595
rect 61271 69549 61339 69595
rect 61385 69549 61453 69595
rect 61499 69549 61567 69595
rect 61613 69549 61681 69595
rect 61727 69549 61795 69595
rect 61841 69549 61909 69595
rect 61955 69549 62023 69595
rect 62069 69549 62137 69595
rect 62183 69549 62251 69595
rect 62297 69549 62365 69595
rect 62411 69549 62479 69595
rect 62525 69549 62593 69595
rect 62639 69549 62707 69595
rect 62753 69549 62821 69595
rect 62867 69549 62935 69595
rect 62981 69549 63049 69595
rect 63095 69549 63163 69595
rect 63209 69549 63277 69595
rect 63323 69549 63391 69595
rect 63437 69549 63505 69595
rect 63551 69549 63619 69595
rect 63665 69549 63733 69595
rect 63779 69549 63847 69595
rect 63893 69549 63961 69595
rect 64007 69549 64075 69595
rect 64121 69549 64189 69595
rect 64235 69549 64303 69595
rect 64349 69549 64417 69595
rect 64463 69549 64531 69595
rect 64577 69549 64645 69595
rect 64691 69549 64759 69595
rect 64805 69549 64873 69595
rect 64919 69549 64987 69595
rect 65033 69549 65101 69595
rect 65147 69549 65215 69595
rect 65261 69549 65329 69595
rect 65375 69549 65443 69595
rect 65489 69549 65557 69595
rect 65603 69549 65671 69595
rect 65717 69549 65785 69595
rect 65831 69549 65899 69595
rect 65945 69549 66013 69595
rect 66059 69549 66127 69595
rect 66173 69549 66241 69595
rect 66287 69549 66355 69595
rect 66401 69549 66469 69595
rect 66515 69549 66583 69595
rect 66629 69549 66697 69595
rect 66743 69549 66811 69595
rect 66857 69549 66925 69595
rect 66971 69549 67039 69595
rect 67085 69549 67153 69595
rect 67199 69549 67267 69595
rect 67313 69549 67381 69595
rect 67427 69549 67495 69595
rect 67541 69549 67609 69595
rect 67655 69549 67723 69595
rect 67769 69549 67837 69595
rect 67883 69549 67951 69595
rect 67997 69549 68065 69595
rect 68111 69549 68179 69595
rect 68225 69549 68293 69595
rect 68339 69549 68407 69595
rect 68453 69549 68521 69595
rect 68567 69549 68635 69595
rect 68681 69549 68749 69595
rect 68795 69549 68863 69595
rect 68909 69549 68977 69595
rect 69023 69549 69091 69595
rect 69137 69549 69205 69595
rect 69251 69549 69319 69595
rect 69365 69549 69433 69595
rect 69479 69549 69490 69595
rect 60188 69481 69490 69549
rect 60188 69435 60199 69481
rect 60245 69435 60313 69481
rect 60359 69435 60427 69481
rect 60473 69435 60541 69481
rect 60587 69435 60655 69481
rect 60701 69435 60769 69481
rect 60815 69435 60883 69481
rect 60929 69435 60997 69481
rect 61043 69435 61111 69481
rect 61157 69435 61225 69481
rect 61271 69435 61339 69481
rect 61385 69435 61453 69481
rect 61499 69435 61567 69481
rect 61613 69435 61681 69481
rect 61727 69435 61795 69481
rect 61841 69435 61909 69481
rect 61955 69435 62023 69481
rect 62069 69435 62137 69481
rect 62183 69435 62251 69481
rect 62297 69435 62365 69481
rect 62411 69435 62479 69481
rect 62525 69435 62593 69481
rect 62639 69435 62707 69481
rect 62753 69435 62821 69481
rect 62867 69435 62935 69481
rect 62981 69435 63049 69481
rect 63095 69435 63163 69481
rect 63209 69435 63277 69481
rect 63323 69435 63391 69481
rect 63437 69435 63505 69481
rect 63551 69435 63619 69481
rect 63665 69435 63733 69481
rect 63779 69435 63847 69481
rect 63893 69435 63961 69481
rect 64007 69435 64075 69481
rect 64121 69435 64189 69481
rect 64235 69435 64303 69481
rect 64349 69435 64417 69481
rect 64463 69435 64531 69481
rect 64577 69435 64645 69481
rect 64691 69435 64759 69481
rect 64805 69435 64873 69481
rect 64919 69435 64987 69481
rect 65033 69435 65101 69481
rect 65147 69435 65215 69481
rect 65261 69435 65329 69481
rect 65375 69435 65443 69481
rect 65489 69435 65557 69481
rect 65603 69435 65671 69481
rect 65717 69435 65785 69481
rect 65831 69435 65899 69481
rect 65945 69435 66013 69481
rect 66059 69435 66127 69481
rect 66173 69435 66241 69481
rect 66287 69435 66355 69481
rect 66401 69435 66469 69481
rect 66515 69435 66583 69481
rect 66629 69435 66697 69481
rect 66743 69435 66811 69481
rect 66857 69435 66925 69481
rect 66971 69435 67039 69481
rect 67085 69435 67153 69481
rect 67199 69435 67267 69481
rect 67313 69435 67381 69481
rect 67427 69435 67495 69481
rect 67541 69435 67609 69481
rect 67655 69435 67723 69481
rect 67769 69435 67837 69481
rect 67883 69435 67951 69481
rect 67997 69435 68065 69481
rect 68111 69435 68179 69481
rect 68225 69435 68293 69481
rect 68339 69435 68407 69481
rect 68453 69435 68521 69481
rect 68567 69435 68635 69481
rect 68681 69435 68749 69481
rect 68795 69435 68863 69481
rect 68909 69435 68977 69481
rect 69023 69435 69091 69481
rect 69137 69435 69205 69481
rect 69251 69435 69319 69481
rect 69365 69435 69433 69481
rect 69479 69435 69490 69481
rect 60188 69367 69490 69435
rect 60188 69321 60199 69367
rect 60245 69321 60313 69367
rect 60359 69321 60427 69367
rect 60473 69321 60541 69367
rect 60587 69321 60655 69367
rect 60701 69321 60769 69367
rect 60815 69321 60883 69367
rect 60929 69321 60997 69367
rect 61043 69321 61111 69367
rect 61157 69321 61225 69367
rect 61271 69321 61339 69367
rect 61385 69321 61453 69367
rect 61499 69321 61567 69367
rect 61613 69321 61681 69367
rect 61727 69321 61795 69367
rect 61841 69321 61909 69367
rect 61955 69321 62023 69367
rect 62069 69321 62137 69367
rect 62183 69321 62251 69367
rect 62297 69321 62365 69367
rect 62411 69321 62479 69367
rect 62525 69321 62593 69367
rect 62639 69321 62707 69367
rect 62753 69321 62821 69367
rect 62867 69321 62935 69367
rect 62981 69321 63049 69367
rect 63095 69321 63163 69367
rect 63209 69321 63277 69367
rect 63323 69321 63391 69367
rect 63437 69321 63505 69367
rect 63551 69321 63619 69367
rect 63665 69321 63733 69367
rect 63779 69321 63847 69367
rect 63893 69321 63961 69367
rect 64007 69321 64075 69367
rect 64121 69321 64189 69367
rect 64235 69321 64303 69367
rect 64349 69321 64417 69367
rect 64463 69321 64531 69367
rect 64577 69321 64645 69367
rect 64691 69321 64759 69367
rect 64805 69321 64873 69367
rect 64919 69321 64987 69367
rect 65033 69321 65101 69367
rect 65147 69321 65215 69367
rect 65261 69321 65329 69367
rect 65375 69321 65443 69367
rect 65489 69321 65557 69367
rect 65603 69321 65671 69367
rect 65717 69321 65785 69367
rect 65831 69321 65899 69367
rect 65945 69321 66013 69367
rect 66059 69321 66127 69367
rect 66173 69321 66241 69367
rect 66287 69321 66355 69367
rect 66401 69321 66469 69367
rect 66515 69321 66583 69367
rect 66629 69321 66697 69367
rect 66743 69321 66811 69367
rect 66857 69321 66925 69367
rect 66971 69321 67039 69367
rect 67085 69321 67153 69367
rect 67199 69321 67267 69367
rect 67313 69321 67381 69367
rect 67427 69321 67495 69367
rect 67541 69321 67609 69367
rect 67655 69321 67723 69367
rect 67769 69321 67837 69367
rect 67883 69321 67951 69367
rect 67997 69321 68065 69367
rect 68111 69321 68179 69367
rect 68225 69321 68293 69367
rect 68339 69321 68407 69367
rect 68453 69321 68521 69367
rect 68567 69321 68635 69367
rect 68681 69321 68749 69367
rect 68795 69321 68863 69367
rect 68909 69321 68977 69367
rect 69023 69321 69091 69367
rect 69137 69321 69205 69367
rect 69251 69321 69319 69367
rect 69365 69321 69433 69367
rect 69479 69321 69490 69367
rect 60188 69253 69490 69321
rect 60188 69207 60199 69253
rect 60245 69207 60313 69253
rect 60359 69207 60427 69253
rect 60473 69207 60541 69253
rect 60587 69207 60655 69253
rect 60701 69207 60769 69253
rect 60815 69207 60883 69253
rect 60929 69207 60997 69253
rect 61043 69207 61111 69253
rect 61157 69207 61225 69253
rect 61271 69207 61339 69253
rect 61385 69207 61453 69253
rect 61499 69207 61567 69253
rect 61613 69207 61681 69253
rect 61727 69207 61795 69253
rect 61841 69207 61909 69253
rect 61955 69207 62023 69253
rect 62069 69207 62137 69253
rect 62183 69207 62251 69253
rect 62297 69207 62365 69253
rect 62411 69207 62479 69253
rect 62525 69207 62593 69253
rect 62639 69207 62707 69253
rect 62753 69207 62821 69253
rect 62867 69207 62935 69253
rect 62981 69207 63049 69253
rect 63095 69207 63163 69253
rect 63209 69207 63277 69253
rect 63323 69207 63391 69253
rect 63437 69207 63505 69253
rect 63551 69207 63619 69253
rect 63665 69207 63733 69253
rect 63779 69207 63847 69253
rect 63893 69207 63961 69253
rect 64007 69207 64075 69253
rect 64121 69207 64189 69253
rect 64235 69207 64303 69253
rect 64349 69207 64417 69253
rect 64463 69207 64531 69253
rect 64577 69207 64645 69253
rect 64691 69207 64759 69253
rect 64805 69207 64873 69253
rect 64919 69207 64987 69253
rect 65033 69207 65101 69253
rect 65147 69207 65215 69253
rect 65261 69207 65329 69253
rect 65375 69207 65443 69253
rect 65489 69207 65557 69253
rect 65603 69207 65671 69253
rect 65717 69207 65785 69253
rect 65831 69207 65899 69253
rect 65945 69207 66013 69253
rect 66059 69207 66127 69253
rect 66173 69207 66241 69253
rect 66287 69207 66355 69253
rect 66401 69207 66469 69253
rect 66515 69207 66583 69253
rect 66629 69207 66697 69253
rect 66743 69207 66811 69253
rect 66857 69207 66925 69253
rect 66971 69207 67039 69253
rect 67085 69207 67153 69253
rect 67199 69207 67267 69253
rect 67313 69207 67381 69253
rect 67427 69207 67495 69253
rect 67541 69207 67609 69253
rect 67655 69207 67723 69253
rect 67769 69207 67837 69253
rect 67883 69207 67951 69253
rect 67997 69207 68065 69253
rect 68111 69207 68179 69253
rect 68225 69207 68293 69253
rect 68339 69207 68407 69253
rect 68453 69207 68521 69253
rect 68567 69207 68635 69253
rect 68681 69207 68749 69253
rect 68795 69207 68863 69253
rect 68909 69207 68977 69253
rect 69023 69207 69091 69253
rect 69137 69207 69205 69253
rect 69251 69207 69319 69253
rect 69365 69207 69433 69253
rect 69479 69207 69490 69253
rect 60188 69139 69490 69207
rect 60188 69093 60199 69139
rect 60245 69093 60313 69139
rect 60359 69093 60427 69139
rect 60473 69093 60541 69139
rect 60587 69093 60655 69139
rect 60701 69093 60769 69139
rect 60815 69093 60883 69139
rect 60929 69093 60997 69139
rect 61043 69093 61111 69139
rect 61157 69093 61225 69139
rect 61271 69093 61339 69139
rect 61385 69093 61453 69139
rect 61499 69093 61567 69139
rect 61613 69093 61681 69139
rect 61727 69093 61795 69139
rect 61841 69093 61909 69139
rect 61955 69093 62023 69139
rect 62069 69093 62137 69139
rect 62183 69093 62251 69139
rect 62297 69093 62365 69139
rect 62411 69093 62479 69139
rect 62525 69093 62593 69139
rect 62639 69093 62707 69139
rect 62753 69093 62821 69139
rect 62867 69093 62935 69139
rect 62981 69093 63049 69139
rect 63095 69093 63163 69139
rect 63209 69093 63277 69139
rect 63323 69093 63391 69139
rect 63437 69093 63505 69139
rect 63551 69093 63619 69139
rect 63665 69093 63733 69139
rect 63779 69093 63847 69139
rect 63893 69093 63961 69139
rect 64007 69093 64075 69139
rect 64121 69093 64189 69139
rect 64235 69093 64303 69139
rect 64349 69093 64417 69139
rect 64463 69093 64531 69139
rect 64577 69093 64645 69139
rect 64691 69093 64759 69139
rect 64805 69093 64873 69139
rect 64919 69093 64987 69139
rect 65033 69093 65101 69139
rect 65147 69093 65215 69139
rect 65261 69093 65329 69139
rect 65375 69093 65443 69139
rect 65489 69093 65557 69139
rect 65603 69093 65671 69139
rect 65717 69093 65785 69139
rect 65831 69093 65899 69139
rect 65945 69093 66013 69139
rect 66059 69093 66127 69139
rect 66173 69093 66241 69139
rect 66287 69093 66355 69139
rect 66401 69093 66469 69139
rect 66515 69093 66583 69139
rect 66629 69093 66697 69139
rect 66743 69093 66811 69139
rect 66857 69093 66925 69139
rect 66971 69093 67039 69139
rect 67085 69093 67153 69139
rect 67199 69093 67267 69139
rect 67313 69093 67381 69139
rect 67427 69093 67495 69139
rect 67541 69093 67609 69139
rect 67655 69093 67723 69139
rect 67769 69093 67837 69139
rect 67883 69093 67951 69139
rect 67997 69093 68065 69139
rect 68111 69093 68179 69139
rect 68225 69093 68293 69139
rect 68339 69093 68407 69139
rect 68453 69093 68521 69139
rect 68567 69093 68635 69139
rect 68681 69093 68749 69139
rect 68795 69093 68863 69139
rect 68909 69093 68977 69139
rect 69023 69093 69091 69139
rect 69137 69093 69205 69139
rect 69251 69093 69319 69139
rect 69365 69093 69433 69139
rect 69479 69093 69490 69139
rect 60188 69025 69490 69093
rect 60188 68979 60199 69025
rect 60245 68979 60313 69025
rect 60359 68979 60427 69025
rect 60473 68979 60541 69025
rect 60587 68979 60655 69025
rect 60701 68979 60769 69025
rect 60815 68979 60883 69025
rect 60929 68979 60997 69025
rect 61043 68979 61111 69025
rect 61157 68979 61225 69025
rect 61271 68979 61339 69025
rect 61385 68979 61453 69025
rect 61499 68979 61567 69025
rect 61613 68979 61681 69025
rect 61727 68979 61795 69025
rect 61841 68979 61909 69025
rect 61955 68979 62023 69025
rect 62069 68979 62137 69025
rect 62183 68979 62251 69025
rect 62297 68979 62365 69025
rect 62411 68979 62479 69025
rect 62525 68979 62593 69025
rect 62639 68979 62707 69025
rect 62753 68979 62821 69025
rect 62867 68979 62935 69025
rect 62981 68979 63049 69025
rect 63095 68979 63163 69025
rect 63209 68979 63277 69025
rect 63323 68979 63391 69025
rect 63437 68979 63505 69025
rect 63551 68979 63619 69025
rect 63665 68979 63733 69025
rect 63779 68979 63847 69025
rect 63893 68979 63961 69025
rect 64007 68979 64075 69025
rect 64121 68979 64189 69025
rect 64235 68979 64303 69025
rect 64349 68979 64417 69025
rect 64463 68979 64531 69025
rect 64577 68979 64645 69025
rect 64691 68979 64759 69025
rect 64805 68979 64873 69025
rect 64919 68979 64987 69025
rect 65033 68979 65101 69025
rect 65147 68979 65215 69025
rect 65261 68979 65329 69025
rect 65375 68979 65443 69025
rect 65489 68979 65557 69025
rect 65603 68979 65671 69025
rect 65717 68979 65785 69025
rect 65831 68979 65899 69025
rect 65945 68979 66013 69025
rect 66059 68979 66127 69025
rect 66173 68979 66241 69025
rect 66287 68979 66355 69025
rect 66401 68979 66469 69025
rect 66515 68979 66583 69025
rect 66629 68979 66697 69025
rect 66743 68979 66811 69025
rect 66857 68979 66925 69025
rect 66971 68979 67039 69025
rect 67085 68979 67153 69025
rect 67199 68979 67267 69025
rect 67313 68979 67381 69025
rect 67427 68979 67495 69025
rect 67541 68979 67609 69025
rect 67655 68979 67723 69025
rect 67769 68979 67837 69025
rect 67883 68979 67951 69025
rect 67997 68979 68065 69025
rect 68111 68979 68179 69025
rect 68225 68979 68293 69025
rect 68339 68979 68407 69025
rect 68453 68979 68521 69025
rect 68567 68979 68635 69025
rect 68681 68979 68749 69025
rect 68795 68979 68863 69025
rect 68909 68979 68977 69025
rect 69023 68979 69091 69025
rect 69137 68979 69205 69025
rect 69251 68979 69319 69025
rect 69365 68979 69433 69025
rect 69479 68979 69490 69025
rect 60188 68968 69490 68979
<< metal2 >>
rect 41230 69040 41920 69720
rect 39940 67850 40460 68400
rect 67990 40330 68400 40820
rect 69180 40330 69680 40850
use ESD_CLAMP_COR  ESD_CLAMP_COR_0
timestamp 1758744525
transform 1 0 13500 0 1 13500
box 0 0 57389 57390
use moscap_corner  moscap_corner_0
timestamp 1758726819
transform 1 0 59877 0 1 56727
box 32 32 10576 12320
use moscap_corner_1  moscap_corner_1_0
timestamp 1758726819
transform 1 0 10870 0 1 43133
box 4904 32 10576 12320
use moscap_corner  moscap_corner_1
timestamp 1758726819
transform 1 0 45978 0 1 16351
box 32 32 10576 12320
use moscap_corner_2  moscap_corner_2_0
timestamp 1758726819
transform 1 0 25298 0 1 28703
box 32 32 10576 12320
use moscap_corner  moscap_corner_2
timestamp 1758726819
transform 1 0 45978 0 1 28703
box 32 32 10576 12320
use moscap_corner  moscap_corner_3
timestamp 1758726819
transform 1 0 41890 0 1 43133
box 32 32 10576 12320
use moscap_corner_3  moscap_corner_3_0
timestamp 1758726819
transform 1 0 35370 0 1 16351
box 2285 32 10576 12320
use moscap_corner  moscap_corner_4
timestamp 1758726819
transform 1 0 35638 0 1 28703
box 32 32 10576 12320
use moscap_corner  moscap_corner_5
timestamp 1758726819
transform 1 0 31550 0 1 43133
box 32 32 10576 12320
use moscap_corner  moscap_corner_6
timestamp 1758726819
transform 1 0 21210 0 1 43133
box 32 32 10576 12320
use moscap_routing  moscap_routing_0
timestamp 1758726819
transform 1 0 60556 0 1 68904
box -47022 -55377 9837 76
<< labels >>
rlabel metal3 s 18632 70151 18632 70151 4 DVSS
port 1 nsew
rlabel metal2 69420 40560 69420 40560 0 VSS
rlabel metal2 67990 40330 68400 40820 0 VDD
rlabel metal2 41230 69040 41920 69720 0 DVSS
rlabel metal2 39940 67850 40460 68400 0 DVDD
<< end >>
