magic
tech gf180mcuD
magscale 1 10
timestamp 1758725296
<< psubdiff >>
rect 1648 933 1682 1005
rect 1638 -214 1672 -142
rect 1990 -1333 2018 -1261
rect 2020 -2426 2048 -2354
<< nsubdiff >>
rect 1648 217 1682 289
rect 1638 -930 1672 -858
rect 1990 -2049 2018 -1977
rect 2020 -3142 2048 -3070
<< metal1 >>
rect 946 929 2560 1086
rect 946 -57 1194 929
rect 2145 812 2197 825
rect 1324 747 1376 759
rect 1649 700 1805 713
rect 1586 653 1649 699
rect 1910 652 2099 698
rect 1649 636 1805 648
rect 2145 643 2197 656
rect 2288 652 2299 704
rect 2455 652 2467 704
rect 1324 578 1376 591
rect 2636 292 2884 1086
rect 1277 131 2884 292
rect 946 -218 2560 -57
rect 946 -1181 1194 -218
rect 2136 -332 2188 -319
rect 1316 -408 1368 -396
rect 1639 -446 1795 -434
rect 1573 -494 1639 -448
rect 1921 -496 2089 -450
rect 1639 -510 1795 -498
rect 2136 -505 2188 -488
rect 2267 -498 2280 -446
rect 2436 -498 2448 -446
rect 1316 -577 1368 -564
rect 2636 -855 2884 131
rect 1266 -1016 2884 -855
rect 946 -1342 2560 -1181
rect 946 -2269 1194 -1342
rect 1971 -1402 2043 -1394
rect 1909 -1407 2098 -1402
rect 1909 -1494 1980 -1407
rect 1455 -1507 1636 -1500
rect 1455 -1559 1470 -1507
rect 1626 -1559 1636 -1507
rect 1455 -1573 1636 -1559
rect 1971 -1563 1980 -1494
rect 2032 -1494 2098 -1407
rect 2369 -1426 2550 -1416
rect 2369 -1478 2381 -1426
rect 2537 -1478 2550 -1426
rect 2369 -1489 2550 -1478
rect 2032 -1563 2043 -1494
rect 1971 -1579 2043 -1563
rect 2366 -1629 2547 -1619
rect 2366 -1681 2374 -1629
rect 2530 -1681 2547 -1629
rect 2366 -1692 2547 -1681
rect 1455 -1709 1636 -1700
rect 1455 -1761 1470 -1709
rect 1626 -1761 1636 -1709
rect 1455 -1773 1636 -1761
rect 1580 -1856 1763 -1850
rect 1580 -1908 1593 -1856
rect 1749 -1908 1763 -1856
rect 1580 -1918 1763 -1908
rect 2249 -1853 2433 -1847
rect 2249 -1905 2261 -1853
rect 2417 -1905 2433 -1853
rect 2249 -1915 2433 -1905
rect 2636 -1974 2884 -1016
rect 1470 -2135 2884 -1974
rect 946 -2430 2560 -2269
rect 946 -3243 1194 -2430
rect 1842 -2708 1855 -2656
rect 2011 -2708 2025 -2656
rect 2217 -2710 2230 -2658
rect 2386 -2710 2398 -2658
rect 1727 -2825 1779 -2793
rect 1727 -3011 1779 -2981
rect 2122 -2825 2174 -2786
rect 2122 -3011 2174 -2981
rect 2636 -3067 2884 -2135
rect 1470 -3223 2884 -3067
rect 1611 -3284 1663 -3272
rect 2122 -3284 2174 -3272
rect 1663 -3346 2122 -3285
rect 1611 -3452 1663 -3440
rect 2460 -3284 2512 -3272
rect 2174 -3346 2460 -3285
rect 2122 -3452 2174 -3440
rect 2246 -3414 2298 -3402
rect 1493 -3496 1545 -3484
rect 1545 -3549 2246 -3498
rect 2460 -3452 2512 -3440
rect 2246 -3582 2298 -3570
rect 1493 -3664 1545 -3652
<< via1 >>
rect 1324 591 1376 747
rect 1649 648 1805 700
rect 2145 656 2197 812
rect 2299 652 2455 704
rect 1316 -564 1368 -408
rect 1639 -498 1795 -446
rect 2136 -488 2188 -332
rect 2280 -498 2436 -446
rect 1470 -1559 1626 -1507
rect 1980 -1563 2032 -1407
rect 2381 -1478 2537 -1426
rect 2374 -1681 2530 -1629
rect 1470 -1761 1626 -1709
rect 1593 -1908 1749 -1856
rect 2261 -1905 2417 -1853
rect 1855 -2708 2011 -2656
rect 2230 -2710 2386 -2658
rect 1727 -2981 1779 -2825
rect 2122 -2981 2174 -2825
rect 1611 -3440 1663 -3284
rect 2122 -3440 2174 -3284
rect 1493 -3652 1545 -3496
rect 2246 -3570 2298 -3414
rect 2460 -3440 2512 -3284
<< metal2 >>
rect 1678 1017 2905 1073
rect 1320 747 1379 760
rect 1320 591 1324 747
rect 1376 591 1379 747
rect 1678 702 1734 1017
rect 1908 905 2793 961
rect 1636 700 1817 702
rect 1636 648 1649 700
rect 1805 648 1817 700
rect 1636 645 1817 648
rect 1320 582 1379 591
rect 1908 582 1964 905
rect 1320 526 1964 582
rect 2136 825 2199 829
rect 2136 812 2200 825
rect 2136 656 2145 812
rect 2197 656 2200 812
rect 2136 641 2200 656
rect 2286 704 2674 709
rect 2286 652 2299 704
rect 2455 652 2674 704
rect 2286 647 2674 652
rect 2136 -319 2199 641
rect 2133 -332 2199 -319
rect 1313 -408 1372 -396
rect 1313 -564 1316 -408
rect 1368 -564 1372 -408
rect 1313 -578 1372 -564
rect 1624 -446 1807 -443
rect 1624 -498 1639 -446
rect 1795 -498 1807 -446
rect 1624 -502 1807 -498
rect 2133 -488 2136 -332
rect 2188 -488 2199 -332
rect 1313 -625 1369 -578
rect 1117 -681 1369 -625
rect 1117 -3186 1173 -681
rect 1624 -813 1680 -502
rect 2133 -504 2199 -488
rect 2268 -446 2448 -442
rect 2268 -498 2280 -446
rect 2436 -498 2448 -446
rect 2268 -501 2448 -498
rect 1230 -869 1680 -813
rect 1230 -3061 1286 -869
rect 2136 -966 2199 -504
rect 1975 -1029 2199 -966
rect 1975 -1394 2038 -1029
rect 2284 -1123 2340 -501
rect 2126 -1179 2340 -1123
rect 1971 -1407 2043 -1394
rect 1342 -1507 1640 -1500
rect 1342 -1559 1470 -1507
rect 1626 -1559 1640 -1507
rect 1342 -1573 1640 -1559
rect 1971 -1563 1980 -1407
rect 2032 -1563 2043 -1407
rect 1342 -2893 1398 -1573
rect 1971 -1579 2043 -1563
rect 1455 -1709 1636 -1700
rect 1455 -1761 1470 -1709
rect 1626 -1761 1636 -1709
rect 1455 -1773 1636 -1761
rect 1455 -2660 1511 -1773
rect 1723 -1850 1783 -1849
rect 1580 -1856 1783 -1850
rect 1580 -1908 1593 -1856
rect 1749 -1908 1783 -1856
rect 1580 -1918 1783 -1908
rect 1455 -2716 1665 -2660
rect 1342 -2949 1547 -2893
rect 1230 -3117 1404 -3061
rect 1117 -3244 1272 -3186
rect 1348 -3269 1404 -3117
rect 1491 -3496 1547 -2949
rect 1609 -3284 1665 -2716
rect 1723 -2825 1783 -1918
rect 2126 -1853 2182 -1179
rect 2618 -1274 2674 647
rect 2254 -1330 2674 -1274
rect 2254 -1627 2310 -1330
rect 2369 -1426 2673 -1416
rect 2369 -1478 2381 -1426
rect 2537 -1478 2673 -1426
rect 2369 -1489 2673 -1478
rect 2366 -1627 2545 -1619
rect 2254 -1629 2545 -1627
rect 2254 -1681 2374 -1629
rect 2530 -1681 2545 -1629
rect 2254 -1683 2545 -1681
rect 2366 -1692 2545 -1683
rect 2249 -1853 2433 -1847
rect 2126 -1905 2261 -1853
rect 2417 -1905 2433 -1853
rect 2126 -1909 2433 -1905
rect 2126 -1932 2182 -1909
rect 2249 -1915 2433 -1909
rect 1969 -1988 2182 -1932
rect 1969 -2653 2025 -1988
rect 2489 -2178 2545 -1692
rect 1842 -2656 2025 -2653
rect 2244 -2234 2545 -2178
rect 2244 -2655 2300 -2234
rect 2617 -2319 2673 -1489
rect 2459 -2375 2673 -2319
rect 1842 -2708 1855 -2656
rect 2011 -2708 2025 -2656
rect 1842 -2712 2025 -2708
rect 1723 -2981 1727 -2825
rect 1779 -2981 1783 -2825
rect 1723 -3032 1783 -2981
rect 1609 -3440 1611 -3284
rect 1663 -3440 1665 -3284
rect 1969 -3416 2025 -2712
rect 2218 -2658 2398 -2655
rect 2218 -2710 2230 -2658
rect 2386 -2710 2398 -2658
rect 2218 -2715 2398 -2710
rect 2118 -2825 2178 -2810
rect 2118 -2981 2122 -2825
rect 2174 -2981 2178 -2825
rect 2118 -3284 2178 -2981
rect 1609 -3472 1665 -3440
rect 2118 -3440 2122 -3284
rect 2174 -3440 2178 -3284
rect 2118 -3455 2178 -3440
rect 2244 -3414 2300 -2715
rect 2459 -3265 2515 -2375
rect 2737 -2508 2793 905
rect 2594 -2574 2793 -2508
rect 2594 -3251 2650 -2574
rect 2849 -2633 2905 1017
rect 2746 -2697 2905 -2633
rect 2746 -3251 2802 -2697
rect 1491 -3652 1493 -3496
rect 1545 -3652 1547 -3496
rect 2244 -3570 2246 -3414
rect 2298 -3570 2300 -3414
rect 2456 -3284 2516 -3265
rect 2456 -3440 2460 -3284
rect 2512 -3440 2516 -3284
rect 2456 -3455 2516 -3440
rect 2244 -3587 2300 -3570
rect 1491 -3664 1547 -3652
use lv_inv  lv_inv_0
timestamp 1758724778
transform -1 0 18104 0 -1 50671
box 16038 50813 16457 51634
use lv_inv  lv_inv_1
timestamp 1758724778
transform -1 0 18114 0 -1 51818
box 16038 50813 16457 51634
use lv_inv  lv_inv_2
timestamp 1758724778
transform -1 0 18480 0 -1 48459
box 16038 50813 16457 51634
use lv_inv  lv_inv_3
timestamp 1758724778
transform -1 0 18086 0 -1 48459
box 16038 50813 16457 51634
use lv_inv  lv_inv_5
timestamp 1758724778
transform -1 0 17714 0 -1 51818
box 16038 50813 16457 51634
use lv_inv  lv_inv_7
timestamp 1758724778
transform -1 0 17704 0 -1 50671
box 16038 50813 16457 51634
use lv_nand  lv_nand_0
timestamp 1758724778
transform -1 0 19464 0 -1 51807
box 16932 50802 17513 51623
use lv_nand  lv_nand_4
timestamp 1758724778
transform -1 0 19454 0 -1 50660
box 16932 50802 17513 51623
use lv_passgate  lv_passgate_0
timestamp 1758724778
transform 1 0 -13799 0 -1 44483
box 15342 45744 15814 46565
use lv_passgate  lv_passgate_1
timestamp 1758724778
transform -1 0 17807 0 -1 44483
box 15342 45744 15814 46565
<< end >>
