magic
tech gf180mcuB
magscale 1 10
timestamp 1758827725
<< metal4 >>
rect 0 63600 1000 65000
rect 0 49200 1000 50600
use GF_NI_BRK5_0  GF_NI_BRK5_0_0 ..
timestamp 1484609607
transform 1 0 0 0 1 0
box -32 13097 1032 69968
<< labels >>
flabel metal4 s 0 63600 1000 65000 0 FreeSans 1600 0 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 0 49200 1000 50600 0 FreeSans 1600 0 0 0 VSS
port 1 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 1000 70000
string LEFclass PAD SPACER
string LEFsite GF_IO_Site
string LEFsymmetry X Y R90
<< end >>
