magic
tech gf180mcuD
magscale 1 10
timestamp 1758724778
<< nwell >>
rect 18187 54691 19183 55985
<< mvnmos >>
rect 18514 53764 18654 54064
rect 18758 53764 18898 54064
<< mvpmos >>
rect 18514 55332 18654 55632
rect 18758 55332 18898 55632
<< mvndiff >>
rect 18426 54051 18514 54064
rect 18426 54005 18439 54051
rect 18485 54005 18514 54051
rect 18426 53937 18514 54005
rect 18426 53891 18439 53937
rect 18485 53891 18514 53937
rect 18426 53823 18514 53891
rect 18426 53777 18439 53823
rect 18485 53777 18514 53823
rect 18426 53764 18514 53777
rect 18654 54051 18758 54064
rect 18654 54005 18683 54051
rect 18729 54005 18758 54051
rect 18654 53937 18758 54005
rect 18654 53891 18683 53937
rect 18729 53891 18758 53937
rect 18654 53823 18758 53891
rect 18654 53777 18683 53823
rect 18729 53777 18758 53823
rect 18654 53764 18758 53777
rect 18898 54051 18988 54064
rect 18898 54005 18927 54051
rect 18973 54005 18988 54051
rect 18898 53937 18988 54005
rect 18898 53891 18927 53937
rect 18973 53891 18988 53937
rect 18898 53823 18988 53891
rect 18898 53777 18927 53823
rect 18973 53777 18988 53823
rect 18898 53764 18988 53777
<< mvpdiff >>
rect 18426 55619 18514 55632
rect 18426 55573 18439 55619
rect 18485 55573 18514 55619
rect 18426 55514 18514 55573
rect 18426 55468 18439 55514
rect 18485 55468 18514 55514
rect 18426 55409 18514 55468
rect 18426 55363 18439 55409
rect 18485 55363 18514 55409
rect 18426 55332 18514 55363
rect 18654 55619 18758 55632
rect 18654 55573 18683 55619
rect 18729 55573 18758 55619
rect 18654 55514 18758 55573
rect 18654 55468 18683 55514
rect 18729 55468 18758 55514
rect 18654 55409 18758 55468
rect 18654 55363 18683 55409
rect 18729 55363 18758 55409
rect 18654 55332 18758 55363
rect 18898 55619 18988 55632
rect 18898 55573 18927 55619
rect 18973 55573 18988 55619
rect 18898 55514 18988 55573
rect 18898 55468 18927 55514
rect 18973 55468 18988 55514
rect 18898 55409 18988 55468
rect 18898 55363 18927 55409
rect 18973 55363 18988 55409
rect 18898 55332 18988 55363
<< mvndiffc >>
rect 18439 54005 18485 54051
rect 18439 53891 18485 53937
rect 18439 53777 18485 53823
rect 18683 54005 18729 54051
rect 18683 53891 18729 53937
rect 18683 53777 18729 53823
rect 18927 54005 18973 54051
rect 18927 53891 18973 53937
rect 18927 53777 18973 53823
<< mvpdiffc >>
rect 18439 55573 18485 55619
rect 18439 55468 18485 55514
rect 18439 55363 18485 55409
rect 18683 55573 18729 55619
rect 18683 55468 18729 55514
rect 18683 55363 18729 55409
rect 18927 55573 18973 55619
rect 18927 55468 18973 55514
rect 18927 55363 18973 55409
<< psubdiff >>
rect 18264 54324 18354 54346
rect 18264 53432 18286 54324
rect 18332 53500 18354 54324
rect 19061 54418 19151 54440
rect 19061 53500 19083 54418
rect 18332 53478 19083 53500
rect 18332 53432 18416 53478
rect 18989 53432 19083 53478
rect 19129 53432 19151 54418
rect 18264 53410 19151 53432
<< nsubdiff >>
rect 18264 55880 19151 55902
rect 18264 54894 18286 55880
rect 18332 55834 18425 55880
rect 19000 55834 19083 55880
rect 18332 55812 19083 55834
rect 18332 54894 18354 55812
rect 18264 54872 18354 54894
rect 19061 54894 19083 55812
rect 19129 54894 19151 55880
rect 19061 54872 19151 54894
<< psubdiffcont >>
rect 18286 53432 18332 54324
rect 18416 53432 18989 53478
rect 19083 53432 19129 54418
<< nsubdiffcont >>
rect 18286 54894 18332 55880
rect 18425 55834 19000 55880
rect 19083 54894 19129 55880
<< polysilicon >>
rect 18514 55632 18654 55676
rect 18758 55632 18898 55676
rect 18514 55272 18654 55332
rect 18514 55257 18688 55272
rect 18514 55195 18560 55257
rect 18672 55195 18688 55257
rect 18514 55181 18688 55195
rect 18758 55130 18898 55332
rect 18528 55116 18898 55130
rect 18528 55056 18544 55116
rect 18747 55056 18898 55116
rect 18528 55040 18898 55056
rect 18504 54786 18898 54830
rect 18504 54687 18523 54786
rect 18644 54687 18898 54786
rect 18504 54667 18898 54687
rect 18502 54527 18654 54544
rect 18502 54420 18515 54527
rect 18639 54420 18654 54527
rect 18502 54386 18654 54420
rect 18514 54064 18654 54386
rect 18758 54064 18898 54667
rect 18514 53720 18654 53764
rect 18758 53720 18898 53764
<< polycontact >>
rect 18560 55195 18672 55257
rect 18544 55056 18747 55116
rect 18523 54687 18644 54786
rect 18515 54420 18639 54527
<< metal1 >>
rect 18275 55880 19144 55891
rect 18275 54894 18286 55880
rect 18332 55834 18425 55880
rect 19000 55834 19083 55880
rect 18332 55823 19083 55834
rect 18332 54894 18343 55823
rect 18424 55619 18500 55632
rect 18424 55573 18439 55619
rect 18485 55573 18500 55619
rect 18424 55514 18500 55573
rect 18424 55468 18439 55514
rect 18485 55468 18500 55514
rect 18424 55409 18500 55468
rect 18424 55363 18439 55409
rect 18485 55363 18500 55409
rect 18424 55129 18500 55363
rect 18668 55619 18745 55823
rect 18668 55573 18683 55619
rect 18729 55573 18745 55619
rect 18668 55514 18745 55573
rect 18668 55468 18683 55514
rect 18729 55468 18745 55514
rect 18668 55409 18745 55468
rect 18668 55363 18683 55409
rect 18729 55363 18745 55409
rect 18668 55328 18745 55363
rect 18912 55619 18988 55632
rect 18912 55573 18927 55619
rect 18973 55573 18988 55619
rect 18912 55514 18988 55573
rect 18912 55468 18927 55514
rect 18973 55468 18988 55514
rect 18912 55409 18988 55468
rect 18912 55363 18927 55409
rect 18973 55363 18988 55409
rect 18912 55272 18988 55363
rect 18547 55257 18988 55272
rect 18547 55195 18560 55257
rect 18672 55195 18988 55257
rect 18547 55178 18988 55195
rect 18424 55116 18805 55129
rect 18424 55056 18544 55116
rect 18747 55056 18805 55116
rect 18424 55043 18805 55056
rect 18275 54883 18343 54894
rect 18394 54786 18655 54820
rect 18394 54687 18523 54786
rect 18644 54687 18655 54786
rect 18394 54663 18655 54687
rect 18394 54527 18655 54543
rect 18394 54420 18515 54527
rect 18639 54420 18655 54527
rect 18394 54386 18655 54420
rect 18275 54324 18343 54335
rect 18275 53432 18286 54324
rect 18332 53489 18343 54324
rect 18729 54208 18805 55043
rect 18424 54132 18805 54208
rect 18424 54051 18500 54132
rect 18424 54005 18439 54051
rect 18485 54005 18500 54051
rect 18424 53937 18500 54005
rect 18424 53891 18439 53937
rect 18485 53891 18500 53937
rect 18424 53823 18500 53891
rect 18424 53777 18439 53823
rect 18485 53777 18500 53823
rect 18424 53764 18500 53777
rect 18668 54051 18743 54064
rect 18668 54005 18683 54051
rect 18729 54005 18743 54051
rect 18668 53937 18743 54005
rect 18668 53891 18683 53937
rect 18729 53891 18743 53937
rect 18668 53823 18743 53891
rect 18668 53777 18683 53823
rect 18729 53777 18743 53823
rect 18668 53489 18743 53777
rect 18912 54051 18988 55178
rect 19068 54894 19083 55823
rect 19129 54894 19144 55880
rect 19068 54883 19144 54894
rect 19072 54418 19140 54429
rect 19072 54329 19083 54418
rect 18912 54005 18927 54051
rect 18973 54005 18988 54051
rect 18912 53937 18988 54005
rect 18912 53891 18927 53937
rect 18973 53891 18988 53937
rect 18912 53823 18988 53891
rect 18912 53777 18927 53823
rect 18973 53777 18988 53823
rect 18912 53764 18988 53777
rect 19068 53489 19083 54329
rect 18332 53478 19083 53489
rect 18332 53432 18416 53478
rect 18989 53432 19083 53478
rect 19129 54329 19140 54418
rect 19129 53432 19144 54329
rect 18275 53421 19144 53432
<< end >>
