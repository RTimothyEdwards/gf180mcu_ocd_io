magic
tech gf180mcuA
magscale 1 10
timestamp 1758829324
<< metal3 >>
rect 0 68400 2000 69678
rect 0 66800 2000 68200
rect 0 65200 2000 66600
rect 0 63600 2000 65000
rect 0 62000 2000 63400
rect 0 60400 2000 61800
rect 0 58800 2000 60200
rect 0 57200 2000 58600
rect 0 55600 2000 57000
rect 0 54000 2000 55400
rect 0 52400 2000 53800
rect 0 50800 2000 52200
rect 0 49200 2000 50600
rect 0 46000 2000 49000
rect 0 42800 2000 45800
rect 0 41200 2000 42600
rect 0 39600 2000 41000
rect 0 36400 2000 39400
rect 0 33200 2000 36200
rect 0 30000 2000 33000
rect 0 26800 2000 29800
rect 0 25200 2000 26600
rect 0 23600 2000 25000
rect 0 20400 2000 23400
rect 0 17200 2000 20200
rect 0 14000 2000 17000
use GF_NI_FILL10_0  GF_NI_FILL10_0_0 ..
timestamp 1484609607
transform 1 0 0 0 1 0
box -32 13097 2032 69968
<< labels >>
flabel metal3 s 0 63600 2000 65000 0 FreeSans 1600 0 0 0 VSS
port 4 nsew ground bidirectional
flabel metal3 s 0 49200 2000 50600 0 FreeSans 1600 0 0 0 VSS
port 4 nsew ground bidirectional
flabel metal3 s 0 50800 2000 52200 0 FreeSans 1600 0 0 0 VDD
port 3 nsew power bidirectional
flabel metal3 s 0 62000 2000 63400 0 FreeSans 1600 0 0 0 VDD
port 3 nsew power bidirectional
flabel metal3 s 0 17200 2000 20200 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal3 s 0 14000 2000 17000 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal3 s 0 20400 2000 23400 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal3 s 0 25200 2000 26600 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal3 s 0 39600 2000 41000 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal3 s 0 46000 2000 49000 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal3 s 0 57200 2000 58600 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal3 s 0 60400 2000 61800 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal3 s 0 65200 2000 66600 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal3 s 0 68400 2000 69678 0 FreeSans 1600 0 0 0 DVSS
port 2 nsew ground bidirectional
flabel metal3 s 0 30000 2000 33000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal3 s 0 26800 2000 29800 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal3 s 0 23600 2000 25000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal3 s 0 58800 2000 60200 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal3 s 0 55600 2000 57000 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal3 s 0 54000 2000 55400 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal3 s 0 52400 2000 53800 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal3 s 0 42800 2000 45800 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal3 s 0 41200 2000 42600 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal3 s 0 36400 2000 39400 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal3 s 0 33200 2000 36200 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
flabel metal3 s 0 66800 2000 68200 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 2000 70000
string LEFclass PAD SPACER
string LEFsite GF_IO_Site
string LEFsymmetry X Y R90
<< end >>
