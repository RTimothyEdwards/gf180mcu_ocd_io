magic
tech gf180mcuD
magscale 1 10
timestamp 1484609607
<< metal2 >>
rect 220 65000 792 69616
rect 0 63600 1000 65000
rect 220 50600 792 63600
rect 0 49200 1000 50600
rect 220 13622 792 49200
<< metal3 >>
rect 158 64886 854 64896
rect 158 64830 168 64886
rect 224 64830 292 64886
rect 348 64830 416 64886
rect 472 64830 540 64886
rect 596 64830 664 64886
rect 720 64830 788 64886
rect 844 64830 854 64886
rect 158 64762 854 64830
rect 158 64706 168 64762
rect 224 64706 292 64762
rect 348 64706 416 64762
rect 472 64706 540 64762
rect 596 64706 664 64762
rect 720 64706 788 64762
rect 844 64706 854 64762
rect 158 64638 854 64706
rect 158 64582 168 64638
rect 224 64582 292 64638
rect 348 64582 416 64638
rect 472 64582 540 64638
rect 596 64582 664 64638
rect 720 64582 788 64638
rect 844 64582 854 64638
rect 158 64514 854 64582
rect 158 64458 168 64514
rect 224 64458 292 64514
rect 348 64458 416 64514
rect 472 64458 540 64514
rect 596 64458 664 64514
rect 720 64458 788 64514
rect 844 64458 854 64514
rect 158 64390 854 64458
rect 158 64334 168 64390
rect 224 64334 292 64390
rect 348 64334 416 64390
rect 472 64334 540 64390
rect 596 64334 664 64390
rect 720 64334 788 64390
rect 844 64334 854 64390
rect 158 64266 854 64334
rect 158 64210 168 64266
rect 224 64210 292 64266
rect 348 64210 416 64266
rect 472 64210 540 64266
rect 596 64210 664 64266
rect 720 64210 788 64266
rect 844 64210 854 64266
rect 158 64142 854 64210
rect 158 64086 168 64142
rect 224 64086 292 64142
rect 348 64086 416 64142
rect 472 64086 540 64142
rect 596 64086 664 64142
rect 720 64086 788 64142
rect 844 64086 854 64142
rect 158 64018 854 64086
rect 158 63962 168 64018
rect 224 63962 292 64018
rect 348 63962 416 64018
rect 472 63962 540 64018
rect 596 63962 664 64018
rect 720 63962 788 64018
rect 844 63962 854 64018
rect 158 63894 854 63962
rect 158 63838 168 63894
rect 224 63838 292 63894
rect 348 63838 416 63894
rect 472 63838 540 63894
rect 596 63838 664 63894
rect 720 63838 788 63894
rect 844 63838 854 63894
rect 158 63770 854 63838
rect 158 63714 168 63770
rect 224 63714 292 63770
rect 348 63714 416 63770
rect 472 63714 540 63770
rect 596 63714 664 63770
rect 720 63714 788 63770
rect 844 63714 854 63770
rect 158 63704 854 63714
rect 150 50480 846 50490
rect 150 50424 160 50480
rect 216 50424 284 50480
rect 340 50424 408 50480
rect 464 50424 532 50480
rect 588 50424 656 50480
rect 712 50424 780 50480
rect 836 50424 846 50480
rect 150 50356 846 50424
rect 150 50300 160 50356
rect 216 50300 284 50356
rect 340 50300 408 50356
rect 464 50300 532 50356
rect 588 50300 656 50356
rect 712 50300 780 50356
rect 836 50300 846 50356
rect 150 50232 846 50300
rect 150 50176 160 50232
rect 216 50176 284 50232
rect 340 50176 408 50232
rect 464 50176 532 50232
rect 588 50176 656 50232
rect 712 50176 780 50232
rect 836 50176 846 50232
rect 150 50108 846 50176
rect 150 50052 160 50108
rect 216 50052 284 50108
rect 340 50052 408 50108
rect 464 50052 532 50108
rect 588 50052 656 50108
rect 712 50052 780 50108
rect 836 50052 846 50108
rect 150 49984 846 50052
rect 150 49928 160 49984
rect 216 49928 284 49984
rect 340 49928 408 49984
rect 464 49928 532 49984
rect 588 49928 656 49984
rect 712 49928 780 49984
rect 836 49928 846 49984
rect 150 49860 846 49928
rect 150 49804 160 49860
rect 216 49804 284 49860
rect 340 49804 408 49860
rect 464 49804 532 49860
rect 588 49804 656 49860
rect 712 49804 780 49860
rect 836 49804 846 49860
rect 150 49736 846 49804
rect 150 49680 160 49736
rect 216 49680 284 49736
rect 340 49680 408 49736
rect 464 49680 532 49736
rect 588 49680 656 49736
rect 712 49680 780 49736
rect 836 49680 846 49736
rect 150 49612 846 49680
rect 150 49556 160 49612
rect 216 49556 284 49612
rect 340 49556 408 49612
rect 464 49556 532 49612
rect 588 49556 656 49612
rect 712 49556 780 49612
rect 836 49556 846 49612
rect 150 49488 846 49556
rect 150 49432 160 49488
rect 216 49432 284 49488
rect 340 49432 408 49488
rect 464 49432 532 49488
rect 588 49432 656 49488
rect 712 49432 780 49488
rect 836 49432 846 49488
rect 150 49364 846 49432
rect 150 49308 160 49364
rect 216 49308 284 49364
rect 340 49308 408 49364
rect 464 49308 532 49364
rect 588 49308 656 49364
rect 712 49308 780 49364
rect 836 49308 846 49364
rect 150 49298 846 49308
<< via3 >>
rect 168 64830 224 64886
rect 292 64830 348 64886
rect 416 64830 472 64886
rect 540 64830 596 64886
rect 664 64830 720 64886
rect 788 64830 844 64886
rect 168 64706 224 64762
rect 292 64706 348 64762
rect 416 64706 472 64762
rect 540 64706 596 64762
rect 664 64706 720 64762
rect 788 64706 844 64762
rect 168 64582 224 64638
rect 292 64582 348 64638
rect 416 64582 472 64638
rect 540 64582 596 64638
rect 664 64582 720 64638
rect 788 64582 844 64638
rect 168 64458 224 64514
rect 292 64458 348 64514
rect 416 64458 472 64514
rect 540 64458 596 64514
rect 664 64458 720 64514
rect 788 64458 844 64514
rect 168 64334 224 64390
rect 292 64334 348 64390
rect 416 64334 472 64390
rect 540 64334 596 64390
rect 664 64334 720 64390
rect 788 64334 844 64390
rect 168 64210 224 64266
rect 292 64210 348 64266
rect 416 64210 472 64266
rect 540 64210 596 64266
rect 664 64210 720 64266
rect 788 64210 844 64266
rect 168 64086 224 64142
rect 292 64086 348 64142
rect 416 64086 472 64142
rect 540 64086 596 64142
rect 664 64086 720 64142
rect 788 64086 844 64142
rect 168 63962 224 64018
rect 292 63962 348 64018
rect 416 63962 472 64018
rect 540 63962 596 64018
rect 664 63962 720 64018
rect 788 63962 844 64018
rect 168 63838 224 63894
rect 292 63838 348 63894
rect 416 63838 472 63894
rect 540 63838 596 63894
rect 664 63838 720 63894
rect 788 63838 844 63894
rect 168 63714 224 63770
rect 292 63714 348 63770
rect 416 63714 472 63770
rect 540 63714 596 63770
rect 664 63714 720 63770
rect 788 63714 844 63770
rect 160 50424 216 50480
rect 284 50424 340 50480
rect 408 50424 464 50480
rect 532 50424 588 50480
rect 656 50424 712 50480
rect 780 50424 836 50480
rect 160 50300 216 50356
rect 284 50300 340 50356
rect 408 50300 464 50356
rect 532 50300 588 50356
rect 656 50300 712 50356
rect 780 50300 836 50356
rect 160 50176 216 50232
rect 284 50176 340 50232
rect 408 50176 464 50232
rect 532 50176 588 50232
rect 656 50176 712 50232
rect 780 50176 836 50232
rect 160 50052 216 50108
rect 284 50052 340 50108
rect 408 50052 464 50108
rect 532 50052 588 50108
rect 656 50052 712 50108
rect 780 50052 836 50108
rect 160 49928 216 49984
rect 284 49928 340 49984
rect 408 49928 464 49984
rect 532 49928 588 49984
rect 656 49928 712 49984
rect 780 49928 836 49984
rect 160 49804 216 49860
rect 284 49804 340 49860
rect 408 49804 464 49860
rect 532 49804 588 49860
rect 656 49804 712 49860
rect 780 49804 836 49860
rect 160 49680 216 49736
rect 284 49680 340 49736
rect 408 49680 464 49736
rect 532 49680 588 49736
rect 656 49680 712 49736
rect 780 49680 836 49736
rect 160 49556 216 49612
rect 284 49556 340 49612
rect 408 49556 464 49612
rect 532 49556 588 49612
rect 656 49556 712 49612
rect 780 49556 836 49612
rect 160 49432 216 49488
rect 284 49432 340 49488
rect 408 49432 464 49488
rect 532 49432 588 49488
rect 656 49432 712 49488
rect 780 49432 836 49488
rect 160 49308 216 49364
rect 284 49308 340 49364
rect 408 49308 464 49364
rect 532 49308 588 49364
rect 656 49308 712 49364
rect 780 49308 836 49364
<< metal4 >>
rect 0 64886 1000 65000
rect 0 64830 168 64886
rect 224 64830 292 64886
rect 348 64830 416 64886
rect 472 64830 540 64886
rect 596 64830 664 64886
rect 720 64830 788 64886
rect 844 64830 1000 64886
rect 0 64762 1000 64830
rect 0 64706 168 64762
rect 224 64706 292 64762
rect 348 64706 416 64762
rect 472 64706 540 64762
rect 596 64706 664 64762
rect 720 64706 788 64762
rect 844 64706 1000 64762
rect 0 64638 1000 64706
rect 0 64582 168 64638
rect 224 64582 292 64638
rect 348 64582 416 64638
rect 472 64582 540 64638
rect 596 64582 664 64638
rect 720 64582 788 64638
rect 844 64582 1000 64638
rect 0 64514 1000 64582
rect 0 64458 168 64514
rect 224 64458 292 64514
rect 348 64458 416 64514
rect 472 64458 540 64514
rect 596 64458 664 64514
rect 720 64458 788 64514
rect 844 64458 1000 64514
rect 0 64390 1000 64458
rect 0 64334 168 64390
rect 224 64334 292 64390
rect 348 64334 416 64390
rect 472 64334 540 64390
rect 596 64334 664 64390
rect 720 64334 788 64390
rect 844 64334 1000 64390
rect 0 64266 1000 64334
rect 0 64210 168 64266
rect 224 64210 292 64266
rect 348 64210 416 64266
rect 472 64210 540 64266
rect 596 64210 664 64266
rect 720 64210 788 64266
rect 844 64210 1000 64266
rect 0 64142 1000 64210
rect 0 64086 168 64142
rect 224 64086 292 64142
rect 348 64086 416 64142
rect 472 64086 540 64142
rect 596 64086 664 64142
rect 720 64086 788 64142
rect 844 64086 1000 64142
rect 0 64018 1000 64086
rect 0 63962 168 64018
rect 224 63962 292 64018
rect 348 63962 416 64018
rect 472 63962 540 64018
rect 596 63962 664 64018
rect 720 63962 788 64018
rect 844 63962 1000 64018
rect 0 63894 1000 63962
rect 0 63838 168 63894
rect 224 63838 292 63894
rect 348 63838 416 63894
rect 472 63838 540 63894
rect 596 63838 664 63894
rect 720 63838 788 63894
rect 844 63838 1000 63894
rect 0 63770 1000 63838
rect 0 63714 168 63770
rect 224 63714 292 63770
rect 348 63714 416 63770
rect 472 63714 540 63770
rect 596 63714 664 63770
rect 720 63714 788 63770
rect 844 63714 1000 63770
rect 0 63600 1000 63714
rect 0 50480 1000 50600
rect 0 50424 160 50480
rect 216 50424 284 50480
rect 340 50424 408 50480
rect 464 50424 532 50480
rect 588 50424 656 50480
rect 712 50424 780 50480
rect 836 50424 1000 50480
rect 0 50356 1000 50424
rect 0 50300 160 50356
rect 216 50300 284 50356
rect 340 50300 408 50356
rect 464 50300 532 50356
rect 588 50300 656 50356
rect 712 50300 780 50356
rect 836 50300 1000 50356
rect 0 50232 1000 50300
rect 0 50176 160 50232
rect 216 50176 284 50232
rect 340 50176 408 50232
rect 464 50176 532 50232
rect 588 50176 656 50232
rect 712 50176 780 50232
rect 836 50176 1000 50232
rect 0 50108 1000 50176
rect 0 50052 160 50108
rect 216 50052 284 50108
rect 340 50052 408 50108
rect 464 50052 532 50108
rect 588 50052 656 50108
rect 712 50052 780 50108
rect 836 50052 1000 50108
rect 0 49984 1000 50052
rect 0 49928 160 49984
rect 216 49928 284 49984
rect 340 49928 408 49984
rect 464 49928 532 49984
rect 588 49928 656 49984
rect 712 49928 780 49984
rect 836 49928 1000 49984
rect 0 49860 1000 49928
rect 0 49804 160 49860
rect 216 49804 284 49860
rect 340 49804 408 49860
rect 464 49804 532 49860
rect 588 49804 656 49860
rect 712 49804 780 49860
rect 836 49804 1000 49860
rect 0 49736 1000 49804
rect 0 49680 160 49736
rect 216 49680 284 49736
rect 340 49680 408 49736
rect 464 49680 532 49736
rect 588 49680 656 49736
rect 712 49680 780 49736
rect 836 49680 1000 49736
rect 0 49612 1000 49680
rect 0 49556 160 49612
rect 216 49556 284 49612
rect 340 49556 408 49612
rect 464 49556 532 49612
rect 588 49556 656 49612
rect 712 49556 780 49612
rect 836 49556 1000 49612
rect 0 49488 1000 49556
rect 0 49432 160 49488
rect 216 49432 284 49488
rect 340 49432 408 49488
rect 464 49432 532 49488
rect 588 49432 656 49488
rect 712 49432 780 49488
rect 836 49432 1000 49488
rect 0 49364 1000 49432
rect 0 49308 160 49364
rect 216 49308 284 49364
rect 340 49308 408 49364
rect 464 49308 532 49364
rect 588 49308 656 49364
rect 712 49308 780 49364
rect 836 49308 1000 49364
rect 0 49200 1000 49308
use GF_NI_BRK5_1  GF_NI_BRK5_1_0
timestamp 1484609607
transform 1 0 0 0 1 0
box -32 13097 1032 69968
<< labels >>
rlabel metal3 s 498 64258 498 64258 4 VSS
port 1 nsew
rlabel metal3 s 510 50023 510 50023 4 VSS
port 1 nsew
rlabel metal4 s 510 50023 510 50023 4 VSS
port 1 nsew
rlabel metal4 s 498 64258 498 64258 4 VSS
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 1000 70000
<< end >>
