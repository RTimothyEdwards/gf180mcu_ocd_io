* NGSPICE file created from gf180mcu_ocd_io__vdd.ext - technology: gf180mcuD

.subckt x5LM_METAL_RAIL_PAD_60 VSUBS Bondpad_5LM_0/m2_n400_0# 5LM_METAL_RAIL_0/VDD
+ 5LM_METAL_RAIL_0/VSS 5LM_METAL_RAIL_0/DVSS 5LM_METAL_RAIL_0/DVDD
.ends

.subckt comp018green_esd_rc_v5p0 VRC VPLUS VMINUS
X0 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X1 a_353_1149# a_13226_869# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X2 a_353_2269# a_13226_1989# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X3 a_353_3389# a_13226_3109# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X4 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X5 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X6 a_353_2829# a_13226_3109# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X7 a_353_1709# a_13226_1989# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X8 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X9 a_353_1709# a_13226_1429# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X10 a_353_2829# a_13226_2549# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X11 VRC a_13226_3669# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X12 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X13 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X14 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X15 VPLUS a_13226_869# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X16 a_353_1149# a_13226_1429# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X17 a_353_2269# a_13226_2549# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
X18 VRC VMINUS cap_nmos_06v0 c_width=25u c_length=10u
X19 a_353_3389# a_13226_3669# VPLUS ppolyf_u r_width=0.8u r_length=63.855u
.ends

.subckt nmos_clamp_20_50_4_DVDD a_582_632# w_n51_n51# a_1237_1481#
X0 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X1 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X2 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=22p pd=0.10088m as=13p ps=50.52u w=50u l=0.7u
X3 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=22p pd=0.10088m as=13p ps=50.52u w=50u l=0.7u
X4 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X5 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X6 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X7 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X8 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X9 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X10 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X11 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X12 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X13 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X14 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X15 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X16 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X17 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X18 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X19 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X20 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X21 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=22p pd=0.10088m as=13p ps=50.52u w=50u l=0.7u
X22 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X23 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X24 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X25 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X26 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X27 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X28 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X29 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X30 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X31 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X32 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X33 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X34 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X35 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X36 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X37 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X38 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X39 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X40 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X41 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X42 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X43 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X44 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=22p ps=0.10088m w=50u l=0.7u
X45 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X46 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X47 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X48 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X49 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X50 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X51 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=22p ps=0.10088m w=50u l=0.7u
X52 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X53 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X54 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X55 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=22p ps=0.10088m w=50u l=0.7u
X56 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X57 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X58 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X59 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X60 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X61 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X62 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X63 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X64 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X65 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X66 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X67 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X68 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X69 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X70 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=22p pd=0.10088m as=13p ps=50.52u w=50u l=0.7u
X71 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X72 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X73 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X74 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X75 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=22p ps=0.10088m w=50u l=0.7u
X76 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X77 w_n51_n51# a_1237_1481# a_582_632# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X78 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
X79 a_582_632# a_1237_1481# w_n51_n51# a_582_632# nfet_06v0 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=0.7u
.ends

.subckt comp018green_esd_clamp_v5p0_DVDD comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VPLUS
Xcomp018green_esd_rc_v5p0_0 comp018green_esd_rc_v5p0_0/VRC comp018green_esd_rc_v5p0_0/VPLUS
+ comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0
Xnmos_clamp_20_50_4_DVDD_0 comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VPLUS
+ a_4685_27917# nmos_clamp_20_50_4_DVDD
X0 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X1 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X2 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X3 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.88u w=5u l=0.7u
X4 a_3781_27917# a_2805_27917# comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X5 comp018green_esd_rc_v5p0_0/VMINUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X6 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X7 a_3781_27917# a_2805_27917# comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.88u w=5u l=0.7u
X8 comp018green_esd_rc_v5p0_0/VMINUS a_2805_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X9 a_3781_27917# a_2805_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X10 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X11 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X12 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X13 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X14 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X15 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X16 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X17 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X18 comp018green_esd_rc_v5p0_0/VMINUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X19 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X20 comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VRC a_2805_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X21 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X22 a_2805_27917# comp018green_esd_rc_v5p0_0/VRC comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=2.2p pd=10.88u as=2.2p ps=10.88u w=5u l=0.7u
X23 comp018green_esd_rc_v5p0_0/VMINUS a_2805_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X24 a_2805_27917# comp018green_esd_rc_v5p0_0/VRC comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.88u w=5u l=0.7u
X25 comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VRC a_2805_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X26 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X27 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X28 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X29 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X30 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=2.2p pd=10.88u as=1.3p ps=5.52u w=5u l=0.7u
X31 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X32 a_3781_27917# a_2805_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=2.2p pd=10.88u as=1.3p ps=5.52u w=5u l=0.7u
X33 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X34 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X35 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X36 comp018green_esd_rc_v5p0_0/VMINUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=2.2p pd=10.88u as=1.3p ps=5.52u w=5u l=0.7u
X37 a_3781_27917# a_2805_27917# comp018green_esd_rc_v5p0_0/VMINUS comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X38 comp018green_esd_rc_v5p0_0/VMINUS a_2805_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VMINUS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X39 a_2805_27917# comp018green_esd_rc_v5p0_0/VRC comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X40 comp018green_esd_rc_v5p0_0/VPLUS a_2805_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X41 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X42 a_4685_27917# a_3781_27917# comp018green_esd_rc_v5p0_0/VPLUS comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X43 comp018green_esd_rc_v5p0_0/VPLUS a_3781_27917# a_4685_27917# comp018green_esd_rc_v5p0_0/VPLUS pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
.ends

.subckt GF_NI_VDD_BASE DVSS DVDD VSS m3_9927_12842# m3_7265_56043# m3_5168_14436#
+ m3_7265_52842# m3_12297_33636# m3_2798_11242# m3_12297_56043# m3_2798_17636# m3_9927_1636#
+ m3_12297_52842# m3_7265_8036# m3_12861_28842# m3_9927_33636# m3_7265_4836# m3_7874_28842#
+ m3_12861_24036# m3_12861_54442# m3_10244_14436# m3_4851_27242# m3_9927_56043# m3_5168_11242#
+ m3_9927_52842# m3_7874_24036# m3_7874_54442# m3_2798_30436# m3_12861_20836# m3_12861_43242#
+ m3_5168_17636# m3_12861_41642# m3_7265_48042# m3_2481_27242# m3_7874_20836# m3_9927_8036#
+ m3_7874_43242# m3_12297_1636# m3_7874_41642# m3_4851_12842# m3_7265_44842# m3_9927_4836#
+ m3_12297_48042# m3_10244_11242# m3_5168_30436# m3_2481_12842# m3_12297_44842# m3_10244_17636#
+ m3_2481_1636# m3_2798_28842# m3_9927_48042# m3_4851_33636# m3_12297_8036# m3_12861_14436#
+ m3_2798_24036# m3_2798_54442# m3_4851_56043# m3_9927_44842# m3_12297_4836# m3_4851_52842#
+ m3_7874_14436# m3_2481_33636# m3_10244_30436# m3_2798_20836# m3_2798_43242# m3_2798_41642#
+ m3_4851_1636# m3_2481_56043# m3_5168_28842# m3_2481_8036# m3_2481_52842# m3_7265_27242#
+ m3_5168_24036# m3_2481_4836# m3_5168_54442# m3_12861_11242# m3_5168_20836# m3_5168_43242#
+ m3_12297_27242# m3_12861_17636# m3_7874_11242# m3_5168_41642# m3_4851_8036# m3_10244_28842#
+ m3_4851_48042# m3_7265_12842# m3_7874_17636# m3_4851_4836# m3_10244_24036# m3_2798_14436#
+ m3_10244_54442# m3_4851_44842# m3_9927_27242# m3_12297_12842# m3_2481_48042# VDD
+ m3_12861_30436# m3_10244_20836# m3_10244_43242# m3_7265_1636# m3_10244_41642# m3_2481_44842#
+ m3_7874_30436# m3_7265_33636#
Xcomp018green_esd_clamp_v5p0_DVDD_0 VSS VDD comp018green_esd_clamp_v5p0_DVDD
X0 VDD VSS cap_nmos_06v0 c_width=15u c_length=15u
D0 VSS VDD diode_nd2ps_06v0 pj=82u area=40p
X1 VDD VSS cap_nmos_06v0 c_width=15u c_length=15u
D1 VSS VDD diode_nd2ps_06v0 pj=82u area=40p
D2 VSS VDD diode_nd2ps_06v0 pj=82u area=40p
D3 VSS VDD diode_nd2ps_06v0 pj=82u area=40p
X2 VDD VSS cap_nmos_06v0 c_width=15u c_length=15u
X3 VDD VSS cap_nmos_06v0 c_width=15u c_length=15u
.ends

.subckt gf180mcu_ocd_io__vdd DVDD DVSS VDD VSS
X5LM_METAL_RAIL_PAD_60_0 VSS VDD VDD VSS DVSS DVDD x5LM_METAL_RAIL_PAD_60
XGF_NI_VDD_BASE_0 DVSS DVDD VSS DVSS DVSS DVDD DVSS DVSS DVDD DVSS DVDD DVSS DVSS
+ DVSS DVDD DVSS DVSS DVDD DVDD DVDD DVDD DVSS DVSS DVDD DVSS DVDD DVDD DVDD DVDD
+ DVDD DVDD DVDD DVSS DVSS DVDD DVSS DVDD DVSS DVDD DVSS DVSS DVSS DVSS DVDD DVDD
+ DVSS DVSS DVDD DVSS DVDD DVSS DVSS DVSS DVDD DVDD DVDD DVSS DVSS DVSS DVSS DVDD
+ DVSS DVDD DVDD DVDD DVDD DVSS DVSS DVDD DVSS DVSS DVSS DVDD DVSS DVDD DVDD DVDD
+ DVDD DVSS DVDD DVDD DVDD DVSS DVDD DVSS DVSS DVDD DVSS DVDD DVDD DVDD DVSS DVSS
+ DVSS DVSS VDD DVDD DVDD DVDD DVSS DVDD DVSS DVDD DVSS GF_NI_VDD_BASE
.ends

